magic
tech sky130A
magscale 1 2
timestamp 1701598240
<< obsli1 >>
rect 1104 2159 84364 85425
<< obsm1 >>
rect 934 2128 84534 85456
<< metal2 >>
rect 21362 0 21418 800
rect 64142 0 64198 800
<< obsm2 >>
rect 938 856 84530 85445
rect 938 800 21306 856
rect 21474 800 64086 856
rect 64254 800 84530 856
<< metal3 >>
rect 84743 80248 85543 80368
rect 84743 79704 85543 79824
rect 84743 79160 85543 79280
rect 84743 78616 85543 78736
rect 84743 78072 85543 78192
rect 84743 77528 85543 77648
rect 84743 76984 85543 77104
rect 84743 76440 85543 76560
rect 84743 75896 85543 76016
rect 84743 75352 85543 75472
rect 84743 74808 85543 74928
rect 84743 74264 85543 74384
rect 84743 73720 85543 73840
rect 84743 73176 85543 73296
rect 84743 72632 85543 72752
rect 84743 72088 85543 72208
rect 84743 71544 85543 71664
rect 84743 71000 85543 71120
rect 84743 70456 85543 70576
rect 84743 69912 85543 70032
rect 84743 69368 85543 69488
rect 84743 68824 85543 68944
rect 84743 68280 85543 68400
rect 84743 67736 85543 67856
rect 84743 67192 85543 67312
rect 84743 66648 85543 66768
rect 84743 66104 85543 66224
rect 0 65560 800 65680
rect 84743 65560 85543 65680
rect 84743 65016 85543 65136
rect 84743 64472 85543 64592
rect 84743 63928 85543 64048
rect 84743 63384 85543 63504
rect 84743 62840 85543 62960
rect 84743 62296 85543 62416
rect 84743 61752 85543 61872
rect 84743 61208 85543 61328
rect 84743 60664 85543 60784
rect 84743 60120 85543 60240
rect 84743 59576 85543 59696
rect 84743 59032 85543 59152
rect 84743 58488 85543 58608
rect 84743 57944 85543 58064
rect 84743 57400 85543 57520
rect 84743 56856 85543 56976
rect 84743 56312 85543 56432
rect 84743 55768 85543 55888
rect 84743 55224 85543 55344
rect 84743 54680 85543 54800
rect 84743 54136 85543 54256
rect 84743 53592 85543 53712
rect 84743 53048 85543 53168
rect 84743 52504 85543 52624
rect 84743 51960 85543 52080
rect 84743 51416 85543 51536
rect 84743 50872 85543 50992
rect 84743 50328 85543 50448
rect 84743 49784 85543 49904
rect 84743 49240 85543 49360
rect 84743 48696 85543 48816
rect 84743 48152 85543 48272
rect 84743 47608 85543 47728
rect 84743 47064 85543 47184
rect 84743 46520 85543 46640
rect 84743 45976 85543 46096
rect 84743 45432 85543 45552
rect 84743 44888 85543 45008
rect 84743 44344 85543 44464
rect 84743 43800 85543 43920
rect 84743 43256 85543 43376
rect 84743 42712 85543 42832
rect 84743 42168 85543 42288
rect 84743 41624 85543 41744
rect 84743 41080 85543 41200
rect 84743 40536 85543 40656
rect 84743 39992 85543 40112
rect 84743 39448 85543 39568
rect 84743 38904 85543 39024
rect 84743 38360 85543 38480
rect 84743 37816 85543 37936
rect 84743 37272 85543 37392
rect 84743 36728 85543 36848
rect 84743 36184 85543 36304
rect 84743 35640 85543 35760
rect 84743 35096 85543 35216
rect 84743 34552 85543 34672
rect 84743 34008 85543 34128
rect 84743 33464 85543 33584
rect 84743 32920 85543 33040
rect 84743 32376 85543 32496
rect 84743 31832 85543 31952
rect 84743 31288 85543 31408
rect 84743 30744 85543 30864
rect 84743 30200 85543 30320
rect 84743 29656 85543 29776
rect 84743 29112 85543 29232
rect 84743 28568 85543 28688
rect 84743 28024 85543 28144
rect 84743 27480 85543 27600
rect 84743 26936 85543 27056
rect 84743 26392 85543 26512
rect 84743 25848 85543 25968
rect 84743 25304 85543 25424
rect 84743 24760 85543 24880
rect 84743 24216 85543 24336
rect 84743 23672 85543 23792
rect 84743 23128 85543 23248
rect 84743 22584 85543 22704
rect 84743 22040 85543 22160
rect 0 21768 800 21888
rect 84743 21496 85543 21616
rect 84743 20952 85543 21072
rect 84743 20408 85543 20528
rect 84743 19864 85543 19984
rect 84743 19320 85543 19440
rect 84743 18776 85543 18896
rect 84743 18232 85543 18352
rect 84743 17688 85543 17808
rect 84743 17144 85543 17264
rect 84743 16600 85543 16720
rect 84743 16056 85543 16176
rect 84743 15512 85543 15632
rect 84743 14968 85543 15088
rect 84743 14424 85543 14544
rect 84743 13880 85543 14000
rect 84743 13336 85543 13456
rect 84743 12792 85543 12912
rect 84743 12248 85543 12368
rect 84743 11704 85543 11824
rect 84743 11160 85543 11280
rect 84743 10616 85543 10736
rect 84743 10072 85543 10192
rect 84743 9528 85543 9648
rect 84743 8984 85543 9104
rect 84743 8440 85543 8560
rect 84743 7896 85543 8016
rect 84743 7352 85543 7472
<< obsm3 >>
rect 800 80448 84743 85441
rect 800 80168 84663 80448
rect 800 79904 84743 80168
rect 800 79624 84663 79904
rect 800 79360 84743 79624
rect 800 79080 84663 79360
rect 800 78816 84743 79080
rect 800 78536 84663 78816
rect 800 78272 84743 78536
rect 800 77992 84663 78272
rect 800 77728 84743 77992
rect 800 77448 84663 77728
rect 800 77184 84743 77448
rect 800 76904 84663 77184
rect 800 76640 84743 76904
rect 800 76360 84663 76640
rect 800 76096 84743 76360
rect 800 75816 84663 76096
rect 800 75552 84743 75816
rect 800 75272 84663 75552
rect 800 75008 84743 75272
rect 800 74728 84663 75008
rect 800 74464 84743 74728
rect 800 74184 84663 74464
rect 800 73920 84743 74184
rect 800 73640 84663 73920
rect 800 73376 84743 73640
rect 800 73096 84663 73376
rect 800 72832 84743 73096
rect 800 72552 84663 72832
rect 800 72288 84743 72552
rect 800 72008 84663 72288
rect 800 71744 84743 72008
rect 800 71464 84663 71744
rect 800 71200 84743 71464
rect 800 70920 84663 71200
rect 800 70656 84743 70920
rect 800 70376 84663 70656
rect 800 70112 84743 70376
rect 800 69832 84663 70112
rect 800 69568 84743 69832
rect 800 69288 84663 69568
rect 800 69024 84743 69288
rect 800 68744 84663 69024
rect 800 68480 84743 68744
rect 800 68200 84663 68480
rect 800 67936 84743 68200
rect 800 67656 84663 67936
rect 800 67392 84743 67656
rect 800 67112 84663 67392
rect 800 66848 84743 67112
rect 800 66568 84663 66848
rect 800 66304 84743 66568
rect 800 66024 84663 66304
rect 800 65760 84743 66024
rect 880 65480 84663 65760
rect 800 65216 84743 65480
rect 800 64936 84663 65216
rect 800 64672 84743 64936
rect 800 64392 84663 64672
rect 800 64128 84743 64392
rect 800 63848 84663 64128
rect 800 63584 84743 63848
rect 800 63304 84663 63584
rect 800 63040 84743 63304
rect 800 62760 84663 63040
rect 800 62496 84743 62760
rect 800 62216 84663 62496
rect 800 61952 84743 62216
rect 800 61672 84663 61952
rect 800 61408 84743 61672
rect 800 61128 84663 61408
rect 800 60864 84743 61128
rect 800 60584 84663 60864
rect 800 60320 84743 60584
rect 800 60040 84663 60320
rect 800 59776 84743 60040
rect 800 59496 84663 59776
rect 800 59232 84743 59496
rect 800 58952 84663 59232
rect 800 58688 84743 58952
rect 800 58408 84663 58688
rect 800 58144 84743 58408
rect 800 57864 84663 58144
rect 800 57600 84743 57864
rect 800 57320 84663 57600
rect 800 57056 84743 57320
rect 800 56776 84663 57056
rect 800 56512 84743 56776
rect 800 56232 84663 56512
rect 800 55968 84743 56232
rect 800 55688 84663 55968
rect 800 55424 84743 55688
rect 800 55144 84663 55424
rect 800 54880 84743 55144
rect 800 54600 84663 54880
rect 800 54336 84743 54600
rect 800 54056 84663 54336
rect 800 53792 84743 54056
rect 800 53512 84663 53792
rect 800 53248 84743 53512
rect 800 52968 84663 53248
rect 800 52704 84743 52968
rect 800 52424 84663 52704
rect 800 52160 84743 52424
rect 800 51880 84663 52160
rect 800 51616 84743 51880
rect 800 51336 84663 51616
rect 800 51072 84743 51336
rect 800 50792 84663 51072
rect 800 50528 84743 50792
rect 800 50248 84663 50528
rect 800 49984 84743 50248
rect 800 49704 84663 49984
rect 800 49440 84743 49704
rect 800 49160 84663 49440
rect 800 48896 84743 49160
rect 800 48616 84663 48896
rect 800 48352 84743 48616
rect 800 48072 84663 48352
rect 800 47808 84743 48072
rect 800 47528 84663 47808
rect 800 47264 84743 47528
rect 800 46984 84663 47264
rect 800 46720 84743 46984
rect 800 46440 84663 46720
rect 800 46176 84743 46440
rect 800 45896 84663 46176
rect 800 45632 84743 45896
rect 800 45352 84663 45632
rect 800 45088 84743 45352
rect 800 44808 84663 45088
rect 800 44544 84743 44808
rect 800 44264 84663 44544
rect 800 44000 84743 44264
rect 800 43720 84663 44000
rect 800 43456 84743 43720
rect 800 43176 84663 43456
rect 800 42912 84743 43176
rect 800 42632 84663 42912
rect 800 42368 84743 42632
rect 800 42088 84663 42368
rect 800 41824 84743 42088
rect 800 41544 84663 41824
rect 800 41280 84743 41544
rect 800 41000 84663 41280
rect 800 40736 84743 41000
rect 800 40456 84663 40736
rect 800 40192 84743 40456
rect 800 39912 84663 40192
rect 800 39648 84743 39912
rect 800 39368 84663 39648
rect 800 39104 84743 39368
rect 800 38824 84663 39104
rect 800 38560 84743 38824
rect 800 38280 84663 38560
rect 800 38016 84743 38280
rect 800 37736 84663 38016
rect 800 37472 84743 37736
rect 800 37192 84663 37472
rect 800 36928 84743 37192
rect 800 36648 84663 36928
rect 800 36384 84743 36648
rect 800 36104 84663 36384
rect 800 35840 84743 36104
rect 800 35560 84663 35840
rect 800 35296 84743 35560
rect 800 35016 84663 35296
rect 800 34752 84743 35016
rect 800 34472 84663 34752
rect 800 34208 84743 34472
rect 800 33928 84663 34208
rect 800 33664 84743 33928
rect 800 33384 84663 33664
rect 800 33120 84743 33384
rect 800 32840 84663 33120
rect 800 32576 84743 32840
rect 800 32296 84663 32576
rect 800 32032 84743 32296
rect 800 31752 84663 32032
rect 800 31488 84743 31752
rect 800 31208 84663 31488
rect 800 30944 84743 31208
rect 800 30664 84663 30944
rect 800 30400 84743 30664
rect 800 30120 84663 30400
rect 800 29856 84743 30120
rect 800 29576 84663 29856
rect 800 29312 84743 29576
rect 800 29032 84663 29312
rect 800 28768 84743 29032
rect 800 28488 84663 28768
rect 800 28224 84743 28488
rect 800 27944 84663 28224
rect 800 27680 84743 27944
rect 800 27400 84663 27680
rect 800 27136 84743 27400
rect 800 26856 84663 27136
rect 800 26592 84743 26856
rect 800 26312 84663 26592
rect 800 26048 84743 26312
rect 800 25768 84663 26048
rect 800 25504 84743 25768
rect 800 25224 84663 25504
rect 800 24960 84743 25224
rect 800 24680 84663 24960
rect 800 24416 84743 24680
rect 800 24136 84663 24416
rect 800 23872 84743 24136
rect 800 23592 84663 23872
rect 800 23328 84743 23592
rect 800 23048 84663 23328
rect 800 22784 84743 23048
rect 800 22504 84663 22784
rect 800 22240 84743 22504
rect 800 21968 84663 22240
rect 880 21960 84663 21968
rect 880 21696 84743 21960
rect 880 21688 84663 21696
rect 800 21416 84663 21688
rect 800 21152 84743 21416
rect 800 20872 84663 21152
rect 800 20608 84743 20872
rect 800 20328 84663 20608
rect 800 20064 84743 20328
rect 800 19784 84663 20064
rect 800 19520 84743 19784
rect 800 19240 84663 19520
rect 800 18976 84743 19240
rect 800 18696 84663 18976
rect 800 18432 84743 18696
rect 800 18152 84663 18432
rect 800 17888 84743 18152
rect 800 17608 84663 17888
rect 800 17344 84743 17608
rect 800 17064 84663 17344
rect 800 16800 84743 17064
rect 800 16520 84663 16800
rect 800 16256 84743 16520
rect 800 15976 84663 16256
rect 800 15712 84743 15976
rect 800 15432 84663 15712
rect 800 15168 84743 15432
rect 800 14888 84663 15168
rect 800 14624 84743 14888
rect 800 14344 84663 14624
rect 800 14080 84743 14344
rect 800 13800 84663 14080
rect 800 13536 84743 13800
rect 800 13256 84663 13536
rect 800 12992 84743 13256
rect 800 12712 84663 12992
rect 800 12448 84743 12712
rect 800 12168 84663 12448
rect 800 11904 84743 12168
rect 800 11624 84663 11904
rect 800 11360 84743 11624
rect 800 11080 84663 11360
rect 800 10816 84743 11080
rect 800 10536 84663 10816
rect 800 10272 84743 10536
rect 800 9992 84663 10272
rect 800 9728 84743 9992
rect 800 9448 84663 9728
rect 800 9184 84743 9448
rect 800 8904 84663 9184
rect 800 8640 84743 8904
rect 800 8360 84663 8640
rect 800 8096 84743 8360
rect 800 7816 84663 8096
rect 800 7552 84743 7816
rect 800 7272 84663 7552
rect 800 2143 84743 7272
<< metal4 >>
rect 4208 2128 4528 85456
rect 19568 2128 19888 85456
rect 34928 2128 35248 85456
rect 50288 2128 50608 85456
rect 65648 2128 65968 85456
rect 81008 2128 81328 85456
<< obsm4 >>
rect 49371 13907 50208 53957
rect 50688 13907 65568 53957
rect 66048 13907 80928 53957
rect 81408 13907 82741 53957
<< labels >>
rlabel metal4 s 19568 2128 19888 85456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 85456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 85456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 85456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 85456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 85456 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 21362 0 21418 800 6 clk
port 3 nsew signal input
rlabel metal3 s 84743 45432 85543 45552 6 reg_dat_di[0]
port 4 nsew signal input
rlabel metal3 s 84743 50872 85543 50992 6 reg_dat_di[10]
port 5 nsew signal input
rlabel metal3 s 84743 51416 85543 51536 6 reg_dat_di[11]
port 6 nsew signal input
rlabel metal3 s 84743 51960 85543 52080 6 reg_dat_di[12]
port 7 nsew signal input
rlabel metal3 s 84743 52504 85543 52624 6 reg_dat_di[13]
port 8 nsew signal input
rlabel metal3 s 84743 53048 85543 53168 6 reg_dat_di[14]
port 9 nsew signal input
rlabel metal3 s 84743 53592 85543 53712 6 reg_dat_di[15]
port 10 nsew signal input
rlabel metal3 s 84743 54136 85543 54256 6 reg_dat_di[16]
port 11 nsew signal input
rlabel metal3 s 84743 54680 85543 54800 6 reg_dat_di[17]
port 12 nsew signal input
rlabel metal3 s 84743 55224 85543 55344 6 reg_dat_di[18]
port 13 nsew signal input
rlabel metal3 s 84743 55768 85543 55888 6 reg_dat_di[19]
port 14 nsew signal input
rlabel metal3 s 84743 45976 85543 46096 6 reg_dat_di[1]
port 15 nsew signal input
rlabel metal3 s 84743 56312 85543 56432 6 reg_dat_di[20]
port 16 nsew signal input
rlabel metal3 s 84743 56856 85543 56976 6 reg_dat_di[21]
port 17 nsew signal input
rlabel metal3 s 84743 57400 85543 57520 6 reg_dat_di[22]
port 18 nsew signal input
rlabel metal3 s 84743 57944 85543 58064 6 reg_dat_di[23]
port 19 nsew signal input
rlabel metal3 s 84743 58488 85543 58608 6 reg_dat_di[24]
port 20 nsew signal input
rlabel metal3 s 84743 59032 85543 59152 6 reg_dat_di[25]
port 21 nsew signal input
rlabel metal3 s 84743 59576 85543 59696 6 reg_dat_di[26]
port 22 nsew signal input
rlabel metal3 s 84743 60120 85543 60240 6 reg_dat_di[27]
port 23 nsew signal input
rlabel metal3 s 84743 60664 85543 60784 6 reg_dat_di[28]
port 24 nsew signal input
rlabel metal3 s 84743 61208 85543 61328 6 reg_dat_di[29]
port 25 nsew signal input
rlabel metal3 s 84743 46520 85543 46640 6 reg_dat_di[2]
port 26 nsew signal input
rlabel metal3 s 84743 61752 85543 61872 6 reg_dat_di[30]
port 27 nsew signal input
rlabel metal3 s 84743 62296 85543 62416 6 reg_dat_di[31]
port 28 nsew signal input
rlabel metal3 s 84743 47064 85543 47184 6 reg_dat_di[3]
port 29 nsew signal input
rlabel metal3 s 84743 47608 85543 47728 6 reg_dat_di[4]
port 30 nsew signal input
rlabel metal3 s 84743 48152 85543 48272 6 reg_dat_di[5]
port 31 nsew signal input
rlabel metal3 s 84743 48696 85543 48816 6 reg_dat_di[6]
port 32 nsew signal input
rlabel metal3 s 84743 49240 85543 49360 6 reg_dat_di[7]
port 33 nsew signal input
rlabel metal3 s 84743 49784 85543 49904 6 reg_dat_di[8]
port 34 nsew signal input
rlabel metal3 s 84743 50328 85543 50448 6 reg_dat_di[9]
port 35 nsew signal input
rlabel metal3 s 84743 62840 85543 62960 6 reg_dat_do[0]
port 36 nsew signal output
rlabel metal3 s 84743 68280 85543 68400 6 reg_dat_do[10]
port 37 nsew signal output
rlabel metal3 s 84743 68824 85543 68944 6 reg_dat_do[11]
port 38 nsew signal output
rlabel metal3 s 84743 69368 85543 69488 6 reg_dat_do[12]
port 39 nsew signal output
rlabel metal3 s 84743 69912 85543 70032 6 reg_dat_do[13]
port 40 nsew signal output
rlabel metal3 s 84743 70456 85543 70576 6 reg_dat_do[14]
port 41 nsew signal output
rlabel metal3 s 84743 71000 85543 71120 6 reg_dat_do[15]
port 42 nsew signal output
rlabel metal3 s 84743 71544 85543 71664 6 reg_dat_do[16]
port 43 nsew signal output
rlabel metal3 s 84743 72088 85543 72208 6 reg_dat_do[17]
port 44 nsew signal output
rlabel metal3 s 84743 72632 85543 72752 6 reg_dat_do[18]
port 45 nsew signal output
rlabel metal3 s 84743 73176 85543 73296 6 reg_dat_do[19]
port 46 nsew signal output
rlabel metal3 s 84743 63384 85543 63504 6 reg_dat_do[1]
port 47 nsew signal output
rlabel metal3 s 84743 73720 85543 73840 6 reg_dat_do[20]
port 48 nsew signal output
rlabel metal3 s 84743 74264 85543 74384 6 reg_dat_do[21]
port 49 nsew signal output
rlabel metal3 s 84743 74808 85543 74928 6 reg_dat_do[22]
port 50 nsew signal output
rlabel metal3 s 84743 75352 85543 75472 6 reg_dat_do[23]
port 51 nsew signal output
rlabel metal3 s 84743 75896 85543 76016 6 reg_dat_do[24]
port 52 nsew signal output
rlabel metal3 s 84743 76440 85543 76560 6 reg_dat_do[25]
port 53 nsew signal output
rlabel metal3 s 84743 76984 85543 77104 6 reg_dat_do[26]
port 54 nsew signal output
rlabel metal3 s 84743 77528 85543 77648 6 reg_dat_do[27]
port 55 nsew signal output
rlabel metal3 s 84743 78072 85543 78192 6 reg_dat_do[28]
port 56 nsew signal output
rlabel metal3 s 84743 78616 85543 78736 6 reg_dat_do[29]
port 57 nsew signal output
rlabel metal3 s 84743 63928 85543 64048 6 reg_dat_do[2]
port 58 nsew signal output
rlabel metal3 s 84743 79160 85543 79280 6 reg_dat_do[30]
port 59 nsew signal output
rlabel metal3 s 84743 79704 85543 79824 6 reg_dat_do[31]
port 60 nsew signal output
rlabel metal3 s 84743 64472 85543 64592 6 reg_dat_do[3]
port 61 nsew signal output
rlabel metal3 s 84743 65016 85543 65136 6 reg_dat_do[4]
port 62 nsew signal output
rlabel metal3 s 84743 65560 85543 65680 6 reg_dat_do[5]
port 63 nsew signal output
rlabel metal3 s 84743 66104 85543 66224 6 reg_dat_do[6]
port 64 nsew signal output
rlabel metal3 s 84743 66648 85543 66768 6 reg_dat_do[7]
port 65 nsew signal output
rlabel metal3 s 84743 67192 85543 67312 6 reg_dat_do[8]
port 66 nsew signal output
rlabel metal3 s 84743 67736 85543 67856 6 reg_dat_do[9]
port 67 nsew signal output
rlabel metal3 s 84743 44888 85543 45008 6 reg_dat_re
port 68 nsew signal input
rlabel metal3 s 84743 80248 85543 80368 6 reg_dat_wait
port 69 nsew signal output
rlabel metal3 s 84743 44344 85543 44464 6 reg_dat_we
port 70 nsew signal input
rlabel metal3 s 84743 9528 85543 9648 6 reg_div_di[0]
port 71 nsew signal input
rlabel metal3 s 84743 14968 85543 15088 6 reg_div_di[10]
port 72 nsew signal input
rlabel metal3 s 84743 15512 85543 15632 6 reg_div_di[11]
port 73 nsew signal input
rlabel metal3 s 84743 16056 85543 16176 6 reg_div_di[12]
port 74 nsew signal input
rlabel metal3 s 84743 16600 85543 16720 6 reg_div_di[13]
port 75 nsew signal input
rlabel metal3 s 84743 17144 85543 17264 6 reg_div_di[14]
port 76 nsew signal input
rlabel metal3 s 84743 17688 85543 17808 6 reg_div_di[15]
port 77 nsew signal input
rlabel metal3 s 84743 18232 85543 18352 6 reg_div_di[16]
port 78 nsew signal input
rlabel metal3 s 84743 18776 85543 18896 6 reg_div_di[17]
port 79 nsew signal input
rlabel metal3 s 84743 19320 85543 19440 6 reg_div_di[18]
port 80 nsew signal input
rlabel metal3 s 84743 19864 85543 19984 6 reg_div_di[19]
port 81 nsew signal input
rlabel metal3 s 84743 10072 85543 10192 6 reg_div_di[1]
port 82 nsew signal input
rlabel metal3 s 84743 20408 85543 20528 6 reg_div_di[20]
port 83 nsew signal input
rlabel metal3 s 84743 20952 85543 21072 6 reg_div_di[21]
port 84 nsew signal input
rlabel metal3 s 84743 21496 85543 21616 6 reg_div_di[22]
port 85 nsew signal input
rlabel metal3 s 84743 22040 85543 22160 6 reg_div_di[23]
port 86 nsew signal input
rlabel metal3 s 84743 22584 85543 22704 6 reg_div_di[24]
port 87 nsew signal input
rlabel metal3 s 84743 23128 85543 23248 6 reg_div_di[25]
port 88 nsew signal input
rlabel metal3 s 84743 23672 85543 23792 6 reg_div_di[26]
port 89 nsew signal input
rlabel metal3 s 84743 24216 85543 24336 6 reg_div_di[27]
port 90 nsew signal input
rlabel metal3 s 84743 24760 85543 24880 6 reg_div_di[28]
port 91 nsew signal input
rlabel metal3 s 84743 25304 85543 25424 6 reg_div_di[29]
port 92 nsew signal input
rlabel metal3 s 84743 10616 85543 10736 6 reg_div_di[2]
port 93 nsew signal input
rlabel metal3 s 84743 25848 85543 25968 6 reg_div_di[30]
port 94 nsew signal input
rlabel metal3 s 84743 26392 85543 26512 6 reg_div_di[31]
port 95 nsew signal input
rlabel metal3 s 84743 11160 85543 11280 6 reg_div_di[3]
port 96 nsew signal input
rlabel metal3 s 84743 11704 85543 11824 6 reg_div_di[4]
port 97 nsew signal input
rlabel metal3 s 84743 12248 85543 12368 6 reg_div_di[5]
port 98 nsew signal input
rlabel metal3 s 84743 12792 85543 12912 6 reg_div_di[6]
port 99 nsew signal input
rlabel metal3 s 84743 13336 85543 13456 6 reg_div_di[7]
port 100 nsew signal input
rlabel metal3 s 84743 13880 85543 14000 6 reg_div_di[8]
port 101 nsew signal input
rlabel metal3 s 84743 14424 85543 14544 6 reg_div_di[9]
port 102 nsew signal input
rlabel metal3 s 84743 26936 85543 27056 6 reg_div_do[0]
port 103 nsew signal output
rlabel metal3 s 84743 32376 85543 32496 6 reg_div_do[10]
port 104 nsew signal output
rlabel metal3 s 84743 32920 85543 33040 6 reg_div_do[11]
port 105 nsew signal output
rlabel metal3 s 84743 33464 85543 33584 6 reg_div_do[12]
port 106 nsew signal output
rlabel metal3 s 84743 34008 85543 34128 6 reg_div_do[13]
port 107 nsew signal output
rlabel metal3 s 84743 34552 85543 34672 6 reg_div_do[14]
port 108 nsew signal output
rlabel metal3 s 84743 35096 85543 35216 6 reg_div_do[15]
port 109 nsew signal output
rlabel metal3 s 84743 35640 85543 35760 6 reg_div_do[16]
port 110 nsew signal output
rlabel metal3 s 84743 36184 85543 36304 6 reg_div_do[17]
port 111 nsew signal output
rlabel metal3 s 84743 36728 85543 36848 6 reg_div_do[18]
port 112 nsew signal output
rlabel metal3 s 84743 37272 85543 37392 6 reg_div_do[19]
port 113 nsew signal output
rlabel metal3 s 84743 27480 85543 27600 6 reg_div_do[1]
port 114 nsew signal output
rlabel metal3 s 84743 37816 85543 37936 6 reg_div_do[20]
port 115 nsew signal output
rlabel metal3 s 84743 38360 85543 38480 6 reg_div_do[21]
port 116 nsew signal output
rlabel metal3 s 84743 38904 85543 39024 6 reg_div_do[22]
port 117 nsew signal output
rlabel metal3 s 84743 39448 85543 39568 6 reg_div_do[23]
port 118 nsew signal output
rlabel metal3 s 84743 39992 85543 40112 6 reg_div_do[24]
port 119 nsew signal output
rlabel metal3 s 84743 40536 85543 40656 6 reg_div_do[25]
port 120 nsew signal output
rlabel metal3 s 84743 41080 85543 41200 6 reg_div_do[26]
port 121 nsew signal output
rlabel metal3 s 84743 41624 85543 41744 6 reg_div_do[27]
port 122 nsew signal output
rlabel metal3 s 84743 42168 85543 42288 6 reg_div_do[28]
port 123 nsew signal output
rlabel metal3 s 84743 42712 85543 42832 6 reg_div_do[29]
port 124 nsew signal output
rlabel metal3 s 84743 28024 85543 28144 6 reg_div_do[2]
port 125 nsew signal output
rlabel metal3 s 84743 43256 85543 43376 6 reg_div_do[30]
port 126 nsew signal output
rlabel metal3 s 84743 43800 85543 43920 6 reg_div_do[31]
port 127 nsew signal output
rlabel metal3 s 84743 28568 85543 28688 6 reg_div_do[3]
port 128 nsew signal output
rlabel metal3 s 84743 29112 85543 29232 6 reg_div_do[4]
port 129 nsew signal output
rlabel metal3 s 84743 29656 85543 29776 6 reg_div_do[5]
port 130 nsew signal output
rlabel metal3 s 84743 30200 85543 30320 6 reg_div_do[6]
port 131 nsew signal output
rlabel metal3 s 84743 30744 85543 30864 6 reg_div_do[7]
port 132 nsew signal output
rlabel metal3 s 84743 31288 85543 31408 6 reg_div_do[8]
port 133 nsew signal output
rlabel metal3 s 84743 31832 85543 31952 6 reg_div_do[9]
port 134 nsew signal output
rlabel metal3 s 84743 7352 85543 7472 6 reg_div_we[0]
port 135 nsew signal input
rlabel metal3 s 84743 7896 85543 8016 6 reg_div_we[1]
port 136 nsew signal input
rlabel metal3 s 84743 8440 85543 8560 6 reg_div_we[2]
port 137 nsew signal input
rlabel metal3 s 84743 8984 85543 9104 6 reg_div_we[3]
port 138 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 resetn
port 139 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 ser_rx
port 140 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 ser_tx
port 141 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 85543 87687
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4772578
string GDS_FILE /openlane/designs/simpleuart/runs/RUN_2023.12.03_10.07.08/results/signoff/simpleuart.magic.gds
string GDS_START 477138
<< end >>

