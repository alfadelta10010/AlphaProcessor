magic
tech sky130A
magscale 1 2
timestamp 1701597199
<< obsli1 >>
rect 1104 2159 96232 96849
<< obsm1 >>
rect 290 2128 96494 98864
<< metal2 >>
rect 4986 98721 5042 99521
rect 5354 98721 5410 99521
rect 5722 98721 5778 99521
rect 6090 98721 6146 99521
rect 6458 98721 6514 99521
rect 6826 98721 6882 99521
rect 7194 98721 7250 99521
rect 7562 98721 7618 99521
rect 7930 98721 7986 99521
rect 8298 98721 8354 99521
rect 8666 98721 8722 99521
rect 9034 98721 9090 99521
rect 9402 98721 9458 99521
rect 9770 98721 9826 99521
rect 10138 98721 10194 99521
rect 10506 98721 10562 99521
rect 10874 98721 10930 99521
rect 11242 98721 11298 99521
rect 11610 98721 11666 99521
rect 11978 98721 12034 99521
rect 12346 98721 12402 99521
rect 12714 98721 12770 99521
rect 13082 98721 13138 99521
rect 13450 98721 13506 99521
rect 13818 98721 13874 99521
rect 14186 98721 14242 99521
rect 14554 98721 14610 99521
rect 14922 98721 14978 99521
rect 15290 98721 15346 99521
rect 15658 98721 15714 99521
rect 16026 98721 16082 99521
rect 16394 98721 16450 99521
rect 16762 98721 16818 99521
rect 17130 98721 17186 99521
rect 17498 98721 17554 99521
rect 17866 98721 17922 99521
rect 18234 98721 18290 99521
rect 18602 98721 18658 99521
rect 18970 98721 19026 99521
rect 19338 98721 19394 99521
rect 19706 98721 19762 99521
rect 20074 98721 20130 99521
rect 20442 98721 20498 99521
rect 20810 98721 20866 99521
rect 21178 98721 21234 99521
rect 21546 98721 21602 99521
rect 21914 98721 21970 99521
rect 22282 98721 22338 99521
rect 22650 98721 22706 99521
rect 23018 98721 23074 99521
rect 23386 98721 23442 99521
rect 23754 98721 23810 99521
rect 24122 98721 24178 99521
rect 24490 98721 24546 99521
rect 24858 98721 24914 99521
rect 25226 98721 25282 99521
rect 25594 98721 25650 99521
rect 25962 98721 26018 99521
rect 26330 98721 26386 99521
rect 26698 98721 26754 99521
rect 27066 98721 27122 99521
rect 27434 98721 27490 99521
rect 27802 98721 27858 99521
rect 28170 98721 28226 99521
rect 28538 98721 28594 99521
rect 28906 98721 28962 99521
rect 29274 98721 29330 99521
rect 29642 98721 29698 99521
rect 30010 98721 30066 99521
rect 30378 98721 30434 99521
rect 30746 98721 30802 99521
rect 31114 98721 31170 99521
rect 31482 98721 31538 99521
rect 31850 98721 31906 99521
rect 32218 98721 32274 99521
rect 32586 98721 32642 99521
rect 32954 98721 33010 99521
rect 33322 98721 33378 99521
rect 33690 98721 33746 99521
rect 34058 98721 34114 99521
rect 34426 98721 34482 99521
rect 34794 98721 34850 99521
rect 35162 98721 35218 99521
rect 35530 98721 35586 99521
rect 35898 98721 35954 99521
rect 36266 98721 36322 99521
rect 36634 98721 36690 99521
rect 37002 98721 37058 99521
rect 37370 98721 37426 99521
rect 37738 98721 37794 99521
rect 38106 98721 38162 99521
rect 38474 98721 38530 99521
rect 38842 98721 38898 99521
rect 39210 98721 39266 99521
rect 39578 98721 39634 99521
rect 39946 98721 40002 99521
rect 40314 98721 40370 99521
rect 40682 98721 40738 99521
rect 41050 98721 41106 99521
rect 41418 98721 41474 99521
rect 41786 98721 41842 99521
rect 42154 98721 42210 99521
rect 42522 98721 42578 99521
rect 42890 98721 42946 99521
rect 43258 98721 43314 99521
rect 43626 98721 43682 99521
rect 43994 98721 44050 99521
rect 44362 98721 44418 99521
rect 44730 98721 44786 99521
rect 45098 98721 45154 99521
rect 45466 98721 45522 99521
rect 45834 98721 45890 99521
rect 46202 98721 46258 99521
rect 46570 98721 46626 99521
rect 46938 98721 46994 99521
rect 47306 98721 47362 99521
rect 47674 98721 47730 99521
rect 48042 98721 48098 99521
rect 48410 98721 48466 99521
rect 48778 98721 48834 99521
rect 49146 98721 49202 99521
rect 49514 98721 49570 99521
rect 49882 98721 49938 99521
rect 50250 98721 50306 99521
rect 50618 98721 50674 99521
rect 50986 98721 51042 99521
rect 51354 98721 51410 99521
rect 51722 98721 51778 99521
rect 52090 98721 52146 99521
rect 52458 98721 52514 99521
rect 52826 98721 52882 99521
rect 53194 98721 53250 99521
rect 53562 98721 53618 99521
rect 53930 98721 53986 99521
rect 54298 98721 54354 99521
rect 54666 98721 54722 99521
rect 55034 98721 55090 99521
rect 55402 98721 55458 99521
rect 55770 98721 55826 99521
rect 56138 98721 56194 99521
rect 56506 98721 56562 99521
rect 56874 98721 56930 99521
rect 57242 98721 57298 99521
rect 57610 98721 57666 99521
rect 57978 98721 58034 99521
rect 58346 98721 58402 99521
rect 58714 98721 58770 99521
rect 59082 98721 59138 99521
rect 59450 98721 59506 99521
rect 59818 98721 59874 99521
rect 60186 98721 60242 99521
rect 60554 98721 60610 99521
rect 60922 98721 60978 99521
rect 61290 98721 61346 99521
rect 61658 98721 61714 99521
rect 62026 98721 62082 99521
rect 62394 98721 62450 99521
rect 62762 98721 62818 99521
rect 63130 98721 63186 99521
rect 63498 98721 63554 99521
rect 63866 98721 63922 99521
rect 64234 98721 64290 99521
rect 64602 98721 64658 99521
rect 64970 98721 65026 99521
rect 65338 98721 65394 99521
rect 65706 98721 65762 99521
rect 66074 98721 66130 99521
rect 66442 98721 66498 99521
rect 66810 98721 66866 99521
rect 67178 98721 67234 99521
rect 67546 98721 67602 99521
rect 67914 98721 67970 99521
rect 68282 98721 68338 99521
rect 68650 98721 68706 99521
rect 69018 98721 69074 99521
rect 69386 98721 69442 99521
rect 69754 98721 69810 99521
rect 70122 98721 70178 99521
rect 70490 98721 70546 99521
rect 70858 98721 70914 99521
rect 71226 98721 71282 99521
rect 71594 98721 71650 99521
rect 71962 98721 72018 99521
rect 72330 98721 72386 99521
rect 72698 98721 72754 99521
rect 73066 98721 73122 99521
rect 73434 98721 73490 99521
rect 73802 98721 73858 99521
rect 74170 98721 74226 99521
rect 74538 98721 74594 99521
rect 74906 98721 74962 99521
rect 75274 98721 75330 99521
rect 75642 98721 75698 99521
rect 76010 98721 76066 99521
rect 76378 98721 76434 99521
rect 76746 98721 76802 99521
rect 77114 98721 77170 99521
rect 77482 98721 77538 99521
rect 77850 98721 77906 99521
rect 78218 98721 78274 99521
rect 78586 98721 78642 99521
rect 78954 98721 79010 99521
rect 79322 98721 79378 99521
rect 79690 98721 79746 99521
rect 80058 98721 80114 99521
rect 80426 98721 80482 99521
rect 80794 98721 80850 99521
rect 81162 98721 81218 99521
rect 81530 98721 81586 99521
rect 81898 98721 81954 99521
rect 82266 98721 82322 99521
rect 82634 98721 82690 99521
rect 83002 98721 83058 99521
rect 83370 98721 83426 99521
rect 83738 98721 83794 99521
rect 84106 98721 84162 99521
rect 84474 98721 84530 99521
rect 84842 98721 84898 99521
rect 85210 98721 85266 99521
rect 85578 98721 85634 99521
rect 85946 98721 86002 99521
rect 86314 98721 86370 99521
rect 86682 98721 86738 99521
rect 87050 98721 87106 99521
rect 87418 98721 87474 99521
rect 87786 98721 87842 99521
rect 88154 98721 88210 99521
rect 88522 98721 88578 99521
rect 88890 98721 88946 99521
rect 89258 98721 89314 99521
rect 89626 98721 89682 99521
rect 89994 98721 90050 99521
rect 90362 98721 90418 99521
rect 90730 98721 90786 99521
rect 91098 98721 91154 99521
rect 91466 98721 91522 99521
rect 91834 98721 91890 99521
rect 92202 98721 92258 99521
rect 24306 0 24362 800
rect 72974 0 73030 800
<< obsm2 >>
rect 296 98665 4930 98870
rect 5098 98665 5298 98870
rect 5466 98665 5666 98870
rect 5834 98665 6034 98870
rect 6202 98665 6402 98870
rect 6570 98665 6770 98870
rect 6938 98665 7138 98870
rect 7306 98665 7506 98870
rect 7674 98665 7874 98870
rect 8042 98665 8242 98870
rect 8410 98665 8610 98870
rect 8778 98665 8978 98870
rect 9146 98665 9346 98870
rect 9514 98665 9714 98870
rect 9882 98665 10082 98870
rect 10250 98665 10450 98870
rect 10618 98665 10818 98870
rect 10986 98665 11186 98870
rect 11354 98665 11554 98870
rect 11722 98665 11922 98870
rect 12090 98665 12290 98870
rect 12458 98665 12658 98870
rect 12826 98665 13026 98870
rect 13194 98665 13394 98870
rect 13562 98665 13762 98870
rect 13930 98665 14130 98870
rect 14298 98665 14498 98870
rect 14666 98665 14866 98870
rect 15034 98665 15234 98870
rect 15402 98665 15602 98870
rect 15770 98665 15970 98870
rect 16138 98665 16338 98870
rect 16506 98665 16706 98870
rect 16874 98665 17074 98870
rect 17242 98665 17442 98870
rect 17610 98665 17810 98870
rect 17978 98665 18178 98870
rect 18346 98665 18546 98870
rect 18714 98665 18914 98870
rect 19082 98665 19282 98870
rect 19450 98665 19650 98870
rect 19818 98665 20018 98870
rect 20186 98665 20386 98870
rect 20554 98665 20754 98870
rect 20922 98665 21122 98870
rect 21290 98665 21490 98870
rect 21658 98665 21858 98870
rect 22026 98665 22226 98870
rect 22394 98665 22594 98870
rect 22762 98665 22962 98870
rect 23130 98665 23330 98870
rect 23498 98665 23698 98870
rect 23866 98665 24066 98870
rect 24234 98665 24434 98870
rect 24602 98665 24802 98870
rect 24970 98665 25170 98870
rect 25338 98665 25538 98870
rect 25706 98665 25906 98870
rect 26074 98665 26274 98870
rect 26442 98665 26642 98870
rect 26810 98665 27010 98870
rect 27178 98665 27378 98870
rect 27546 98665 27746 98870
rect 27914 98665 28114 98870
rect 28282 98665 28482 98870
rect 28650 98665 28850 98870
rect 29018 98665 29218 98870
rect 29386 98665 29586 98870
rect 29754 98665 29954 98870
rect 30122 98665 30322 98870
rect 30490 98665 30690 98870
rect 30858 98665 31058 98870
rect 31226 98665 31426 98870
rect 31594 98665 31794 98870
rect 31962 98665 32162 98870
rect 32330 98665 32530 98870
rect 32698 98665 32898 98870
rect 33066 98665 33266 98870
rect 33434 98665 33634 98870
rect 33802 98665 34002 98870
rect 34170 98665 34370 98870
rect 34538 98665 34738 98870
rect 34906 98665 35106 98870
rect 35274 98665 35474 98870
rect 35642 98665 35842 98870
rect 36010 98665 36210 98870
rect 36378 98665 36578 98870
rect 36746 98665 36946 98870
rect 37114 98665 37314 98870
rect 37482 98665 37682 98870
rect 37850 98665 38050 98870
rect 38218 98665 38418 98870
rect 38586 98665 38786 98870
rect 38954 98665 39154 98870
rect 39322 98665 39522 98870
rect 39690 98665 39890 98870
rect 40058 98665 40258 98870
rect 40426 98665 40626 98870
rect 40794 98665 40994 98870
rect 41162 98665 41362 98870
rect 41530 98665 41730 98870
rect 41898 98665 42098 98870
rect 42266 98665 42466 98870
rect 42634 98665 42834 98870
rect 43002 98665 43202 98870
rect 43370 98665 43570 98870
rect 43738 98665 43938 98870
rect 44106 98665 44306 98870
rect 44474 98665 44674 98870
rect 44842 98665 45042 98870
rect 45210 98665 45410 98870
rect 45578 98665 45778 98870
rect 45946 98665 46146 98870
rect 46314 98665 46514 98870
rect 46682 98665 46882 98870
rect 47050 98665 47250 98870
rect 47418 98665 47618 98870
rect 47786 98665 47986 98870
rect 48154 98665 48354 98870
rect 48522 98665 48722 98870
rect 48890 98665 49090 98870
rect 49258 98665 49458 98870
rect 49626 98665 49826 98870
rect 49994 98665 50194 98870
rect 50362 98665 50562 98870
rect 50730 98665 50930 98870
rect 51098 98665 51298 98870
rect 51466 98665 51666 98870
rect 51834 98665 52034 98870
rect 52202 98665 52402 98870
rect 52570 98665 52770 98870
rect 52938 98665 53138 98870
rect 53306 98665 53506 98870
rect 53674 98665 53874 98870
rect 54042 98665 54242 98870
rect 54410 98665 54610 98870
rect 54778 98665 54978 98870
rect 55146 98665 55346 98870
rect 55514 98665 55714 98870
rect 55882 98665 56082 98870
rect 56250 98665 56450 98870
rect 56618 98665 56818 98870
rect 56986 98665 57186 98870
rect 57354 98665 57554 98870
rect 57722 98665 57922 98870
rect 58090 98665 58290 98870
rect 58458 98665 58658 98870
rect 58826 98665 59026 98870
rect 59194 98665 59394 98870
rect 59562 98665 59762 98870
rect 59930 98665 60130 98870
rect 60298 98665 60498 98870
rect 60666 98665 60866 98870
rect 61034 98665 61234 98870
rect 61402 98665 61602 98870
rect 61770 98665 61970 98870
rect 62138 98665 62338 98870
rect 62506 98665 62706 98870
rect 62874 98665 63074 98870
rect 63242 98665 63442 98870
rect 63610 98665 63810 98870
rect 63978 98665 64178 98870
rect 64346 98665 64546 98870
rect 64714 98665 64914 98870
rect 65082 98665 65282 98870
rect 65450 98665 65650 98870
rect 65818 98665 66018 98870
rect 66186 98665 66386 98870
rect 66554 98665 66754 98870
rect 66922 98665 67122 98870
rect 67290 98665 67490 98870
rect 67658 98665 67858 98870
rect 68026 98665 68226 98870
rect 68394 98665 68594 98870
rect 68762 98665 68962 98870
rect 69130 98665 69330 98870
rect 69498 98665 69698 98870
rect 69866 98665 70066 98870
rect 70234 98665 70434 98870
rect 70602 98665 70802 98870
rect 70970 98665 71170 98870
rect 71338 98665 71538 98870
rect 71706 98665 71906 98870
rect 72074 98665 72274 98870
rect 72442 98665 72642 98870
rect 72810 98665 73010 98870
rect 73178 98665 73378 98870
rect 73546 98665 73746 98870
rect 73914 98665 74114 98870
rect 74282 98665 74482 98870
rect 74650 98665 74850 98870
rect 75018 98665 75218 98870
rect 75386 98665 75586 98870
rect 75754 98665 75954 98870
rect 76122 98665 76322 98870
rect 76490 98665 76690 98870
rect 76858 98665 77058 98870
rect 77226 98665 77426 98870
rect 77594 98665 77794 98870
rect 77962 98665 78162 98870
rect 78330 98665 78530 98870
rect 78698 98665 78898 98870
rect 79066 98665 79266 98870
rect 79434 98665 79634 98870
rect 79802 98665 80002 98870
rect 80170 98665 80370 98870
rect 80538 98665 80738 98870
rect 80906 98665 81106 98870
rect 81274 98665 81474 98870
rect 81642 98665 81842 98870
rect 82010 98665 82210 98870
rect 82378 98665 82578 98870
rect 82746 98665 82946 98870
rect 83114 98665 83314 98870
rect 83482 98665 83682 98870
rect 83850 98665 84050 98870
rect 84218 98665 84418 98870
rect 84586 98665 84786 98870
rect 84954 98665 85154 98870
rect 85322 98665 85522 98870
rect 85690 98665 85890 98870
rect 86058 98665 86258 98870
rect 86426 98665 86626 98870
rect 86794 98665 86994 98870
rect 87162 98665 87362 98870
rect 87530 98665 87730 98870
rect 87898 98665 88098 98870
rect 88266 98665 88466 98870
rect 88634 98665 88834 98870
rect 89002 98665 89202 98870
rect 89370 98665 89570 98870
rect 89738 98665 89938 98870
rect 90106 98665 90306 98870
rect 90474 98665 90674 98870
rect 90842 98665 91042 98870
rect 91210 98665 91410 98870
rect 91578 98665 91778 98870
rect 91946 98665 92146 98870
rect 92314 98665 96490 98870
rect 296 856 96490 98665
rect 296 800 24250 856
rect 24418 800 72918 856
rect 73086 800 96490 856
<< metal3 >>
rect 96577 96024 97377 96144
rect 96577 93032 97377 93152
rect 0 91128 800 91248
rect 0 90312 800 90432
rect 96577 90040 97377 90160
rect 0 89496 800 89616
rect 0 88680 800 88800
rect 0 87864 800 87984
rect 0 87048 800 87168
rect 96577 87048 97377 87168
rect 0 86232 800 86352
rect 0 85416 800 85536
rect 0 84600 800 84720
rect 96577 84056 97377 84176
rect 0 83784 800 83904
rect 0 82968 800 83088
rect 0 82152 800 82272
rect 0 81336 800 81456
rect 96577 81064 97377 81184
rect 0 80520 800 80640
rect 0 79704 800 79824
rect 0 78888 800 79008
rect 0 78072 800 78192
rect 96577 78072 97377 78192
rect 0 77256 800 77376
rect 0 76440 800 76560
rect 0 75624 800 75744
rect 96577 75080 97377 75200
rect 0 74808 800 74928
rect 0 73992 800 74112
rect 0 73176 800 73296
rect 0 72360 800 72480
rect 96577 72088 97377 72208
rect 0 71544 800 71664
rect 0 70728 800 70848
rect 0 69912 800 70032
rect 0 69096 800 69216
rect 96577 69096 97377 69216
rect 0 68280 800 68400
rect 0 67464 800 67584
rect 0 66648 800 66768
rect 96577 66104 97377 66224
rect 0 65832 800 65952
rect 0 65016 800 65136
rect 0 64200 800 64320
rect 0 63384 800 63504
rect 96577 63112 97377 63232
rect 0 62568 800 62688
rect 0 61752 800 61872
rect 0 60936 800 61056
rect 0 60120 800 60240
rect 96577 60120 97377 60240
rect 0 59304 800 59424
rect 0 58488 800 58608
rect 0 57672 800 57792
rect 96577 57128 97377 57248
rect 0 56856 800 56976
rect 0 56040 800 56160
rect 0 55224 800 55344
rect 0 54408 800 54528
rect 96577 54136 97377 54256
rect 0 53592 800 53712
rect 0 52776 800 52896
rect 0 51960 800 52080
rect 0 51144 800 51264
rect 96577 51144 97377 51264
rect 0 50328 800 50448
rect 0 49512 800 49632
rect 0 48696 800 48816
rect 96577 48152 97377 48272
rect 0 47880 800 48000
rect 0 47064 800 47184
rect 0 46248 800 46368
rect 0 45432 800 45552
rect 96577 45160 97377 45280
rect 0 44616 800 44736
rect 0 43800 800 43920
rect 0 42984 800 43104
rect 0 42168 800 42288
rect 96577 42168 97377 42288
rect 0 41352 800 41472
rect 0 40536 800 40656
rect 0 39720 800 39840
rect 96577 39176 97377 39296
rect 0 38904 800 39024
rect 0 38088 800 38208
rect 0 37272 800 37392
rect 0 36456 800 36576
rect 96577 36184 97377 36304
rect 0 35640 800 35760
rect 0 34824 800 34944
rect 0 34008 800 34128
rect 0 33192 800 33312
rect 96577 33192 97377 33312
rect 0 32376 800 32496
rect 0 31560 800 31680
rect 0 30744 800 30864
rect 96577 30200 97377 30320
rect 0 29928 800 30048
rect 0 29112 800 29232
rect 0 28296 800 28416
rect 0 27480 800 27600
rect 96577 27208 97377 27328
rect 0 26664 800 26784
rect 0 25848 800 25968
rect 0 25032 800 25152
rect 0 24216 800 24336
rect 96577 24216 97377 24336
rect 0 23400 800 23520
rect 0 22584 800 22704
rect 0 21768 800 21888
rect 96577 21224 97377 21344
rect 0 20952 800 21072
rect 0 20136 800 20256
rect 0 19320 800 19440
rect 0 18504 800 18624
rect 96577 18232 97377 18352
rect 0 17688 800 17808
rect 0 16872 800 16992
rect 0 16056 800 16176
rect 0 15240 800 15360
rect 96577 15240 97377 15360
rect 0 14424 800 14544
rect 0 13608 800 13728
rect 0 12792 800 12912
rect 96577 12248 97377 12368
rect 0 11976 800 12096
rect 0 11160 800 11280
rect 0 10344 800 10464
rect 0 9528 800 9648
rect 96577 9256 97377 9376
rect 0 8712 800 8832
rect 0 7896 800 8016
rect 96577 6264 97377 6384
rect 96577 3272 97377 3392
<< obsm3 >>
rect 54 96224 96577 98700
rect 54 95944 96497 96224
rect 54 93232 96577 95944
rect 54 92952 96497 93232
rect 54 91328 96577 92952
rect 880 91048 96577 91328
rect 54 90512 96577 91048
rect 880 90240 96577 90512
rect 880 90232 96497 90240
rect 54 89960 96497 90232
rect 54 89696 96577 89960
rect 880 89416 96577 89696
rect 54 88880 96577 89416
rect 880 88600 96577 88880
rect 54 88064 96577 88600
rect 880 87784 96577 88064
rect 54 87248 96577 87784
rect 880 86968 96497 87248
rect 54 86432 96577 86968
rect 880 86152 96577 86432
rect 54 85616 96577 86152
rect 880 85336 96577 85616
rect 54 84800 96577 85336
rect 880 84520 96577 84800
rect 54 84256 96577 84520
rect 54 83984 96497 84256
rect 880 83976 96497 83984
rect 880 83704 96577 83976
rect 54 83168 96577 83704
rect 880 82888 96577 83168
rect 54 82352 96577 82888
rect 880 82072 96577 82352
rect 54 81536 96577 82072
rect 880 81264 96577 81536
rect 880 81256 96497 81264
rect 54 80984 96497 81256
rect 54 80720 96577 80984
rect 880 80440 96577 80720
rect 54 79904 96577 80440
rect 880 79624 96577 79904
rect 54 79088 96577 79624
rect 880 78808 96577 79088
rect 54 78272 96577 78808
rect 880 77992 96497 78272
rect 54 77456 96577 77992
rect 880 77176 96577 77456
rect 54 76640 96577 77176
rect 880 76360 96577 76640
rect 54 75824 96577 76360
rect 880 75544 96577 75824
rect 54 75280 96577 75544
rect 54 75008 96497 75280
rect 880 75000 96497 75008
rect 880 74728 96577 75000
rect 54 74192 96577 74728
rect 880 73912 96577 74192
rect 54 73376 96577 73912
rect 880 73096 96577 73376
rect 54 72560 96577 73096
rect 880 72288 96577 72560
rect 880 72280 96497 72288
rect 54 72008 96497 72280
rect 54 71744 96577 72008
rect 880 71464 96577 71744
rect 54 70928 96577 71464
rect 880 70648 96577 70928
rect 54 70112 96577 70648
rect 880 69832 96577 70112
rect 54 69296 96577 69832
rect 880 69016 96497 69296
rect 54 68480 96577 69016
rect 880 68200 96577 68480
rect 54 67664 96577 68200
rect 880 67384 96577 67664
rect 54 66848 96577 67384
rect 880 66568 96577 66848
rect 54 66304 96577 66568
rect 54 66032 96497 66304
rect 880 66024 96497 66032
rect 880 65752 96577 66024
rect 54 65216 96577 65752
rect 880 64936 96577 65216
rect 54 64400 96577 64936
rect 880 64120 96577 64400
rect 54 63584 96577 64120
rect 880 63312 96577 63584
rect 880 63304 96497 63312
rect 54 63032 96497 63304
rect 54 62768 96577 63032
rect 880 62488 96577 62768
rect 54 61952 96577 62488
rect 880 61672 96577 61952
rect 54 61136 96577 61672
rect 880 60856 96577 61136
rect 54 60320 96577 60856
rect 880 60040 96497 60320
rect 54 59504 96577 60040
rect 880 59224 96577 59504
rect 54 58688 96577 59224
rect 880 58408 96577 58688
rect 54 57872 96577 58408
rect 880 57592 96577 57872
rect 54 57328 96577 57592
rect 54 57056 96497 57328
rect 880 57048 96497 57056
rect 880 56776 96577 57048
rect 54 56240 96577 56776
rect 880 55960 96577 56240
rect 54 55424 96577 55960
rect 880 55144 96577 55424
rect 54 54608 96577 55144
rect 880 54336 96577 54608
rect 880 54328 96497 54336
rect 54 54056 96497 54328
rect 54 53792 96577 54056
rect 880 53512 96577 53792
rect 54 52976 96577 53512
rect 880 52696 96577 52976
rect 54 52160 96577 52696
rect 880 51880 96577 52160
rect 54 51344 96577 51880
rect 880 51064 96497 51344
rect 54 50528 96577 51064
rect 880 50248 96577 50528
rect 54 49712 96577 50248
rect 880 49432 96577 49712
rect 54 48896 96577 49432
rect 880 48616 96577 48896
rect 54 48352 96577 48616
rect 54 48080 96497 48352
rect 880 48072 96497 48080
rect 880 47800 96577 48072
rect 54 47264 96577 47800
rect 880 46984 96577 47264
rect 54 46448 96577 46984
rect 880 46168 96577 46448
rect 54 45632 96577 46168
rect 880 45360 96577 45632
rect 880 45352 96497 45360
rect 54 45080 96497 45352
rect 54 44816 96577 45080
rect 880 44536 96577 44816
rect 54 44000 96577 44536
rect 880 43720 96577 44000
rect 54 43184 96577 43720
rect 880 42904 96577 43184
rect 54 42368 96577 42904
rect 880 42088 96497 42368
rect 54 41552 96577 42088
rect 880 41272 96577 41552
rect 54 40736 96577 41272
rect 880 40456 96577 40736
rect 54 39920 96577 40456
rect 880 39640 96577 39920
rect 54 39376 96577 39640
rect 54 39104 96497 39376
rect 880 39096 96497 39104
rect 880 38824 96577 39096
rect 54 38288 96577 38824
rect 880 38008 96577 38288
rect 54 37472 96577 38008
rect 880 37192 96577 37472
rect 54 36656 96577 37192
rect 880 36384 96577 36656
rect 880 36376 96497 36384
rect 54 36104 96497 36376
rect 54 35840 96577 36104
rect 880 35560 96577 35840
rect 54 35024 96577 35560
rect 880 34744 96577 35024
rect 54 34208 96577 34744
rect 880 33928 96577 34208
rect 54 33392 96577 33928
rect 880 33112 96497 33392
rect 54 32576 96577 33112
rect 880 32296 96577 32576
rect 54 31760 96577 32296
rect 880 31480 96577 31760
rect 54 30944 96577 31480
rect 880 30664 96577 30944
rect 54 30400 96577 30664
rect 54 30128 96497 30400
rect 880 30120 96497 30128
rect 880 29848 96577 30120
rect 54 29312 96577 29848
rect 880 29032 96577 29312
rect 54 28496 96577 29032
rect 880 28216 96577 28496
rect 54 27680 96577 28216
rect 880 27408 96577 27680
rect 880 27400 96497 27408
rect 54 27128 96497 27400
rect 54 26864 96577 27128
rect 880 26584 96577 26864
rect 54 26048 96577 26584
rect 880 25768 96577 26048
rect 54 25232 96577 25768
rect 880 24952 96577 25232
rect 54 24416 96577 24952
rect 880 24136 96497 24416
rect 54 23600 96577 24136
rect 880 23320 96577 23600
rect 54 22784 96577 23320
rect 880 22504 96577 22784
rect 54 21968 96577 22504
rect 880 21688 96577 21968
rect 54 21424 96577 21688
rect 54 21152 96497 21424
rect 880 21144 96497 21152
rect 880 20872 96577 21144
rect 54 20336 96577 20872
rect 880 20056 96577 20336
rect 54 19520 96577 20056
rect 880 19240 96577 19520
rect 54 18704 96577 19240
rect 880 18432 96577 18704
rect 880 18424 96497 18432
rect 54 18152 96497 18424
rect 54 17888 96577 18152
rect 880 17608 96577 17888
rect 54 17072 96577 17608
rect 880 16792 96577 17072
rect 54 16256 96577 16792
rect 880 15976 96577 16256
rect 54 15440 96577 15976
rect 880 15160 96497 15440
rect 54 14624 96577 15160
rect 880 14344 96577 14624
rect 54 13808 96577 14344
rect 880 13528 96577 13808
rect 54 12992 96577 13528
rect 880 12712 96577 12992
rect 54 12448 96577 12712
rect 54 12176 96497 12448
rect 880 12168 96497 12176
rect 880 11896 96577 12168
rect 54 11360 96577 11896
rect 880 11080 96577 11360
rect 54 10544 96577 11080
rect 880 10264 96577 10544
rect 54 9728 96577 10264
rect 880 9456 96577 9728
rect 880 9448 96497 9456
rect 54 9176 96497 9448
rect 54 8912 96577 9176
rect 880 8632 96577 8912
rect 54 8096 96577 8632
rect 880 7816 96577 8096
rect 54 6464 96577 7816
rect 54 6184 96497 6464
rect 54 3472 96577 6184
rect 54 3192 96497 3472
rect 54 2143 96577 3192
<< metal4 >>
rect 4208 2128 4528 96880
rect 19568 2128 19888 96880
rect 34928 2128 35248 96880
rect 50288 2128 50608 96880
rect 65648 2128 65968 96880
rect 81008 2128 81328 96880
<< obsm4 >>
rect 59 96960 92493 98701
rect 59 2619 4128 96960
rect 4608 2619 19488 96960
rect 19968 2619 34848 96960
rect 35328 2619 50208 96960
rect 50688 2619 65568 96960
rect 66048 2619 80928 96960
rect 81408 2619 92493 96960
<< obsm5 >>
rect 300 21260 86548 96380
<< labels >>
rlabel metal4 s 19568 2128 19888 96880 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 96880 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 96880 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 96880 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 96880 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 96880 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 72974 0 73030 800 6 clk
port 3 nsew signal input
rlabel metal2 s 31482 98721 31538 99521 6 cpi_insn[0]
port 4 nsew signal output
rlabel metal2 s 35162 98721 35218 99521 6 cpi_insn[10]
port 5 nsew signal output
rlabel metal2 s 35530 98721 35586 99521 6 cpi_insn[11]
port 6 nsew signal output
rlabel metal2 s 35898 98721 35954 99521 6 cpi_insn[12]
port 7 nsew signal output
rlabel metal2 s 36266 98721 36322 99521 6 cpi_insn[13]
port 8 nsew signal output
rlabel metal2 s 36634 98721 36690 99521 6 cpi_insn[14]
port 9 nsew signal output
rlabel metal2 s 37002 98721 37058 99521 6 cpi_insn[15]
port 10 nsew signal output
rlabel metal2 s 37370 98721 37426 99521 6 cpi_insn[16]
port 11 nsew signal output
rlabel metal2 s 37738 98721 37794 99521 6 cpi_insn[17]
port 12 nsew signal output
rlabel metal2 s 38106 98721 38162 99521 6 cpi_insn[18]
port 13 nsew signal output
rlabel metal2 s 38474 98721 38530 99521 6 cpi_insn[19]
port 14 nsew signal output
rlabel metal2 s 31850 98721 31906 99521 6 cpi_insn[1]
port 15 nsew signal output
rlabel metal2 s 38842 98721 38898 99521 6 cpi_insn[20]
port 16 nsew signal output
rlabel metal2 s 39210 98721 39266 99521 6 cpi_insn[21]
port 17 nsew signal output
rlabel metal2 s 39578 98721 39634 99521 6 cpi_insn[22]
port 18 nsew signal output
rlabel metal2 s 39946 98721 40002 99521 6 cpi_insn[23]
port 19 nsew signal output
rlabel metal2 s 40314 98721 40370 99521 6 cpi_insn[24]
port 20 nsew signal output
rlabel metal2 s 40682 98721 40738 99521 6 cpi_insn[25]
port 21 nsew signal output
rlabel metal2 s 41050 98721 41106 99521 6 cpi_insn[26]
port 22 nsew signal output
rlabel metal2 s 41418 98721 41474 99521 6 cpi_insn[27]
port 23 nsew signal output
rlabel metal2 s 41786 98721 41842 99521 6 cpi_insn[28]
port 24 nsew signal output
rlabel metal2 s 42154 98721 42210 99521 6 cpi_insn[29]
port 25 nsew signal output
rlabel metal2 s 32218 98721 32274 99521 6 cpi_insn[2]
port 26 nsew signal output
rlabel metal2 s 42522 98721 42578 99521 6 cpi_insn[30]
port 27 nsew signal output
rlabel metal2 s 42890 98721 42946 99521 6 cpi_insn[31]
port 28 nsew signal output
rlabel metal2 s 32586 98721 32642 99521 6 cpi_insn[3]
port 29 nsew signal output
rlabel metal2 s 32954 98721 33010 99521 6 cpi_insn[4]
port 30 nsew signal output
rlabel metal2 s 33322 98721 33378 99521 6 cpi_insn[5]
port 31 nsew signal output
rlabel metal2 s 33690 98721 33746 99521 6 cpi_insn[6]
port 32 nsew signal output
rlabel metal2 s 34058 98721 34114 99521 6 cpi_insn[7]
port 33 nsew signal output
rlabel metal2 s 34426 98721 34482 99521 6 cpi_insn[8]
port 34 nsew signal output
rlabel metal2 s 34794 98721 34850 99521 6 cpi_insn[9]
port 35 nsew signal output
rlabel metal2 s 43258 98721 43314 99521 6 cpi_rs1[0]
port 36 nsew signal output
rlabel metal2 s 46938 98721 46994 99521 6 cpi_rs1[10]
port 37 nsew signal output
rlabel metal2 s 47306 98721 47362 99521 6 cpi_rs1[11]
port 38 nsew signal output
rlabel metal2 s 47674 98721 47730 99521 6 cpi_rs1[12]
port 39 nsew signal output
rlabel metal2 s 48042 98721 48098 99521 6 cpi_rs1[13]
port 40 nsew signal output
rlabel metal2 s 48410 98721 48466 99521 6 cpi_rs1[14]
port 41 nsew signal output
rlabel metal2 s 48778 98721 48834 99521 6 cpi_rs1[15]
port 42 nsew signal output
rlabel metal2 s 49146 98721 49202 99521 6 cpi_rs1[16]
port 43 nsew signal output
rlabel metal2 s 49514 98721 49570 99521 6 cpi_rs1[17]
port 44 nsew signal output
rlabel metal2 s 49882 98721 49938 99521 6 cpi_rs1[18]
port 45 nsew signal output
rlabel metal2 s 50250 98721 50306 99521 6 cpi_rs1[19]
port 46 nsew signal output
rlabel metal2 s 43626 98721 43682 99521 6 cpi_rs1[1]
port 47 nsew signal output
rlabel metal2 s 50618 98721 50674 99521 6 cpi_rs1[20]
port 48 nsew signal output
rlabel metal2 s 50986 98721 51042 99521 6 cpi_rs1[21]
port 49 nsew signal output
rlabel metal2 s 51354 98721 51410 99521 6 cpi_rs1[22]
port 50 nsew signal output
rlabel metal2 s 51722 98721 51778 99521 6 cpi_rs1[23]
port 51 nsew signal output
rlabel metal2 s 52090 98721 52146 99521 6 cpi_rs1[24]
port 52 nsew signal output
rlabel metal2 s 52458 98721 52514 99521 6 cpi_rs1[25]
port 53 nsew signal output
rlabel metal2 s 52826 98721 52882 99521 6 cpi_rs1[26]
port 54 nsew signal output
rlabel metal2 s 53194 98721 53250 99521 6 cpi_rs1[27]
port 55 nsew signal output
rlabel metal2 s 53562 98721 53618 99521 6 cpi_rs1[28]
port 56 nsew signal output
rlabel metal2 s 53930 98721 53986 99521 6 cpi_rs1[29]
port 57 nsew signal output
rlabel metal2 s 43994 98721 44050 99521 6 cpi_rs1[2]
port 58 nsew signal output
rlabel metal2 s 54298 98721 54354 99521 6 cpi_rs1[30]
port 59 nsew signal output
rlabel metal2 s 54666 98721 54722 99521 6 cpi_rs1[31]
port 60 nsew signal output
rlabel metal2 s 44362 98721 44418 99521 6 cpi_rs1[3]
port 61 nsew signal output
rlabel metal2 s 44730 98721 44786 99521 6 cpi_rs1[4]
port 62 nsew signal output
rlabel metal2 s 45098 98721 45154 99521 6 cpi_rs1[5]
port 63 nsew signal output
rlabel metal2 s 45466 98721 45522 99521 6 cpi_rs1[6]
port 64 nsew signal output
rlabel metal2 s 45834 98721 45890 99521 6 cpi_rs1[7]
port 65 nsew signal output
rlabel metal2 s 46202 98721 46258 99521 6 cpi_rs1[8]
port 66 nsew signal output
rlabel metal2 s 46570 98721 46626 99521 6 cpi_rs1[9]
port 67 nsew signal output
rlabel metal2 s 55034 98721 55090 99521 6 cpi_rs2[0]
port 68 nsew signal output
rlabel metal2 s 58714 98721 58770 99521 6 cpi_rs2[10]
port 69 nsew signal output
rlabel metal2 s 59082 98721 59138 99521 6 cpi_rs2[11]
port 70 nsew signal output
rlabel metal2 s 59450 98721 59506 99521 6 cpi_rs2[12]
port 71 nsew signal output
rlabel metal2 s 59818 98721 59874 99521 6 cpi_rs2[13]
port 72 nsew signal output
rlabel metal2 s 60186 98721 60242 99521 6 cpi_rs2[14]
port 73 nsew signal output
rlabel metal2 s 60554 98721 60610 99521 6 cpi_rs2[15]
port 74 nsew signal output
rlabel metal2 s 60922 98721 60978 99521 6 cpi_rs2[16]
port 75 nsew signal output
rlabel metal2 s 61290 98721 61346 99521 6 cpi_rs2[17]
port 76 nsew signal output
rlabel metal2 s 61658 98721 61714 99521 6 cpi_rs2[18]
port 77 nsew signal output
rlabel metal2 s 62026 98721 62082 99521 6 cpi_rs2[19]
port 78 nsew signal output
rlabel metal2 s 55402 98721 55458 99521 6 cpi_rs2[1]
port 79 nsew signal output
rlabel metal2 s 62394 98721 62450 99521 6 cpi_rs2[20]
port 80 nsew signal output
rlabel metal2 s 62762 98721 62818 99521 6 cpi_rs2[21]
port 81 nsew signal output
rlabel metal2 s 63130 98721 63186 99521 6 cpi_rs2[22]
port 82 nsew signal output
rlabel metal2 s 63498 98721 63554 99521 6 cpi_rs2[23]
port 83 nsew signal output
rlabel metal2 s 63866 98721 63922 99521 6 cpi_rs2[24]
port 84 nsew signal output
rlabel metal2 s 64234 98721 64290 99521 6 cpi_rs2[25]
port 85 nsew signal output
rlabel metal2 s 64602 98721 64658 99521 6 cpi_rs2[26]
port 86 nsew signal output
rlabel metal2 s 64970 98721 65026 99521 6 cpi_rs2[27]
port 87 nsew signal output
rlabel metal2 s 65338 98721 65394 99521 6 cpi_rs2[28]
port 88 nsew signal output
rlabel metal2 s 65706 98721 65762 99521 6 cpi_rs2[29]
port 89 nsew signal output
rlabel metal2 s 55770 98721 55826 99521 6 cpi_rs2[2]
port 90 nsew signal output
rlabel metal2 s 66074 98721 66130 99521 6 cpi_rs2[30]
port 91 nsew signal output
rlabel metal2 s 66442 98721 66498 99521 6 cpi_rs2[31]
port 92 nsew signal output
rlabel metal2 s 56138 98721 56194 99521 6 cpi_rs2[3]
port 93 nsew signal output
rlabel metal2 s 56506 98721 56562 99521 6 cpi_rs2[4]
port 94 nsew signal output
rlabel metal2 s 56874 98721 56930 99521 6 cpi_rs2[5]
port 95 nsew signal output
rlabel metal2 s 57242 98721 57298 99521 6 cpi_rs2[6]
port 96 nsew signal output
rlabel metal2 s 57610 98721 57666 99521 6 cpi_rs2[7]
port 97 nsew signal output
rlabel metal2 s 57978 98721 58034 99521 6 cpi_rs2[8]
port 98 nsew signal output
rlabel metal2 s 58346 98721 58402 99521 6 cpi_rs2[9]
port 99 nsew signal output
rlabel metal2 s 31114 98721 31170 99521 6 cpi_valid
port 100 nsew signal output
rlabel metal2 s 66810 98721 66866 99521 6 cpi_wait
port 101 nsew signal input
rlabel metal2 s 67178 98721 67234 99521 6 eoi[0]
port 102 nsew signal output
rlabel metal2 s 70858 98721 70914 99521 6 eoi[10]
port 103 nsew signal output
rlabel metal2 s 71226 98721 71282 99521 6 eoi[11]
port 104 nsew signal output
rlabel metal2 s 71594 98721 71650 99521 6 eoi[12]
port 105 nsew signal output
rlabel metal2 s 71962 98721 72018 99521 6 eoi[13]
port 106 nsew signal output
rlabel metal2 s 72330 98721 72386 99521 6 eoi[14]
port 107 nsew signal output
rlabel metal2 s 72698 98721 72754 99521 6 eoi[15]
port 108 nsew signal output
rlabel metal2 s 73066 98721 73122 99521 6 eoi[16]
port 109 nsew signal output
rlabel metal2 s 73434 98721 73490 99521 6 eoi[17]
port 110 nsew signal output
rlabel metal2 s 73802 98721 73858 99521 6 eoi[18]
port 111 nsew signal output
rlabel metal2 s 74170 98721 74226 99521 6 eoi[19]
port 112 nsew signal output
rlabel metal2 s 67546 98721 67602 99521 6 eoi[1]
port 113 nsew signal output
rlabel metal2 s 74538 98721 74594 99521 6 eoi[20]
port 114 nsew signal output
rlabel metal2 s 74906 98721 74962 99521 6 eoi[21]
port 115 nsew signal output
rlabel metal2 s 75274 98721 75330 99521 6 eoi[22]
port 116 nsew signal output
rlabel metal2 s 75642 98721 75698 99521 6 eoi[23]
port 117 nsew signal output
rlabel metal2 s 76010 98721 76066 99521 6 eoi[24]
port 118 nsew signal output
rlabel metal2 s 76378 98721 76434 99521 6 eoi[25]
port 119 nsew signal output
rlabel metal2 s 76746 98721 76802 99521 6 eoi[26]
port 120 nsew signal output
rlabel metal2 s 77114 98721 77170 99521 6 eoi[27]
port 121 nsew signal output
rlabel metal2 s 77482 98721 77538 99521 6 eoi[28]
port 122 nsew signal output
rlabel metal2 s 77850 98721 77906 99521 6 eoi[29]
port 123 nsew signal output
rlabel metal2 s 67914 98721 67970 99521 6 eoi[2]
port 124 nsew signal output
rlabel metal2 s 78218 98721 78274 99521 6 eoi[30]
port 125 nsew signal output
rlabel metal2 s 78586 98721 78642 99521 6 eoi[31]
port 126 nsew signal output
rlabel metal2 s 68282 98721 68338 99521 6 eoi[3]
port 127 nsew signal output
rlabel metal2 s 68650 98721 68706 99521 6 eoi[4]
port 128 nsew signal output
rlabel metal2 s 69018 98721 69074 99521 6 eoi[5]
port 129 nsew signal output
rlabel metal2 s 69386 98721 69442 99521 6 eoi[6]
port 130 nsew signal output
rlabel metal2 s 69754 98721 69810 99521 6 eoi[7]
port 131 nsew signal output
rlabel metal2 s 70122 98721 70178 99521 6 eoi[8]
port 132 nsew signal output
rlabel metal2 s 70490 98721 70546 99521 6 eoi[9]
port 133 nsew signal output
rlabel metal3 s 96577 3272 97377 3392 6 irq[0]
port 134 nsew signal input
rlabel metal3 s 96577 33192 97377 33312 6 irq[10]
port 135 nsew signal input
rlabel metal3 s 96577 36184 97377 36304 6 irq[11]
port 136 nsew signal input
rlabel metal3 s 96577 39176 97377 39296 6 irq[12]
port 137 nsew signal input
rlabel metal3 s 96577 42168 97377 42288 6 irq[13]
port 138 nsew signal input
rlabel metal3 s 96577 45160 97377 45280 6 irq[14]
port 139 nsew signal input
rlabel metal3 s 96577 48152 97377 48272 6 irq[15]
port 140 nsew signal input
rlabel metal3 s 96577 51144 97377 51264 6 irq[16]
port 141 nsew signal input
rlabel metal3 s 96577 54136 97377 54256 6 irq[17]
port 142 nsew signal input
rlabel metal3 s 96577 57128 97377 57248 6 irq[18]
port 143 nsew signal input
rlabel metal3 s 96577 60120 97377 60240 6 irq[19]
port 144 nsew signal input
rlabel metal3 s 96577 6264 97377 6384 6 irq[1]
port 145 nsew signal input
rlabel metal3 s 96577 63112 97377 63232 6 irq[20]
port 146 nsew signal input
rlabel metal3 s 96577 66104 97377 66224 6 irq[21]
port 147 nsew signal input
rlabel metal3 s 96577 69096 97377 69216 6 irq[22]
port 148 nsew signal input
rlabel metal3 s 96577 72088 97377 72208 6 irq[23]
port 149 nsew signal input
rlabel metal3 s 96577 75080 97377 75200 6 irq[24]
port 150 nsew signal input
rlabel metal3 s 96577 78072 97377 78192 6 irq[25]
port 151 nsew signal input
rlabel metal3 s 96577 81064 97377 81184 6 irq[26]
port 152 nsew signal input
rlabel metal3 s 96577 84056 97377 84176 6 irq[27]
port 153 nsew signal input
rlabel metal3 s 96577 87048 97377 87168 6 irq[28]
port 154 nsew signal input
rlabel metal3 s 96577 90040 97377 90160 6 irq[29]
port 155 nsew signal input
rlabel metal3 s 96577 9256 97377 9376 6 irq[2]
port 156 nsew signal input
rlabel metal3 s 96577 93032 97377 93152 6 irq[30]
port 157 nsew signal input
rlabel metal3 s 96577 96024 97377 96144 6 irq[31]
port 158 nsew signal input
rlabel metal3 s 96577 12248 97377 12368 6 irq[3]
port 159 nsew signal input
rlabel metal3 s 96577 15240 97377 15360 6 irq[4]
port 160 nsew signal input
rlabel metal3 s 96577 18232 97377 18352 6 irq[5]
port 161 nsew signal input
rlabel metal3 s 96577 21224 97377 21344 6 irq[6]
port 162 nsew signal input
rlabel metal3 s 96577 24216 97377 24336 6 irq[7]
port 163 nsew signal input
rlabel metal3 s 96577 27208 97377 27328 6 irq[8]
port 164 nsew signal input
rlabel metal3 s 96577 30200 97377 30320 6 irq[9]
port 165 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 mem_addr[0]
port 166 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 mem_addr[10]
port 167 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 mem_addr[11]
port 168 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 mem_addr[12]
port 169 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 mem_addr[13]
port 170 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 mem_addr[14]
port 171 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 mem_addr[15]
port 172 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 mem_addr[16]
port 173 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 mem_addr[17]
port 174 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 mem_addr[18]
port 175 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 mem_addr[19]
port 176 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 mem_addr[1]
port 177 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 mem_addr[20]
port 178 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 mem_addr[21]
port 179 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 mem_addr[22]
port 180 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 mem_addr[23]
port 181 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 mem_addr[24]
port 182 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 mem_addr[25]
port 183 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 mem_addr[26]
port 184 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 mem_addr[27]
port 185 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 mem_addr[28]
port 186 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 mem_addr[29]
port 187 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 mem_addr[2]
port 188 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 mem_addr[30]
port 189 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 mem_addr[31]
port 190 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 mem_addr[3]
port 191 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 mem_addr[4]
port 192 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 mem_addr[5]
port 193 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 mem_addr[6]
port 194 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 mem_addr[7]
port 195 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 mem_addr[8]
port 196 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 mem_addr[9]
port 197 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 mem_instr
port 198 nsew signal output
rlabel metal2 s 17866 98721 17922 99521 6 mem_la_addr[0]
port 199 nsew signal output
rlabel metal2 s 21546 98721 21602 99521 6 mem_la_addr[10]
port 200 nsew signal output
rlabel metal2 s 21914 98721 21970 99521 6 mem_la_addr[11]
port 201 nsew signal output
rlabel metal2 s 22282 98721 22338 99521 6 mem_la_addr[12]
port 202 nsew signal output
rlabel metal2 s 22650 98721 22706 99521 6 mem_la_addr[13]
port 203 nsew signal output
rlabel metal2 s 23018 98721 23074 99521 6 mem_la_addr[14]
port 204 nsew signal output
rlabel metal2 s 23386 98721 23442 99521 6 mem_la_addr[15]
port 205 nsew signal output
rlabel metal2 s 23754 98721 23810 99521 6 mem_la_addr[16]
port 206 nsew signal output
rlabel metal2 s 24122 98721 24178 99521 6 mem_la_addr[17]
port 207 nsew signal output
rlabel metal2 s 24490 98721 24546 99521 6 mem_la_addr[18]
port 208 nsew signal output
rlabel metal2 s 24858 98721 24914 99521 6 mem_la_addr[19]
port 209 nsew signal output
rlabel metal2 s 18234 98721 18290 99521 6 mem_la_addr[1]
port 210 nsew signal output
rlabel metal2 s 25226 98721 25282 99521 6 mem_la_addr[20]
port 211 nsew signal output
rlabel metal2 s 25594 98721 25650 99521 6 mem_la_addr[21]
port 212 nsew signal output
rlabel metal2 s 25962 98721 26018 99521 6 mem_la_addr[22]
port 213 nsew signal output
rlabel metal2 s 26330 98721 26386 99521 6 mem_la_addr[23]
port 214 nsew signal output
rlabel metal2 s 26698 98721 26754 99521 6 mem_la_addr[24]
port 215 nsew signal output
rlabel metal2 s 27066 98721 27122 99521 6 mem_la_addr[25]
port 216 nsew signal output
rlabel metal2 s 27434 98721 27490 99521 6 mem_la_addr[26]
port 217 nsew signal output
rlabel metal2 s 27802 98721 27858 99521 6 mem_la_addr[27]
port 218 nsew signal output
rlabel metal2 s 28170 98721 28226 99521 6 mem_la_addr[28]
port 219 nsew signal output
rlabel metal2 s 28538 98721 28594 99521 6 mem_la_addr[29]
port 220 nsew signal output
rlabel metal2 s 18602 98721 18658 99521 6 mem_la_addr[2]
port 221 nsew signal output
rlabel metal2 s 28906 98721 28962 99521 6 mem_la_addr[30]
port 222 nsew signal output
rlabel metal2 s 29274 98721 29330 99521 6 mem_la_addr[31]
port 223 nsew signal output
rlabel metal2 s 18970 98721 19026 99521 6 mem_la_addr[3]
port 224 nsew signal output
rlabel metal2 s 19338 98721 19394 99521 6 mem_la_addr[4]
port 225 nsew signal output
rlabel metal2 s 19706 98721 19762 99521 6 mem_la_addr[5]
port 226 nsew signal output
rlabel metal2 s 20074 98721 20130 99521 6 mem_la_addr[6]
port 227 nsew signal output
rlabel metal2 s 20442 98721 20498 99521 6 mem_la_addr[7]
port 228 nsew signal output
rlabel metal2 s 20810 98721 20866 99521 6 mem_la_addr[8]
port 229 nsew signal output
rlabel metal2 s 21178 98721 21234 99521 6 mem_la_addr[9]
port 230 nsew signal output
rlabel metal2 s 5354 98721 5410 99521 6 mem_la_read
port 231 nsew signal output
rlabel metal2 s 6090 98721 6146 99521 6 mem_la_wdata[0]
port 232 nsew signal output
rlabel metal2 s 9770 98721 9826 99521 6 mem_la_wdata[10]
port 233 nsew signal output
rlabel metal2 s 10138 98721 10194 99521 6 mem_la_wdata[11]
port 234 nsew signal output
rlabel metal2 s 10506 98721 10562 99521 6 mem_la_wdata[12]
port 235 nsew signal output
rlabel metal2 s 10874 98721 10930 99521 6 mem_la_wdata[13]
port 236 nsew signal output
rlabel metal2 s 11242 98721 11298 99521 6 mem_la_wdata[14]
port 237 nsew signal output
rlabel metal2 s 11610 98721 11666 99521 6 mem_la_wdata[15]
port 238 nsew signal output
rlabel metal2 s 11978 98721 12034 99521 6 mem_la_wdata[16]
port 239 nsew signal output
rlabel metal2 s 12346 98721 12402 99521 6 mem_la_wdata[17]
port 240 nsew signal output
rlabel metal2 s 12714 98721 12770 99521 6 mem_la_wdata[18]
port 241 nsew signal output
rlabel metal2 s 13082 98721 13138 99521 6 mem_la_wdata[19]
port 242 nsew signal output
rlabel metal2 s 6458 98721 6514 99521 6 mem_la_wdata[1]
port 243 nsew signal output
rlabel metal2 s 13450 98721 13506 99521 6 mem_la_wdata[20]
port 244 nsew signal output
rlabel metal2 s 13818 98721 13874 99521 6 mem_la_wdata[21]
port 245 nsew signal output
rlabel metal2 s 14186 98721 14242 99521 6 mem_la_wdata[22]
port 246 nsew signal output
rlabel metal2 s 14554 98721 14610 99521 6 mem_la_wdata[23]
port 247 nsew signal output
rlabel metal2 s 14922 98721 14978 99521 6 mem_la_wdata[24]
port 248 nsew signal output
rlabel metal2 s 15290 98721 15346 99521 6 mem_la_wdata[25]
port 249 nsew signal output
rlabel metal2 s 15658 98721 15714 99521 6 mem_la_wdata[26]
port 250 nsew signal output
rlabel metal2 s 16026 98721 16082 99521 6 mem_la_wdata[27]
port 251 nsew signal output
rlabel metal2 s 16394 98721 16450 99521 6 mem_la_wdata[28]
port 252 nsew signal output
rlabel metal2 s 16762 98721 16818 99521 6 mem_la_wdata[29]
port 253 nsew signal output
rlabel metal2 s 6826 98721 6882 99521 6 mem_la_wdata[2]
port 254 nsew signal output
rlabel metal2 s 17130 98721 17186 99521 6 mem_la_wdata[30]
port 255 nsew signal output
rlabel metal2 s 17498 98721 17554 99521 6 mem_la_wdata[31]
port 256 nsew signal output
rlabel metal2 s 7194 98721 7250 99521 6 mem_la_wdata[3]
port 257 nsew signal output
rlabel metal2 s 7562 98721 7618 99521 6 mem_la_wdata[4]
port 258 nsew signal output
rlabel metal2 s 7930 98721 7986 99521 6 mem_la_wdata[5]
port 259 nsew signal output
rlabel metal2 s 8298 98721 8354 99521 6 mem_la_wdata[6]
port 260 nsew signal output
rlabel metal2 s 8666 98721 8722 99521 6 mem_la_wdata[7]
port 261 nsew signal output
rlabel metal2 s 9034 98721 9090 99521 6 mem_la_wdata[8]
port 262 nsew signal output
rlabel metal2 s 9402 98721 9458 99521 6 mem_la_wdata[9]
port 263 nsew signal output
rlabel metal2 s 5722 98721 5778 99521 6 mem_la_write
port 264 nsew signal output
rlabel metal2 s 29642 98721 29698 99521 6 mem_la_wstrb[0]
port 265 nsew signal output
rlabel metal2 s 30010 98721 30066 99521 6 mem_la_wstrb[1]
port 266 nsew signal output
rlabel metal2 s 30378 98721 30434 99521 6 mem_la_wstrb[2]
port 267 nsew signal output
rlabel metal2 s 30746 98721 30802 99521 6 mem_la_wstrb[3]
port 268 nsew signal output
rlabel metal3 s 0 65832 800 65952 6 mem_rdata[0]
port 269 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 mem_rdata[10]
port 270 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 mem_rdata[11]
port 271 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 mem_rdata[12]
port 272 nsew signal input
rlabel metal3 s 0 76440 800 76560 6 mem_rdata[13]
port 273 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 mem_rdata[14]
port 274 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 mem_rdata[15]
port 275 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 mem_rdata[16]
port 276 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 mem_rdata[17]
port 277 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 mem_rdata[18]
port 278 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 mem_rdata[19]
port 279 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 mem_rdata[1]
port 280 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 mem_rdata[20]
port 281 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 mem_rdata[21]
port 282 nsew signal input
rlabel metal3 s 0 83784 800 83904 6 mem_rdata[22]
port 283 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 mem_rdata[23]
port 284 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 mem_rdata[24]
port 285 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 mem_rdata[25]
port 286 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 mem_rdata[26]
port 287 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 mem_rdata[27]
port 288 nsew signal input
rlabel metal3 s 0 88680 800 88800 6 mem_rdata[28]
port 289 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 mem_rdata[29]
port 290 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 mem_rdata[2]
port 291 nsew signal input
rlabel metal3 s 0 90312 800 90432 6 mem_rdata[30]
port 292 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 mem_rdata[31]
port 293 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 mem_rdata[3]
port 294 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 mem_rdata[4]
port 295 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 mem_rdata[5]
port 296 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 mem_rdata[6]
port 297 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 mem_rdata[7]
port 298 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 mem_rdata[8]
port 299 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 mem_rdata[9]
port 300 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 mem_ready
port 301 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 mem_valid
port 302 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 mem_wdata[0]
port 303 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 mem_wdata[10]
port 304 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 mem_wdata[11]
port 305 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 mem_wdata[12]
port 306 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 mem_wdata[13]
port 307 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 mem_wdata[14]
port 308 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 mem_wdata[15]
port 309 nsew signal output
rlabel metal3 s 0 49512 800 49632 6 mem_wdata[16]
port 310 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 mem_wdata[17]
port 311 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 mem_wdata[18]
port 312 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 mem_wdata[19]
port 313 nsew signal output
rlabel metal3 s 0 37272 800 37392 6 mem_wdata[1]
port 314 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 mem_wdata[20]
port 315 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 mem_wdata[21]
port 316 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 mem_wdata[22]
port 317 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 mem_wdata[23]
port 318 nsew signal output
rlabel metal3 s 0 56040 800 56160 6 mem_wdata[24]
port 319 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 mem_wdata[25]
port 320 nsew signal output
rlabel metal3 s 0 57672 800 57792 6 mem_wdata[26]
port 321 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 mem_wdata[27]
port 322 nsew signal output
rlabel metal3 s 0 59304 800 59424 6 mem_wdata[28]
port 323 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 mem_wdata[29]
port 324 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 mem_wdata[2]
port 325 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 mem_wdata[30]
port 326 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 mem_wdata[31]
port 327 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 mem_wdata[3]
port 328 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 mem_wdata[4]
port 329 nsew signal output
rlabel metal3 s 0 40536 800 40656 6 mem_wdata[5]
port 330 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 mem_wdata[6]
port 331 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 mem_wdata[7]
port 332 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 mem_wdata[8]
port 333 nsew signal output
rlabel metal3 s 0 43800 800 43920 6 mem_wdata[9]
port 334 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 mem_wstrb[0]
port 335 nsew signal output
rlabel metal3 s 0 63384 800 63504 6 mem_wstrb[1]
port 336 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 mem_wstrb[2]
port 337 nsew signal output
rlabel metal3 s 0 65016 800 65136 6 mem_wstrb[3]
port 338 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 resetn
port 339 nsew signal input
rlabel metal2 s 79322 98721 79378 99521 6 trace_data[0]
port 340 nsew signal output
rlabel metal2 s 83002 98721 83058 99521 6 trace_data[10]
port 341 nsew signal output
rlabel metal2 s 83370 98721 83426 99521 6 trace_data[11]
port 342 nsew signal output
rlabel metal2 s 83738 98721 83794 99521 6 trace_data[12]
port 343 nsew signal output
rlabel metal2 s 84106 98721 84162 99521 6 trace_data[13]
port 344 nsew signal output
rlabel metal2 s 84474 98721 84530 99521 6 trace_data[14]
port 345 nsew signal output
rlabel metal2 s 84842 98721 84898 99521 6 trace_data[15]
port 346 nsew signal output
rlabel metal2 s 85210 98721 85266 99521 6 trace_data[16]
port 347 nsew signal output
rlabel metal2 s 85578 98721 85634 99521 6 trace_data[17]
port 348 nsew signal output
rlabel metal2 s 85946 98721 86002 99521 6 trace_data[18]
port 349 nsew signal output
rlabel metal2 s 86314 98721 86370 99521 6 trace_data[19]
port 350 nsew signal output
rlabel metal2 s 79690 98721 79746 99521 6 trace_data[1]
port 351 nsew signal output
rlabel metal2 s 86682 98721 86738 99521 6 trace_data[20]
port 352 nsew signal output
rlabel metal2 s 87050 98721 87106 99521 6 trace_data[21]
port 353 nsew signal output
rlabel metal2 s 87418 98721 87474 99521 6 trace_data[22]
port 354 nsew signal output
rlabel metal2 s 87786 98721 87842 99521 6 trace_data[23]
port 355 nsew signal output
rlabel metal2 s 88154 98721 88210 99521 6 trace_data[24]
port 356 nsew signal output
rlabel metal2 s 88522 98721 88578 99521 6 trace_data[25]
port 357 nsew signal output
rlabel metal2 s 88890 98721 88946 99521 6 trace_data[26]
port 358 nsew signal output
rlabel metal2 s 89258 98721 89314 99521 6 trace_data[27]
port 359 nsew signal output
rlabel metal2 s 89626 98721 89682 99521 6 trace_data[28]
port 360 nsew signal output
rlabel metal2 s 89994 98721 90050 99521 6 trace_data[29]
port 361 nsew signal output
rlabel metal2 s 80058 98721 80114 99521 6 trace_data[2]
port 362 nsew signal output
rlabel metal2 s 90362 98721 90418 99521 6 trace_data[30]
port 363 nsew signal output
rlabel metal2 s 90730 98721 90786 99521 6 trace_data[31]
port 364 nsew signal output
rlabel metal2 s 91098 98721 91154 99521 6 trace_data[32]
port 365 nsew signal output
rlabel metal2 s 91466 98721 91522 99521 6 trace_data[33]
port 366 nsew signal output
rlabel metal2 s 91834 98721 91890 99521 6 trace_data[34]
port 367 nsew signal output
rlabel metal2 s 92202 98721 92258 99521 6 trace_data[35]
port 368 nsew signal output
rlabel metal2 s 80426 98721 80482 99521 6 trace_data[3]
port 369 nsew signal output
rlabel metal2 s 80794 98721 80850 99521 6 trace_data[4]
port 370 nsew signal output
rlabel metal2 s 81162 98721 81218 99521 6 trace_data[5]
port 371 nsew signal output
rlabel metal2 s 81530 98721 81586 99521 6 trace_data[6]
port 372 nsew signal output
rlabel metal2 s 81898 98721 81954 99521 6 trace_data[7]
port 373 nsew signal output
rlabel metal2 s 82266 98721 82322 99521 6 trace_data[8]
port 374 nsew signal output
rlabel metal2 s 82634 98721 82690 99521 6 trace_data[9]
port 375 nsew signal output
rlabel metal2 s 78954 98721 79010 99521 6 trace_valid
port 376 nsew signal output
rlabel metal2 s 4986 98721 5042 99521 6 trap
port 377 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 97377 99521
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 39544006
string GDS_FILE /openlane/designs/alphacore/runs/RUN_2023.12.03_09.03.48/results/signoff/alphacore.magic.gds
string GDS_START 1198914
<< end >>

