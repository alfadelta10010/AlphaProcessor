magic
tech sky130A
magscale 1 2
timestamp 1701553136
<< nwell >>
rect 1066 175429 175390 175995
rect 1066 174341 175390 174907
rect 1066 173253 175390 173819
rect 1066 172165 175390 172731
rect 1066 171077 175390 171643
rect 1066 169989 175390 170555
rect 1066 168901 175390 169467
rect 1066 167813 175390 168379
rect 1066 166725 175390 167291
rect 1066 165637 175390 166203
rect 1066 164549 175390 165115
rect 1066 163461 175390 164027
rect 1066 162373 175390 162939
rect 1066 161285 175390 161851
rect 1066 160197 175390 160763
rect 1066 159109 175390 159675
rect 1066 158021 175390 158587
rect 1066 156933 175390 157499
rect 1066 155845 175390 156411
rect 1066 154757 175390 155323
rect 1066 153669 175390 154235
rect 1066 152581 175390 153147
rect 1066 151493 175390 152059
rect 1066 150405 175390 150971
rect 1066 149317 175390 149883
rect 1066 148229 175390 148795
rect 1066 147141 175390 147707
rect 1066 146053 175390 146619
rect 1066 144965 175390 145531
rect 1066 143877 175390 144443
rect 1066 142789 175390 143355
rect 1066 141701 175390 142267
rect 1066 140613 175390 141179
rect 1066 139525 175390 140091
rect 1066 138437 175390 139003
rect 1066 137349 175390 137915
rect 1066 136261 175390 136827
rect 1066 135173 175390 135739
rect 1066 134085 175390 134651
rect 1066 132997 175390 133563
rect 1066 131909 175390 132475
rect 1066 130821 175390 131387
rect 1066 129733 175390 130299
rect 1066 128645 175390 129211
rect 1066 127557 175390 128123
rect 1066 126469 175390 127035
rect 1066 125381 175390 125947
rect 1066 124293 175390 124859
rect 1066 123205 175390 123771
rect 1066 122117 175390 122683
rect 1066 121029 175390 121595
rect 1066 119941 175390 120507
rect 1066 118853 175390 119419
rect 1066 117765 175390 118331
rect 1066 116677 175390 117243
rect 1066 115589 175390 116155
rect 1066 114501 175390 115067
rect 1066 113413 175390 113979
rect 1066 112325 175390 112891
rect 1066 111237 175390 111803
rect 1066 110149 175390 110715
rect 1066 109061 175390 109627
rect 1066 107973 175390 108539
rect 1066 106885 175390 107451
rect 1066 105797 175390 106363
rect 1066 104709 175390 105275
rect 1066 103621 175390 104187
rect 1066 102533 175390 103099
rect 1066 101445 175390 102011
rect 1066 100357 175390 100923
rect 1066 99269 175390 99835
rect 1066 98181 175390 98747
rect 1066 97093 175390 97659
rect 1066 96005 175390 96571
rect 1066 94917 175390 95483
rect 1066 93829 175390 94395
rect 1066 92741 175390 93307
rect 1066 91653 175390 92219
rect 1066 90565 175390 91131
rect 1066 89477 175390 90043
rect 1066 88389 175390 88955
rect 1066 87301 175390 87867
rect 1066 86213 175390 86779
rect 1066 85125 175390 85691
rect 1066 84037 175390 84603
rect 1066 82949 175390 83515
rect 1066 81861 175390 82427
rect 1066 80773 175390 81339
rect 1066 79685 175390 80251
rect 1066 78597 175390 79163
rect 1066 77509 175390 78075
rect 1066 76421 175390 76987
rect 1066 75333 175390 75899
rect 1066 74245 175390 74811
rect 1066 73157 175390 73723
rect 1066 72069 175390 72635
rect 1066 70981 175390 71547
rect 1066 69893 175390 70459
rect 1066 68805 175390 69371
rect 1066 67717 175390 68283
rect 1066 66629 175390 67195
rect 1066 65541 175390 66107
rect 1066 64453 175390 65019
rect 1066 63365 175390 63931
rect 1066 62277 175390 62843
rect 1066 61189 175390 61755
rect 1066 60101 175390 60667
rect 1066 59013 175390 59579
rect 1066 57925 175390 58491
rect 1066 56837 175390 57403
rect 1066 55749 175390 56315
rect 1066 54661 175390 55227
rect 1066 53573 175390 54139
rect 1066 52485 175390 53051
rect 1066 51397 175390 51963
rect 1066 50309 175390 50875
rect 1066 49221 175390 49787
rect 1066 48133 175390 48699
rect 1066 47045 175390 47611
rect 1066 45957 175390 46523
rect 1066 44869 175390 45435
rect 1066 43781 175390 44347
rect 1066 42693 175390 43259
rect 1066 41605 175390 42171
rect 1066 40517 175390 41083
rect 1066 39429 175390 39995
rect 1066 38341 175390 38907
rect 1066 37253 175390 37819
rect 1066 36165 175390 36731
rect 1066 35077 175390 35643
rect 1066 33989 175390 34555
rect 1066 32901 175390 33467
rect 1066 31813 175390 32379
rect 1066 30725 175390 31291
rect 1066 29637 175390 30203
rect 1066 28549 175390 29115
rect 1066 27461 175390 28027
rect 1066 26373 175390 26939
rect 1066 25285 175390 25851
rect 1066 24197 175390 24763
rect 1066 23109 175390 23675
rect 1066 22021 175390 22587
rect 1066 20933 175390 21499
rect 1066 19845 175390 20411
rect 1066 18757 175390 19323
rect 1066 17669 175390 18235
rect 1066 16581 175390 17147
rect 1066 15493 175390 16059
rect 1066 14405 175390 14971
rect 1066 13317 175390 13883
rect 1066 12229 175390 12795
rect 1066 11141 175390 11707
rect 1066 10053 175390 10619
rect 1066 8965 175390 9531
rect 1066 7877 175390 8443
rect 1066 6789 175390 7355
rect 1066 5701 175390 6267
rect 1066 4613 175390 5179
rect 1066 3525 175390 4091
rect 1066 2437 175390 3003
<< obsli1 >>
rect 1104 2159 175352 176273
<< obsm1 >>
rect 1104 2128 175614 176384
<< metal2 >>
rect 88154 0 88210 800
<< obsm2 >>
rect 1400 856 175610 176390
rect 1400 800 88098 856
rect 88266 800 175610 856
<< metal3 >>
rect 175715 173816 176515 173936
rect 175715 171912 176515 172032
rect 175715 170008 176515 170128
rect 175715 168104 176515 168224
rect 175715 166200 176515 166320
rect 175715 164296 176515 164416
rect 175715 162392 176515 162512
rect 175715 160488 176515 160608
rect 175715 158584 176515 158704
rect 175715 156680 176515 156800
rect 175715 154776 176515 154896
rect 175715 152872 176515 152992
rect 175715 150968 176515 151088
rect 175715 149064 176515 149184
rect 175715 147160 176515 147280
rect 175715 145256 176515 145376
rect 175715 143352 176515 143472
rect 175715 141448 176515 141568
rect 175715 139544 176515 139664
rect 175715 137640 176515 137760
rect 175715 135736 176515 135856
rect 175715 133832 176515 133952
rect 175715 131928 176515 132048
rect 175715 130024 176515 130144
rect 175715 128120 176515 128240
rect 175715 126216 176515 126336
rect 175715 124312 176515 124432
rect 175715 122408 176515 122528
rect 175715 120504 176515 120624
rect 175715 118600 176515 118720
rect 175715 116696 176515 116816
rect 175715 114792 176515 114912
rect 175715 112888 176515 113008
rect 175715 110984 176515 111104
rect 175715 109080 176515 109200
rect 175715 107176 176515 107296
rect 175715 105272 176515 105392
rect 175715 103368 176515 103488
rect 175715 101464 176515 101584
rect 175715 99560 176515 99680
rect 175715 97656 176515 97776
rect 175715 95752 176515 95872
rect 175715 93848 176515 93968
rect 175715 91944 176515 92064
rect 175715 90040 176515 90160
rect 175715 88136 176515 88256
rect 175715 86232 176515 86352
rect 175715 84328 176515 84448
rect 175715 82424 176515 82544
rect 175715 80520 176515 80640
rect 175715 78616 176515 78736
rect 175715 76712 176515 76832
rect 175715 74808 176515 74928
rect 175715 72904 176515 73024
rect 175715 71000 176515 71120
rect 175715 69096 176515 69216
rect 175715 67192 176515 67312
rect 175715 65288 176515 65408
rect 175715 63384 176515 63504
rect 175715 61480 176515 61600
rect 175715 59576 176515 59696
rect 175715 57672 176515 57792
rect 175715 55768 176515 55888
rect 175715 53864 176515 53984
rect 175715 51960 176515 52080
rect 175715 50056 176515 50176
rect 175715 48152 176515 48272
rect 175715 46248 176515 46368
rect 175715 44344 176515 44464
rect 175715 42440 176515 42560
rect 175715 40536 176515 40656
rect 175715 38632 176515 38752
rect 175715 36728 176515 36848
rect 175715 34824 176515 34944
rect 175715 32920 176515 33040
rect 175715 31016 176515 31136
rect 175715 29112 176515 29232
rect 175715 27208 176515 27328
rect 175715 25304 176515 25424
rect 175715 23400 176515 23520
rect 175715 21496 176515 21616
rect 175715 19592 176515 19712
rect 175715 17688 176515 17808
rect 175715 15784 176515 15904
rect 175715 13880 176515 14000
rect 175715 11976 176515 12096
rect 175715 10072 176515 10192
rect 175715 8168 176515 8288
rect 175715 6264 176515 6384
rect 175715 4360 176515 4480
<< obsm3 >>
rect 4210 174016 175715 176289
rect 4210 173736 175635 174016
rect 4210 172112 175715 173736
rect 4210 171832 175635 172112
rect 4210 170208 175715 171832
rect 4210 169928 175635 170208
rect 4210 168304 175715 169928
rect 4210 168024 175635 168304
rect 4210 166400 175715 168024
rect 4210 166120 175635 166400
rect 4210 164496 175715 166120
rect 4210 164216 175635 164496
rect 4210 162592 175715 164216
rect 4210 162312 175635 162592
rect 4210 160688 175715 162312
rect 4210 160408 175635 160688
rect 4210 158784 175715 160408
rect 4210 158504 175635 158784
rect 4210 156880 175715 158504
rect 4210 156600 175635 156880
rect 4210 154976 175715 156600
rect 4210 154696 175635 154976
rect 4210 153072 175715 154696
rect 4210 152792 175635 153072
rect 4210 151168 175715 152792
rect 4210 150888 175635 151168
rect 4210 149264 175715 150888
rect 4210 148984 175635 149264
rect 4210 147360 175715 148984
rect 4210 147080 175635 147360
rect 4210 145456 175715 147080
rect 4210 145176 175635 145456
rect 4210 143552 175715 145176
rect 4210 143272 175635 143552
rect 4210 141648 175715 143272
rect 4210 141368 175635 141648
rect 4210 139744 175715 141368
rect 4210 139464 175635 139744
rect 4210 137840 175715 139464
rect 4210 137560 175635 137840
rect 4210 135936 175715 137560
rect 4210 135656 175635 135936
rect 4210 134032 175715 135656
rect 4210 133752 175635 134032
rect 4210 132128 175715 133752
rect 4210 131848 175635 132128
rect 4210 130224 175715 131848
rect 4210 129944 175635 130224
rect 4210 128320 175715 129944
rect 4210 128040 175635 128320
rect 4210 126416 175715 128040
rect 4210 126136 175635 126416
rect 4210 124512 175715 126136
rect 4210 124232 175635 124512
rect 4210 122608 175715 124232
rect 4210 122328 175635 122608
rect 4210 120704 175715 122328
rect 4210 120424 175635 120704
rect 4210 118800 175715 120424
rect 4210 118520 175635 118800
rect 4210 116896 175715 118520
rect 4210 116616 175635 116896
rect 4210 114992 175715 116616
rect 4210 114712 175635 114992
rect 4210 113088 175715 114712
rect 4210 112808 175635 113088
rect 4210 111184 175715 112808
rect 4210 110904 175635 111184
rect 4210 109280 175715 110904
rect 4210 109000 175635 109280
rect 4210 107376 175715 109000
rect 4210 107096 175635 107376
rect 4210 105472 175715 107096
rect 4210 105192 175635 105472
rect 4210 103568 175715 105192
rect 4210 103288 175635 103568
rect 4210 101664 175715 103288
rect 4210 101384 175635 101664
rect 4210 99760 175715 101384
rect 4210 99480 175635 99760
rect 4210 97856 175715 99480
rect 4210 97576 175635 97856
rect 4210 95952 175715 97576
rect 4210 95672 175635 95952
rect 4210 94048 175715 95672
rect 4210 93768 175635 94048
rect 4210 92144 175715 93768
rect 4210 91864 175635 92144
rect 4210 90240 175715 91864
rect 4210 89960 175635 90240
rect 4210 88336 175715 89960
rect 4210 88056 175635 88336
rect 4210 86432 175715 88056
rect 4210 86152 175635 86432
rect 4210 84528 175715 86152
rect 4210 84248 175635 84528
rect 4210 82624 175715 84248
rect 4210 82344 175635 82624
rect 4210 80720 175715 82344
rect 4210 80440 175635 80720
rect 4210 78816 175715 80440
rect 4210 78536 175635 78816
rect 4210 76912 175715 78536
rect 4210 76632 175635 76912
rect 4210 75008 175715 76632
rect 4210 74728 175635 75008
rect 4210 73104 175715 74728
rect 4210 72824 175635 73104
rect 4210 71200 175715 72824
rect 4210 70920 175635 71200
rect 4210 69296 175715 70920
rect 4210 69016 175635 69296
rect 4210 67392 175715 69016
rect 4210 67112 175635 67392
rect 4210 65488 175715 67112
rect 4210 65208 175635 65488
rect 4210 63584 175715 65208
rect 4210 63304 175635 63584
rect 4210 61680 175715 63304
rect 4210 61400 175635 61680
rect 4210 59776 175715 61400
rect 4210 59496 175635 59776
rect 4210 57872 175715 59496
rect 4210 57592 175635 57872
rect 4210 55968 175715 57592
rect 4210 55688 175635 55968
rect 4210 54064 175715 55688
rect 4210 53784 175635 54064
rect 4210 52160 175715 53784
rect 4210 51880 175635 52160
rect 4210 50256 175715 51880
rect 4210 49976 175635 50256
rect 4210 48352 175715 49976
rect 4210 48072 175635 48352
rect 4210 46448 175715 48072
rect 4210 46168 175635 46448
rect 4210 44544 175715 46168
rect 4210 44264 175635 44544
rect 4210 42640 175715 44264
rect 4210 42360 175635 42640
rect 4210 40736 175715 42360
rect 4210 40456 175635 40736
rect 4210 38832 175715 40456
rect 4210 38552 175635 38832
rect 4210 36928 175715 38552
rect 4210 36648 175635 36928
rect 4210 35024 175715 36648
rect 4210 34744 175635 35024
rect 4210 33120 175715 34744
rect 4210 32840 175635 33120
rect 4210 31216 175715 32840
rect 4210 30936 175635 31216
rect 4210 29312 175715 30936
rect 4210 29032 175635 29312
rect 4210 27408 175715 29032
rect 4210 27128 175635 27408
rect 4210 25504 175715 27128
rect 4210 25224 175635 25504
rect 4210 23600 175715 25224
rect 4210 23320 175635 23600
rect 4210 21696 175715 23320
rect 4210 21416 175635 21696
rect 4210 19792 175715 21416
rect 4210 19512 175635 19792
rect 4210 17888 175715 19512
rect 4210 17608 175635 17888
rect 4210 15984 175715 17608
rect 4210 15704 175635 15984
rect 4210 14080 175715 15704
rect 4210 13800 175635 14080
rect 4210 12176 175715 13800
rect 4210 11896 175635 12176
rect 4210 10272 175715 11896
rect 4210 9992 175635 10272
rect 4210 8368 175715 9992
rect 4210 8088 175635 8368
rect 4210 6464 175715 8088
rect 4210 6184 175635 6464
rect 4210 4560 175715 6184
rect 4210 4280 175635 4560
rect 4210 2143 175715 4280
<< metal4 >>
rect 4208 2128 4528 176304
rect 19568 2128 19888 176304
rect 34928 2128 35248 176304
rect 50288 2128 50608 176304
rect 65648 2128 65968 176304
rect 81008 2128 81328 176304
rect 96368 2128 96688 176304
rect 111728 2128 112048 176304
rect 127088 2128 127408 176304
rect 142448 2128 142768 176304
rect 157808 2128 158128 176304
rect 173168 2128 173488 176304
<< obsm4 >>
rect 13859 3435 19488 173229
rect 19968 3435 34848 173229
rect 35328 3435 50208 173229
rect 50688 3435 65568 173229
rect 66048 3435 80928 173229
rect 81408 3435 96288 173229
rect 96768 3435 111648 173229
rect 112128 3435 127008 173229
rect 127488 3435 142368 173229
rect 142848 3435 157728 173229
rect 158208 3435 173088 173229
rect 173568 3435 173821 173229
<< obsm5 >>
rect 26060 20580 169532 154860
<< labels >>
rlabel metal4 s 19568 2128 19888 176304 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 176304 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 176304 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 176304 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 176304 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 176304 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 176304 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 176304 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 176304 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 176304 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 176304 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 176304 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 175715 11976 176515 12096 6 addr[0]
port 3 nsew signal input
rlabel metal3 s 175715 31016 176515 31136 6 addr[10]
port 4 nsew signal input
rlabel metal3 s 175715 32920 176515 33040 6 addr[11]
port 5 nsew signal input
rlabel metal3 s 175715 34824 176515 34944 6 addr[12]
port 6 nsew signal input
rlabel metal3 s 175715 36728 176515 36848 6 addr[13]
port 7 nsew signal input
rlabel metal3 s 175715 38632 176515 38752 6 addr[14]
port 8 nsew signal input
rlabel metal3 s 175715 40536 176515 40656 6 addr[15]
port 9 nsew signal input
rlabel metal3 s 175715 42440 176515 42560 6 addr[16]
port 10 nsew signal input
rlabel metal3 s 175715 44344 176515 44464 6 addr[17]
port 11 nsew signal input
rlabel metal3 s 175715 46248 176515 46368 6 addr[18]
port 12 nsew signal input
rlabel metal3 s 175715 48152 176515 48272 6 addr[19]
port 13 nsew signal input
rlabel metal3 s 175715 13880 176515 14000 6 addr[1]
port 14 nsew signal input
rlabel metal3 s 175715 50056 176515 50176 6 addr[20]
port 15 nsew signal input
rlabel metal3 s 175715 51960 176515 52080 6 addr[21]
port 16 nsew signal input
rlabel metal3 s 175715 15784 176515 15904 6 addr[2]
port 17 nsew signal input
rlabel metal3 s 175715 17688 176515 17808 6 addr[3]
port 18 nsew signal input
rlabel metal3 s 175715 19592 176515 19712 6 addr[4]
port 19 nsew signal input
rlabel metal3 s 175715 21496 176515 21616 6 addr[5]
port 20 nsew signal input
rlabel metal3 s 175715 23400 176515 23520 6 addr[6]
port 21 nsew signal input
rlabel metal3 s 175715 25304 176515 25424 6 addr[7]
port 22 nsew signal input
rlabel metal3 s 175715 27208 176515 27328 6 addr[8]
port 23 nsew signal input
rlabel metal3 s 175715 29112 176515 29232 6 addr[9]
port 24 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 clk
port 25 nsew signal input
rlabel metal3 s 175715 114792 176515 114912 6 rdata[0]
port 26 nsew signal output
rlabel metal3 s 175715 133832 176515 133952 6 rdata[10]
port 27 nsew signal output
rlabel metal3 s 175715 135736 176515 135856 6 rdata[11]
port 28 nsew signal output
rlabel metal3 s 175715 137640 176515 137760 6 rdata[12]
port 29 nsew signal output
rlabel metal3 s 175715 139544 176515 139664 6 rdata[13]
port 30 nsew signal output
rlabel metal3 s 175715 141448 176515 141568 6 rdata[14]
port 31 nsew signal output
rlabel metal3 s 175715 143352 176515 143472 6 rdata[15]
port 32 nsew signal output
rlabel metal3 s 175715 145256 176515 145376 6 rdata[16]
port 33 nsew signal output
rlabel metal3 s 175715 147160 176515 147280 6 rdata[17]
port 34 nsew signal output
rlabel metal3 s 175715 149064 176515 149184 6 rdata[18]
port 35 nsew signal output
rlabel metal3 s 175715 150968 176515 151088 6 rdata[19]
port 36 nsew signal output
rlabel metal3 s 175715 116696 176515 116816 6 rdata[1]
port 37 nsew signal output
rlabel metal3 s 175715 152872 176515 152992 6 rdata[20]
port 38 nsew signal output
rlabel metal3 s 175715 154776 176515 154896 6 rdata[21]
port 39 nsew signal output
rlabel metal3 s 175715 156680 176515 156800 6 rdata[22]
port 40 nsew signal output
rlabel metal3 s 175715 158584 176515 158704 6 rdata[23]
port 41 nsew signal output
rlabel metal3 s 175715 160488 176515 160608 6 rdata[24]
port 42 nsew signal output
rlabel metal3 s 175715 162392 176515 162512 6 rdata[25]
port 43 nsew signal output
rlabel metal3 s 175715 164296 176515 164416 6 rdata[26]
port 44 nsew signal output
rlabel metal3 s 175715 166200 176515 166320 6 rdata[27]
port 45 nsew signal output
rlabel metal3 s 175715 168104 176515 168224 6 rdata[28]
port 46 nsew signal output
rlabel metal3 s 175715 170008 176515 170128 6 rdata[29]
port 47 nsew signal output
rlabel metal3 s 175715 118600 176515 118720 6 rdata[2]
port 48 nsew signal output
rlabel metal3 s 175715 171912 176515 172032 6 rdata[30]
port 49 nsew signal output
rlabel metal3 s 175715 173816 176515 173936 6 rdata[31]
port 50 nsew signal output
rlabel metal3 s 175715 120504 176515 120624 6 rdata[3]
port 51 nsew signal output
rlabel metal3 s 175715 122408 176515 122528 6 rdata[4]
port 52 nsew signal output
rlabel metal3 s 175715 124312 176515 124432 6 rdata[5]
port 53 nsew signal output
rlabel metal3 s 175715 126216 176515 126336 6 rdata[6]
port 54 nsew signal output
rlabel metal3 s 175715 128120 176515 128240 6 rdata[7]
port 55 nsew signal output
rlabel metal3 s 175715 130024 176515 130144 6 rdata[8]
port 56 nsew signal output
rlabel metal3 s 175715 131928 176515 132048 6 rdata[9]
port 57 nsew signal output
rlabel metal3 s 175715 53864 176515 53984 6 wdata[0]
port 58 nsew signal input
rlabel metal3 s 175715 72904 176515 73024 6 wdata[10]
port 59 nsew signal input
rlabel metal3 s 175715 74808 176515 74928 6 wdata[11]
port 60 nsew signal input
rlabel metal3 s 175715 76712 176515 76832 6 wdata[12]
port 61 nsew signal input
rlabel metal3 s 175715 78616 176515 78736 6 wdata[13]
port 62 nsew signal input
rlabel metal3 s 175715 80520 176515 80640 6 wdata[14]
port 63 nsew signal input
rlabel metal3 s 175715 82424 176515 82544 6 wdata[15]
port 64 nsew signal input
rlabel metal3 s 175715 84328 176515 84448 6 wdata[16]
port 65 nsew signal input
rlabel metal3 s 175715 86232 176515 86352 6 wdata[17]
port 66 nsew signal input
rlabel metal3 s 175715 88136 176515 88256 6 wdata[18]
port 67 nsew signal input
rlabel metal3 s 175715 90040 176515 90160 6 wdata[19]
port 68 nsew signal input
rlabel metal3 s 175715 55768 176515 55888 6 wdata[1]
port 69 nsew signal input
rlabel metal3 s 175715 91944 176515 92064 6 wdata[20]
port 70 nsew signal input
rlabel metal3 s 175715 93848 176515 93968 6 wdata[21]
port 71 nsew signal input
rlabel metal3 s 175715 95752 176515 95872 6 wdata[22]
port 72 nsew signal input
rlabel metal3 s 175715 97656 176515 97776 6 wdata[23]
port 73 nsew signal input
rlabel metal3 s 175715 99560 176515 99680 6 wdata[24]
port 74 nsew signal input
rlabel metal3 s 175715 101464 176515 101584 6 wdata[25]
port 75 nsew signal input
rlabel metal3 s 175715 103368 176515 103488 6 wdata[26]
port 76 nsew signal input
rlabel metal3 s 175715 105272 176515 105392 6 wdata[27]
port 77 nsew signal input
rlabel metal3 s 175715 107176 176515 107296 6 wdata[28]
port 78 nsew signal input
rlabel metal3 s 175715 109080 176515 109200 6 wdata[29]
port 79 nsew signal input
rlabel metal3 s 175715 57672 176515 57792 6 wdata[2]
port 80 nsew signal input
rlabel metal3 s 175715 110984 176515 111104 6 wdata[30]
port 81 nsew signal input
rlabel metal3 s 175715 112888 176515 113008 6 wdata[31]
port 82 nsew signal input
rlabel metal3 s 175715 59576 176515 59696 6 wdata[3]
port 83 nsew signal input
rlabel metal3 s 175715 61480 176515 61600 6 wdata[4]
port 84 nsew signal input
rlabel metal3 s 175715 63384 176515 63504 6 wdata[5]
port 85 nsew signal input
rlabel metal3 s 175715 65288 176515 65408 6 wdata[6]
port 86 nsew signal input
rlabel metal3 s 175715 67192 176515 67312 6 wdata[7]
port 87 nsew signal input
rlabel metal3 s 175715 69096 176515 69216 6 wdata[8]
port 88 nsew signal input
rlabel metal3 s 175715 71000 176515 71120 6 wdata[9]
port 89 nsew signal input
rlabel metal3 s 175715 4360 176515 4480 6 wen[0]
port 90 nsew signal input
rlabel metal3 s 175715 6264 176515 6384 6 wen[1]
port 91 nsew signal input
rlabel metal3 s 175715 8168 176515 8288 6 wen[2]
port 92 nsew signal input
rlabel metal3 s 175715 10072 176515 10192 6 wen[3]
port 93 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 176515 178659
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 83539458
string GDS_FILE /openlane/designs/alphasoc_mem/runs/RUN_2023.12.02_20.46.33/results/signoff/alphasoc_mem.magic.gds
string GDS_START 338600
<< end >>

