VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alphasoc_mem
  CLASS BLOCK ;
  FOREIGN alphasoc_mem ;
  ORIGIN 0.000 0.000 ;
  SIZE 882.575 BY 893.295 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 881.520 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 881.520 ;
    END
  END VPWR
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 59.880 882.575 60.480 ;
    END
  END addr[0]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 155.080 882.575 155.680 ;
    END
  END addr[10]
  PIN addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 164.600 882.575 165.200 ;
    END
  END addr[11]
  PIN addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 174.120 882.575 174.720 ;
    END
  END addr[12]
  PIN addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 183.640 882.575 184.240 ;
    END
  END addr[13]
  PIN addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 193.160 882.575 193.760 ;
    END
  END addr[14]
  PIN addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 202.680 882.575 203.280 ;
    END
  END addr[15]
  PIN addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 212.200 882.575 212.800 ;
    END
  END addr[16]
  PIN addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 221.720 882.575 222.320 ;
    END
  END addr[17]
  PIN addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 231.240 882.575 231.840 ;
    END
  END addr[18]
  PIN addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 240.760 882.575 241.360 ;
    END
  END addr[19]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 69.400 882.575 70.000 ;
    END
  END addr[1]
  PIN addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 250.280 882.575 250.880 ;
    END
  END addr[20]
  PIN addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 259.800 882.575 260.400 ;
    END
  END addr[21]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 78.920 882.575 79.520 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 88.440 882.575 89.040 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 97.960 882.575 98.560 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 107.480 882.575 108.080 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 117.000 882.575 117.600 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 126.520 882.575 127.120 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 136.040 882.575 136.640 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 878.575 145.560 882.575 146.160 ;
    END
  END addr[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END clk
  PIN rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 573.960 882.575 574.560 ;
    END
  END rdata[0]
  PIN rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 669.160 882.575 669.760 ;
    END
  END rdata[10]
  PIN rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 678.680 882.575 679.280 ;
    END
  END rdata[11]
  PIN rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 688.200 882.575 688.800 ;
    END
  END rdata[12]
  PIN rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 697.720 882.575 698.320 ;
    END
  END rdata[13]
  PIN rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 707.240 882.575 707.840 ;
    END
  END rdata[14]
  PIN rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 716.760 882.575 717.360 ;
    END
  END rdata[15]
  PIN rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 726.280 882.575 726.880 ;
    END
  END rdata[16]
  PIN rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 735.800 882.575 736.400 ;
    END
  END rdata[17]
  PIN rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 745.320 882.575 745.920 ;
    END
  END rdata[18]
  PIN rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 754.840 882.575 755.440 ;
    END
  END rdata[19]
  PIN rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 583.480 882.575 584.080 ;
    END
  END rdata[1]
  PIN rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 764.360 882.575 764.960 ;
    END
  END rdata[20]
  PIN rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 773.880 882.575 774.480 ;
    END
  END rdata[21]
  PIN rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 783.400 882.575 784.000 ;
    END
  END rdata[22]
  PIN rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 792.920 882.575 793.520 ;
    END
  END rdata[23]
  PIN rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 802.440 882.575 803.040 ;
    END
  END rdata[24]
  PIN rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 811.960 882.575 812.560 ;
    END
  END rdata[25]
  PIN rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 821.480 882.575 822.080 ;
    END
  END rdata[26]
  PIN rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 831.000 882.575 831.600 ;
    END
  END rdata[27]
  PIN rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 840.520 882.575 841.120 ;
    END
  END rdata[28]
  PIN rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 850.040 882.575 850.640 ;
    END
  END rdata[29]
  PIN rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 593.000 882.575 593.600 ;
    END
  END rdata[2]
  PIN rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 859.560 882.575 860.160 ;
    END
  END rdata[30]
  PIN rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 869.080 882.575 869.680 ;
    END
  END rdata[31]
  PIN rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 602.520 882.575 603.120 ;
    END
  END rdata[3]
  PIN rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 612.040 882.575 612.640 ;
    END
  END rdata[4]
  PIN rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 621.560 882.575 622.160 ;
    END
  END rdata[5]
  PIN rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 631.080 882.575 631.680 ;
    END
  END rdata[6]
  PIN rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 640.600 882.575 641.200 ;
    END
  END rdata[7]
  PIN rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 650.120 882.575 650.720 ;
    END
  END rdata[8]
  PIN rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 878.575 659.640 882.575 660.240 ;
    END
  END rdata[9]
  PIN wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 269.320 882.575 269.920 ;
    END
  END wdata[0]
  PIN wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 364.520 882.575 365.120 ;
    END
  END wdata[10]
  PIN wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 374.040 882.575 374.640 ;
    END
  END wdata[11]
  PIN wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 383.560 882.575 384.160 ;
    END
  END wdata[12]
  PIN wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 393.080 882.575 393.680 ;
    END
  END wdata[13]
  PIN wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 402.600 882.575 403.200 ;
    END
  END wdata[14]
  PIN wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 412.120 882.575 412.720 ;
    END
  END wdata[15]
  PIN wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 421.640 882.575 422.240 ;
    END
  END wdata[16]
  PIN wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 431.160 882.575 431.760 ;
    END
  END wdata[17]
  PIN wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 440.680 882.575 441.280 ;
    END
  END wdata[18]
  PIN wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 450.200 882.575 450.800 ;
    END
  END wdata[19]
  PIN wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 278.840 882.575 279.440 ;
    END
  END wdata[1]
  PIN wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 459.720 882.575 460.320 ;
    END
  END wdata[20]
  PIN wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 469.240 882.575 469.840 ;
    END
  END wdata[21]
  PIN wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 478.760 882.575 479.360 ;
    END
  END wdata[22]
  PIN wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 488.280 882.575 488.880 ;
    END
  END wdata[23]
  PIN wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 497.800 882.575 498.400 ;
    END
  END wdata[24]
  PIN wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 507.320 882.575 507.920 ;
    END
  END wdata[25]
  PIN wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 516.840 882.575 517.440 ;
    END
  END wdata[26]
  PIN wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 526.360 882.575 526.960 ;
    END
  END wdata[27]
  PIN wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 535.880 882.575 536.480 ;
    END
  END wdata[28]
  PIN wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 545.400 882.575 546.000 ;
    END
  END wdata[29]
  PIN wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 288.360 882.575 288.960 ;
    END
  END wdata[2]
  PIN wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 554.920 882.575 555.520 ;
    END
  END wdata[30]
  PIN wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 564.440 882.575 565.040 ;
    END
  END wdata[31]
  PIN wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 297.880 882.575 298.480 ;
    END
  END wdata[3]
  PIN wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 307.400 882.575 308.000 ;
    END
  END wdata[4]
  PIN wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 316.920 882.575 317.520 ;
    END
  END wdata[5]
  PIN wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 326.440 882.575 327.040 ;
    END
  END wdata[6]
  PIN wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 335.960 882.575 336.560 ;
    END
  END wdata[7]
  PIN wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 345.480 882.575 346.080 ;
    END
  END wdata[8]
  PIN wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 355.000 882.575 355.600 ;
    END
  END wdata[9]
  PIN wen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 21.800 882.575 22.400 ;
    END
  END wen[0]
  PIN wen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 31.320 882.575 31.920 ;
    END
  END wen[1]
  PIN wen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 878.575 40.840 882.575 41.440 ;
    END
  END wen[2]
  PIN wen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 878.575 50.360 882.575 50.960 ;
    END
  END wen[3]
  OBS
      LAYER nwell ;
        RECT 5.330 877.145 876.950 879.975 ;
        RECT 5.330 871.705 876.950 874.535 ;
        RECT 5.330 866.265 876.950 869.095 ;
        RECT 5.330 860.825 876.950 863.655 ;
        RECT 5.330 855.385 876.950 858.215 ;
        RECT 5.330 849.945 876.950 852.775 ;
        RECT 5.330 844.505 876.950 847.335 ;
        RECT 5.330 839.065 876.950 841.895 ;
        RECT 5.330 833.625 876.950 836.455 ;
        RECT 5.330 828.185 876.950 831.015 ;
        RECT 5.330 822.745 876.950 825.575 ;
        RECT 5.330 817.305 876.950 820.135 ;
        RECT 5.330 811.865 876.950 814.695 ;
        RECT 5.330 806.425 876.950 809.255 ;
        RECT 5.330 800.985 876.950 803.815 ;
        RECT 5.330 795.545 876.950 798.375 ;
        RECT 5.330 790.105 876.950 792.935 ;
        RECT 5.330 784.665 876.950 787.495 ;
        RECT 5.330 779.225 876.950 782.055 ;
        RECT 5.330 773.785 876.950 776.615 ;
        RECT 5.330 768.345 876.950 771.175 ;
        RECT 5.330 762.905 876.950 765.735 ;
        RECT 5.330 757.465 876.950 760.295 ;
        RECT 5.330 752.025 876.950 754.855 ;
        RECT 5.330 746.585 876.950 749.415 ;
        RECT 5.330 741.145 876.950 743.975 ;
        RECT 5.330 735.705 876.950 738.535 ;
        RECT 5.330 730.265 876.950 733.095 ;
        RECT 5.330 724.825 876.950 727.655 ;
        RECT 5.330 719.385 876.950 722.215 ;
        RECT 5.330 713.945 876.950 716.775 ;
        RECT 5.330 708.505 876.950 711.335 ;
        RECT 5.330 703.065 876.950 705.895 ;
        RECT 5.330 697.625 876.950 700.455 ;
        RECT 5.330 692.185 876.950 695.015 ;
        RECT 5.330 686.745 876.950 689.575 ;
        RECT 5.330 681.305 876.950 684.135 ;
        RECT 5.330 675.865 876.950 678.695 ;
        RECT 5.330 670.425 876.950 673.255 ;
        RECT 5.330 664.985 876.950 667.815 ;
        RECT 5.330 659.545 876.950 662.375 ;
        RECT 5.330 654.105 876.950 656.935 ;
        RECT 5.330 648.665 876.950 651.495 ;
        RECT 5.330 643.225 876.950 646.055 ;
        RECT 5.330 637.785 876.950 640.615 ;
        RECT 5.330 632.345 876.950 635.175 ;
        RECT 5.330 626.905 876.950 629.735 ;
        RECT 5.330 621.465 876.950 624.295 ;
        RECT 5.330 616.025 876.950 618.855 ;
        RECT 5.330 610.585 876.950 613.415 ;
        RECT 5.330 605.145 876.950 607.975 ;
        RECT 5.330 599.705 876.950 602.535 ;
        RECT 5.330 594.265 876.950 597.095 ;
        RECT 5.330 588.825 876.950 591.655 ;
        RECT 5.330 583.385 876.950 586.215 ;
        RECT 5.330 577.945 876.950 580.775 ;
        RECT 5.330 572.505 876.950 575.335 ;
        RECT 5.330 567.065 876.950 569.895 ;
        RECT 5.330 561.625 876.950 564.455 ;
        RECT 5.330 556.185 876.950 559.015 ;
        RECT 5.330 550.745 876.950 553.575 ;
        RECT 5.330 545.305 876.950 548.135 ;
        RECT 5.330 539.865 876.950 542.695 ;
        RECT 5.330 534.425 876.950 537.255 ;
        RECT 5.330 528.985 876.950 531.815 ;
        RECT 5.330 523.545 876.950 526.375 ;
        RECT 5.330 518.105 876.950 520.935 ;
        RECT 5.330 512.665 876.950 515.495 ;
        RECT 5.330 507.225 876.950 510.055 ;
        RECT 5.330 501.785 876.950 504.615 ;
        RECT 5.330 496.345 876.950 499.175 ;
        RECT 5.330 490.905 876.950 493.735 ;
        RECT 5.330 485.465 876.950 488.295 ;
        RECT 5.330 480.025 876.950 482.855 ;
        RECT 5.330 474.585 876.950 477.415 ;
        RECT 5.330 469.145 876.950 471.975 ;
        RECT 5.330 463.705 876.950 466.535 ;
        RECT 5.330 458.265 876.950 461.095 ;
        RECT 5.330 452.825 876.950 455.655 ;
        RECT 5.330 447.385 876.950 450.215 ;
        RECT 5.330 441.945 876.950 444.775 ;
        RECT 5.330 436.505 876.950 439.335 ;
        RECT 5.330 431.065 876.950 433.895 ;
        RECT 5.330 425.625 876.950 428.455 ;
        RECT 5.330 420.185 876.950 423.015 ;
        RECT 5.330 414.745 876.950 417.575 ;
        RECT 5.330 409.305 876.950 412.135 ;
        RECT 5.330 403.865 876.950 406.695 ;
        RECT 5.330 398.425 876.950 401.255 ;
        RECT 5.330 392.985 876.950 395.815 ;
        RECT 5.330 387.545 876.950 390.375 ;
        RECT 5.330 382.105 876.950 384.935 ;
        RECT 5.330 376.665 876.950 379.495 ;
        RECT 5.330 371.225 876.950 374.055 ;
        RECT 5.330 365.785 876.950 368.615 ;
        RECT 5.330 360.345 876.950 363.175 ;
        RECT 5.330 354.905 876.950 357.735 ;
        RECT 5.330 349.465 876.950 352.295 ;
        RECT 5.330 344.025 876.950 346.855 ;
        RECT 5.330 338.585 876.950 341.415 ;
        RECT 5.330 333.145 876.950 335.975 ;
        RECT 5.330 327.705 876.950 330.535 ;
        RECT 5.330 322.265 876.950 325.095 ;
        RECT 5.330 316.825 876.950 319.655 ;
        RECT 5.330 311.385 876.950 314.215 ;
        RECT 5.330 305.945 876.950 308.775 ;
        RECT 5.330 300.505 876.950 303.335 ;
        RECT 5.330 295.065 876.950 297.895 ;
        RECT 5.330 289.625 876.950 292.455 ;
        RECT 5.330 284.185 876.950 287.015 ;
        RECT 5.330 278.745 876.950 281.575 ;
        RECT 5.330 273.305 876.950 276.135 ;
        RECT 5.330 267.865 876.950 270.695 ;
        RECT 5.330 262.425 876.950 265.255 ;
        RECT 5.330 256.985 876.950 259.815 ;
        RECT 5.330 251.545 876.950 254.375 ;
        RECT 5.330 246.105 876.950 248.935 ;
        RECT 5.330 240.665 876.950 243.495 ;
        RECT 5.330 235.225 876.950 238.055 ;
        RECT 5.330 229.785 876.950 232.615 ;
        RECT 5.330 224.345 876.950 227.175 ;
        RECT 5.330 218.905 876.950 221.735 ;
        RECT 5.330 213.465 876.950 216.295 ;
        RECT 5.330 208.025 876.950 210.855 ;
        RECT 5.330 202.585 876.950 205.415 ;
        RECT 5.330 197.145 876.950 199.975 ;
        RECT 5.330 191.705 876.950 194.535 ;
        RECT 5.330 186.265 876.950 189.095 ;
        RECT 5.330 180.825 876.950 183.655 ;
        RECT 5.330 175.385 876.950 178.215 ;
        RECT 5.330 169.945 876.950 172.775 ;
        RECT 5.330 164.505 876.950 167.335 ;
        RECT 5.330 159.065 876.950 161.895 ;
        RECT 5.330 153.625 876.950 156.455 ;
        RECT 5.330 148.185 876.950 151.015 ;
        RECT 5.330 142.745 876.950 145.575 ;
        RECT 5.330 137.305 876.950 140.135 ;
        RECT 5.330 131.865 876.950 134.695 ;
        RECT 5.330 126.425 876.950 129.255 ;
        RECT 5.330 120.985 876.950 123.815 ;
        RECT 5.330 115.545 876.950 118.375 ;
        RECT 5.330 110.105 876.950 112.935 ;
        RECT 5.330 104.665 876.950 107.495 ;
        RECT 5.330 99.225 876.950 102.055 ;
        RECT 5.330 93.785 876.950 96.615 ;
        RECT 5.330 88.345 876.950 91.175 ;
        RECT 5.330 82.905 876.950 85.735 ;
        RECT 5.330 77.465 876.950 80.295 ;
        RECT 5.330 72.025 876.950 74.855 ;
        RECT 5.330 66.585 876.950 69.415 ;
        RECT 5.330 61.145 876.950 63.975 ;
        RECT 5.330 55.705 876.950 58.535 ;
        RECT 5.330 50.265 876.950 53.095 ;
        RECT 5.330 44.825 876.950 47.655 ;
        RECT 5.330 39.385 876.950 42.215 ;
        RECT 5.330 33.945 876.950 36.775 ;
        RECT 5.330 28.505 876.950 31.335 ;
        RECT 5.330 23.065 876.950 25.895 ;
        RECT 5.330 17.625 876.950 20.455 ;
        RECT 5.330 12.185 876.950 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 876.760 881.365 ;
      LAYER met1 ;
        RECT 5.520 10.640 878.070 881.920 ;
      LAYER met2 ;
        RECT 7.000 4.280 878.050 881.950 ;
        RECT 7.000 4.000 440.490 4.280 ;
        RECT 441.330 4.000 878.050 4.280 ;
      LAYER met3 ;
        RECT 21.050 870.080 878.575 881.445 ;
        RECT 21.050 868.680 878.175 870.080 ;
        RECT 21.050 860.560 878.575 868.680 ;
        RECT 21.050 859.160 878.175 860.560 ;
        RECT 21.050 851.040 878.575 859.160 ;
        RECT 21.050 849.640 878.175 851.040 ;
        RECT 21.050 841.520 878.575 849.640 ;
        RECT 21.050 840.120 878.175 841.520 ;
        RECT 21.050 832.000 878.575 840.120 ;
        RECT 21.050 830.600 878.175 832.000 ;
        RECT 21.050 822.480 878.575 830.600 ;
        RECT 21.050 821.080 878.175 822.480 ;
        RECT 21.050 812.960 878.575 821.080 ;
        RECT 21.050 811.560 878.175 812.960 ;
        RECT 21.050 803.440 878.575 811.560 ;
        RECT 21.050 802.040 878.175 803.440 ;
        RECT 21.050 793.920 878.575 802.040 ;
        RECT 21.050 792.520 878.175 793.920 ;
        RECT 21.050 784.400 878.575 792.520 ;
        RECT 21.050 783.000 878.175 784.400 ;
        RECT 21.050 774.880 878.575 783.000 ;
        RECT 21.050 773.480 878.175 774.880 ;
        RECT 21.050 765.360 878.575 773.480 ;
        RECT 21.050 763.960 878.175 765.360 ;
        RECT 21.050 755.840 878.575 763.960 ;
        RECT 21.050 754.440 878.175 755.840 ;
        RECT 21.050 746.320 878.575 754.440 ;
        RECT 21.050 744.920 878.175 746.320 ;
        RECT 21.050 736.800 878.575 744.920 ;
        RECT 21.050 735.400 878.175 736.800 ;
        RECT 21.050 727.280 878.575 735.400 ;
        RECT 21.050 725.880 878.175 727.280 ;
        RECT 21.050 717.760 878.575 725.880 ;
        RECT 21.050 716.360 878.175 717.760 ;
        RECT 21.050 708.240 878.575 716.360 ;
        RECT 21.050 706.840 878.175 708.240 ;
        RECT 21.050 698.720 878.575 706.840 ;
        RECT 21.050 697.320 878.175 698.720 ;
        RECT 21.050 689.200 878.575 697.320 ;
        RECT 21.050 687.800 878.175 689.200 ;
        RECT 21.050 679.680 878.575 687.800 ;
        RECT 21.050 678.280 878.175 679.680 ;
        RECT 21.050 670.160 878.575 678.280 ;
        RECT 21.050 668.760 878.175 670.160 ;
        RECT 21.050 660.640 878.575 668.760 ;
        RECT 21.050 659.240 878.175 660.640 ;
        RECT 21.050 651.120 878.575 659.240 ;
        RECT 21.050 649.720 878.175 651.120 ;
        RECT 21.050 641.600 878.575 649.720 ;
        RECT 21.050 640.200 878.175 641.600 ;
        RECT 21.050 632.080 878.575 640.200 ;
        RECT 21.050 630.680 878.175 632.080 ;
        RECT 21.050 622.560 878.575 630.680 ;
        RECT 21.050 621.160 878.175 622.560 ;
        RECT 21.050 613.040 878.575 621.160 ;
        RECT 21.050 611.640 878.175 613.040 ;
        RECT 21.050 603.520 878.575 611.640 ;
        RECT 21.050 602.120 878.175 603.520 ;
        RECT 21.050 594.000 878.575 602.120 ;
        RECT 21.050 592.600 878.175 594.000 ;
        RECT 21.050 584.480 878.575 592.600 ;
        RECT 21.050 583.080 878.175 584.480 ;
        RECT 21.050 574.960 878.575 583.080 ;
        RECT 21.050 573.560 878.175 574.960 ;
        RECT 21.050 565.440 878.575 573.560 ;
        RECT 21.050 564.040 878.175 565.440 ;
        RECT 21.050 555.920 878.575 564.040 ;
        RECT 21.050 554.520 878.175 555.920 ;
        RECT 21.050 546.400 878.575 554.520 ;
        RECT 21.050 545.000 878.175 546.400 ;
        RECT 21.050 536.880 878.575 545.000 ;
        RECT 21.050 535.480 878.175 536.880 ;
        RECT 21.050 527.360 878.575 535.480 ;
        RECT 21.050 525.960 878.175 527.360 ;
        RECT 21.050 517.840 878.575 525.960 ;
        RECT 21.050 516.440 878.175 517.840 ;
        RECT 21.050 508.320 878.575 516.440 ;
        RECT 21.050 506.920 878.175 508.320 ;
        RECT 21.050 498.800 878.575 506.920 ;
        RECT 21.050 497.400 878.175 498.800 ;
        RECT 21.050 489.280 878.575 497.400 ;
        RECT 21.050 487.880 878.175 489.280 ;
        RECT 21.050 479.760 878.575 487.880 ;
        RECT 21.050 478.360 878.175 479.760 ;
        RECT 21.050 470.240 878.575 478.360 ;
        RECT 21.050 468.840 878.175 470.240 ;
        RECT 21.050 460.720 878.575 468.840 ;
        RECT 21.050 459.320 878.175 460.720 ;
        RECT 21.050 451.200 878.575 459.320 ;
        RECT 21.050 449.800 878.175 451.200 ;
        RECT 21.050 441.680 878.575 449.800 ;
        RECT 21.050 440.280 878.175 441.680 ;
        RECT 21.050 432.160 878.575 440.280 ;
        RECT 21.050 430.760 878.175 432.160 ;
        RECT 21.050 422.640 878.575 430.760 ;
        RECT 21.050 421.240 878.175 422.640 ;
        RECT 21.050 413.120 878.575 421.240 ;
        RECT 21.050 411.720 878.175 413.120 ;
        RECT 21.050 403.600 878.575 411.720 ;
        RECT 21.050 402.200 878.175 403.600 ;
        RECT 21.050 394.080 878.575 402.200 ;
        RECT 21.050 392.680 878.175 394.080 ;
        RECT 21.050 384.560 878.575 392.680 ;
        RECT 21.050 383.160 878.175 384.560 ;
        RECT 21.050 375.040 878.575 383.160 ;
        RECT 21.050 373.640 878.175 375.040 ;
        RECT 21.050 365.520 878.575 373.640 ;
        RECT 21.050 364.120 878.175 365.520 ;
        RECT 21.050 356.000 878.575 364.120 ;
        RECT 21.050 354.600 878.175 356.000 ;
        RECT 21.050 346.480 878.575 354.600 ;
        RECT 21.050 345.080 878.175 346.480 ;
        RECT 21.050 336.960 878.575 345.080 ;
        RECT 21.050 335.560 878.175 336.960 ;
        RECT 21.050 327.440 878.575 335.560 ;
        RECT 21.050 326.040 878.175 327.440 ;
        RECT 21.050 317.920 878.575 326.040 ;
        RECT 21.050 316.520 878.175 317.920 ;
        RECT 21.050 308.400 878.575 316.520 ;
        RECT 21.050 307.000 878.175 308.400 ;
        RECT 21.050 298.880 878.575 307.000 ;
        RECT 21.050 297.480 878.175 298.880 ;
        RECT 21.050 289.360 878.575 297.480 ;
        RECT 21.050 287.960 878.175 289.360 ;
        RECT 21.050 279.840 878.575 287.960 ;
        RECT 21.050 278.440 878.175 279.840 ;
        RECT 21.050 270.320 878.575 278.440 ;
        RECT 21.050 268.920 878.175 270.320 ;
        RECT 21.050 260.800 878.575 268.920 ;
        RECT 21.050 259.400 878.175 260.800 ;
        RECT 21.050 251.280 878.575 259.400 ;
        RECT 21.050 249.880 878.175 251.280 ;
        RECT 21.050 241.760 878.575 249.880 ;
        RECT 21.050 240.360 878.175 241.760 ;
        RECT 21.050 232.240 878.575 240.360 ;
        RECT 21.050 230.840 878.175 232.240 ;
        RECT 21.050 222.720 878.575 230.840 ;
        RECT 21.050 221.320 878.175 222.720 ;
        RECT 21.050 213.200 878.575 221.320 ;
        RECT 21.050 211.800 878.175 213.200 ;
        RECT 21.050 203.680 878.575 211.800 ;
        RECT 21.050 202.280 878.175 203.680 ;
        RECT 21.050 194.160 878.575 202.280 ;
        RECT 21.050 192.760 878.175 194.160 ;
        RECT 21.050 184.640 878.575 192.760 ;
        RECT 21.050 183.240 878.175 184.640 ;
        RECT 21.050 175.120 878.575 183.240 ;
        RECT 21.050 173.720 878.175 175.120 ;
        RECT 21.050 165.600 878.575 173.720 ;
        RECT 21.050 164.200 878.175 165.600 ;
        RECT 21.050 156.080 878.575 164.200 ;
        RECT 21.050 154.680 878.175 156.080 ;
        RECT 21.050 146.560 878.575 154.680 ;
        RECT 21.050 145.160 878.175 146.560 ;
        RECT 21.050 137.040 878.575 145.160 ;
        RECT 21.050 135.640 878.175 137.040 ;
        RECT 21.050 127.520 878.575 135.640 ;
        RECT 21.050 126.120 878.175 127.520 ;
        RECT 21.050 118.000 878.575 126.120 ;
        RECT 21.050 116.600 878.175 118.000 ;
        RECT 21.050 108.480 878.575 116.600 ;
        RECT 21.050 107.080 878.175 108.480 ;
        RECT 21.050 98.960 878.575 107.080 ;
        RECT 21.050 97.560 878.175 98.960 ;
        RECT 21.050 89.440 878.575 97.560 ;
        RECT 21.050 88.040 878.175 89.440 ;
        RECT 21.050 79.920 878.575 88.040 ;
        RECT 21.050 78.520 878.175 79.920 ;
        RECT 21.050 70.400 878.575 78.520 ;
        RECT 21.050 69.000 878.175 70.400 ;
        RECT 21.050 60.880 878.575 69.000 ;
        RECT 21.050 59.480 878.175 60.880 ;
        RECT 21.050 51.360 878.575 59.480 ;
        RECT 21.050 49.960 878.175 51.360 ;
        RECT 21.050 41.840 878.575 49.960 ;
        RECT 21.050 40.440 878.175 41.840 ;
        RECT 21.050 32.320 878.575 40.440 ;
        RECT 21.050 30.920 878.175 32.320 ;
        RECT 21.050 22.800 878.575 30.920 ;
        RECT 21.050 21.400 878.175 22.800 ;
        RECT 21.050 10.715 878.575 21.400 ;
      LAYER met4 ;
        RECT 69.295 17.175 97.440 866.145 ;
        RECT 99.840 17.175 174.240 866.145 ;
        RECT 176.640 17.175 251.040 866.145 ;
        RECT 253.440 17.175 327.840 866.145 ;
        RECT 330.240 17.175 404.640 866.145 ;
        RECT 407.040 17.175 481.440 866.145 ;
        RECT 483.840 17.175 558.240 866.145 ;
        RECT 560.640 17.175 635.040 866.145 ;
        RECT 637.440 17.175 711.840 866.145 ;
        RECT 714.240 17.175 788.640 866.145 ;
        RECT 791.040 17.175 865.440 866.145 ;
        RECT 867.840 17.175 869.105 866.145 ;
      LAYER met5 ;
        RECT 130.300 102.900 847.660 774.300 ;
  END
END alphasoc_mem
END LIBRARY

