VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spimemio
  CLASS BLOCK ;
  FOREIGN spimemio ;
  ORIGIN 0.000 0.000 ;
  SIZE 465.515 BY 476.235 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 465.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 465.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 465.360 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 465.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 465.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 465.360 ;
    END
  END VPWR
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 257.080 465.515 257.680 ;
    END
  END addr[0]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 284.280 465.515 284.880 ;
    END
  END addr[10]
  PIN addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 287.000 465.515 287.600 ;
    END
  END addr[11]
  PIN addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 289.720 465.515 290.320 ;
    END
  END addr[12]
  PIN addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 292.440 465.515 293.040 ;
    END
  END addr[13]
  PIN addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 295.160 465.515 295.760 ;
    END
  END addr[14]
  PIN addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 297.880 465.515 298.480 ;
    END
  END addr[15]
  PIN addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 300.600 465.515 301.200 ;
    END
  END addr[16]
  PIN addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 303.320 465.515 303.920 ;
    END
  END addr[17]
  PIN addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 306.040 465.515 306.640 ;
    END
  END addr[18]
  PIN addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 308.760 465.515 309.360 ;
    END
  END addr[19]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 259.800 465.515 260.400 ;
    END
  END addr[1]
  PIN addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 311.480 465.515 312.080 ;
    END
  END addr[20]
  PIN addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 314.200 465.515 314.800 ;
    END
  END addr[21]
  PIN addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 316.920 465.515 317.520 ;
    END
  END addr[22]
  PIN addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 319.640 465.515 320.240 ;
    END
  END addr[23]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 262.520 465.515 263.120 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 265.240 465.515 265.840 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 267.960 465.515 268.560 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 270.680 465.515 271.280 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 273.400 465.515 274.000 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 276.120 465.515 276.720 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 278.840 465.515 279.440 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 281.560 465.515 282.160 ;
    END
  END addr[9]
  PIN cfgreg_di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 80.280 465.515 80.880 ;
    END
  END cfgreg_di[0]
  PIN cfgreg_di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 107.480 465.515 108.080 ;
    END
  END cfgreg_di[10]
  PIN cfgreg_di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 110.200 465.515 110.800 ;
    END
  END cfgreg_di[11]
  PIN cfgreg_di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 112.920 465.515 113.520 ;
    END
  END cfgreg_di[12]
  PIN cfgreg_di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 115.640 465.515 116.240 ;
    END
  END cfgreg_di[13]
  PIN cfgreg_di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 118.360 465.515 118.960 ;
    END
  END cfgreg_di[14]
  PIN cfgreg_di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 121.080 465.515 121.680 ;
    END
  END cfgreg_di[15]
  PIN cfgreg_di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 123.800 465.515 124.400 ;
    END
  END cfgreg_di[16]
  PIN cfgreg_di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 126.520 465.515 127.120 ;
    END
  END cfgreg_di[17]
  PIN cfgreg_di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 129.240 465.515 129.840 ;
    END
  END cfgreg_di[18]
  PIN cfgreg_di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 131.960 465.515 132.560 ;
    END
  END cfgreg_di[19]
  PIN cfgreg_di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 83.000 465.515 83.600 ;
    END
  END cfgreg_di[1]
  PIN cfgreg_di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 134.680 465.515 135.280 ;
    END
  END cfgreg_di[20]
  PIN cfgreg_di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 137.400 465.515 138.000 ;
    END
  END cfgreg_di[21]
  PIN cfgreg_di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 140.120 465.515 140.720 ;
    END
  END cfgreg_di[22]
  PIN cfgreg_di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 142.840 465.515 143.440 ;
    END
  END cfgreg_di[23]
  PIN cfgreg_di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 145.560 465.515 146.160 ;
    END
  END cfgreg_di[24]
  PIN cfgreg_di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 148.280 465.515 148.880 ;
    END
  END cfgreg_di[25]
  PIN cfgreg_di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 151.000 465.515 151.600 ;
    END
  END cfgreg_di[26]
  PIN cfgreg_di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 153.720 465.515 154.320 ;
    END
  END cfgreg_di[27]
  PIN cfgreg_di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 156.440 465.515 157.040 ;
    END
  END cfgreg_di[28]
  PIN cfgreg_di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 159.160 465.515 159.760 ;
    END
  END cfgreg_di[29]
  PIN cfgreg_di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 85.720 465.515 86.320 ;
    END
  END cfgreg_di[2]
  PIN cfgreg_di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 161.880 465.515 162.480 ;
    END
  END cfgreg_di[30]
  PIN cfgreg_di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 164.600 465.515 165.200 ;
    END
  END cfgreg_di[31]
  PIN cfgreg_di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 88.440 465.515 89.040 ;
    END
  END cfgreg_di[3]
  PIN cfgreg_di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 91.160 465.515 91.760 ;
    END
  END cfgreg_di[4]
  PIN cfgreg_di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 93.880 465.515 94.480 ;
    END
  END cfgreg_di[5]
  PIN cfgreg_di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 96.600 465.515 97.200 ;
    END
  END cfgreg_di[6]
  PIN cfgreg_di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 99.320 465.515 99.920 ;
    END
  END cfgreg_di[7]
  PIN cfgreg_di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 102.040 465.515 102.640 ;
    END
  END cfgreg_di[8]
  PIN cfgreg_di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 461.515 104.760 465.515 105.360 ;
    END
  END cfgreg_di[9]
  PIN cfgreg_do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 167.320 465.515 167.920 ;
    END
  END cfgreg_do[0]
  PIN cfgreg_do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 194.520 465.515 195.120 ;
    END
  END cfgreg_do[10]
  PIN cfgreg_do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 197.240 465.515 197.840 ;
    END
  END cfgreg_do[11]
  PIN cfgreg_do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 199.960 465.515 200.560 ;
    END
  END cfgreg_do[12]
  PIN cfgreg_do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 202.680 465.515 203.280 ;
    END
  END cfgreg_do[13]
  PIN cfgreg_do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 205.400 465.515 206.000 ;
    END
  END cfgreg_do[14]
  PIN cfgreg_do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 208.120 465.515 208.720 ;
    END
  END cfgreg_do[15]
  PIN cfgreg_do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 210.840 465.515 211.440 ;
    END
  END cfgreg_do[16]
  PIN cfgreg_do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 213.560 465.515 214.160 ;
    END
  END cfgreg_do[17]
  PIN cfgreg_do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 216.280 465.515 216.880 ;
    END
  END cfgreg_do[18]
  PIN cfgreg_do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 219.000 465.515 219.600 ;
    END
  END cfgreg_do[19]
  PIN cfgreg_do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 170.040 465.515 170.640 ;
    END
  END cfgreg_do[1]
  PIN cfgreg_do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 221.720 465.515 222.320 ;
    END
  END cfgreg_do[20]
  PIN cfgreg_do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 224.440 465.515 225.040 ;
    END
  END cfgreg_do[21]
  PIN cfgreg_do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 227.160 465.515 227.760 ;
    END
  END cfgreg_do[22]
  PIN cfgreg_do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 229.880 465.515 230.480 ;
    END
  END cfgreg_do[23]
  PIN cfgreg_do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 232.600 465.515 233.200 ;
    END
  END cfgreg_do[24]
  PIN cfgreg_do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 235.320 465.515 235.920 ;
    END
  END cfgreg_do[25]
  PIN cfgreg_do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 238.040 465.515 238.640 ;
    END
  END cfgreg_do[26]
  PIN cfgreg_do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 240.760 465.515 241.360 ;
    END
  END cfgreg_do[27]
  PIN cfgreg_do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 243.480 465.515 244.080 ;
    END
  END cfgreg_do[28]
  PIN cfgreg_do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 246.200 465.515 246.800 ;
    END
  END cfgreg_do[29]
  PIN cfgreg_do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 172.760 465.515 173.360 ;
    END
  END cfgreg_do[2]
  PIN cfgreg_do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 248.920 465.515 249.520 ;
    END
  END cfgreg_do[30]
  PIN cfgreg_do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 251.640 465.515 252.240 ;
    END
  END cfgreg_do[31]
  PIN cfgreg_do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 175.480 465.515 176.080 ;
    END
  END cfgreg_do[3]
  PIN cfgreg_do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 178.200 465.515 178.800 ;
    END
  END cfgreg_do[4]
  PIN cfgreg_do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 180.920 465.515 181.520 ;
    END
  END cfgreg_do[5]
  PIN cfgreg_do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 183.640 465.515 184.240 ;
    END
  END cfgreg_do[6]
  PIN cfgreg_do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 461.515 186.360 465.515 186.960 ;
    END
  END cfgreg_do[7]
  PIN cfgreg_do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 189.080 465.515 189.680 ;
    END
  END cfgreg_do[8]
  PIN cfgreg_do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 191.800 465.515 192.400 ;
    END
  END cfgreg_do[9]
  PIN cfgreg_we[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 69.400 465.515 70.000 ;
    END
  END cfgreg_we[0]
  PIN cfgreg_we[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 72.120 465.515 72.720 ;
    END
  END cfgreg_we[1]
  PIN cfgreg_we[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 74.840 465.515 75.440 ;
    END
  END cfgreg_we[2]
  PIN cfgreg_we[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 77.560 465.515 78.160 ;
    END
  END cfgreg_we[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END clk
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END flash_clk
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END flash_csb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END flash_io0_do
  PIN flash_io0_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END flash_io0_oe
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END flash_io1_do
  PIN flash_io1_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END flash_io1_oe
  PIN flash_io2_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END flash_io2_di
  PIN flash_io2_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END flash_io2_do
  PIN flash_io2_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END flash_io2_oe
  PIN flash_io3_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END flash_io3_di
  PIN flash_io3_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END flash_io3_do
  PIN flash_io3_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END flash_io3_oe
  PIN rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 322.360 465.515 322.960 ;
    END
  END rdata[0]
  PIN rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 349.560 465.515 350.160 ;
    END
  END rdata[10]
  PIN rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 352.280 465.515 352.880 ;
    END
  END rdata[11]
  PIN rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 355.000 465.515 355.600 ;
    END
  END rdata[12]
  PIN rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 357.720 465.515 358.320 ;
    END
  END rdata[13]
  PIN rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 360.440 465.515 361.040 ;
    END
  END rdata[14]
  PIN rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 363.160 465.515 363.760 ;
    END
  END rdata[15]
  PIN rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 365.880 465.515 366.480 ;
    END
  END rdata[16]
  PIN rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 368.600 465.515 369.200 ;
    END
  END rdata[17]
  PIN rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 371.320 465.515 371.920 ;
    END
  END rdata[18]
  PIN rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 374.040 465.515 374.640 ;
    END
  END rdata[19]
  PIN rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 325.080 465.515 325.680 ;
    END
  END rdata[1]
  PIN rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 376.760 465.515 377.360 ;
    END
  END rdata[20]
  PIN rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 379.480 465.515 380.080 ;
    END
  END rdata[21]
  PIN rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 382.200 465.515 382.800 ;
    END
  END rdata[22]
  PIN rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 384.920 465.515 385.520 ;
    END
  END rdata[23]
  PIN rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 387.640 465.515 388.240 ;
    END
  END rdata[24]
  PIN rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 390.360 465.515 390.960 ;
    END
  END rdata[25]
  PIN rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 393.080 465.515 393.680 ;
    END
  END rdata[26]
  PIN rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 395.800 465.515 396.400 ;
    END
  END rdata[27]
  PIN rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 398.520 465.515 399.120 ;
    END
  END rdata[28]
  PIN rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 401.240 465.515 401.840 ;
    END
  END rdata[29]
  PIN rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 327.800 465.515 328.400 ;
    END
  END rdata[2]
  PIN rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 403.960 465.515 404.560 ;
    END
  END rdata[30]
  PIN rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 406.680 465.515 407.280 ;
    END
  END rdata[31]
  PIN rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 330.520 465.515 331.120 ;
    END
  END rdata[3]
  PIN rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 333.240 465.515 333.840 ;
    END
  END rdata[4]
  PIN rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 335.960 465.515 336.560 ;
    END
  END rdata[5]
  PIN rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 338.680 465.515 339.280 ;
    END
  END rdata[6]
  PIN rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 341.400 465.515 342.000 ;
    END
  END rdata[7]
  PIN rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 344.120 465.515 344.720 ;
    END
  END rdata[8]
  PIN rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 346.840 465.515 347.440 ;
    END
  END rdata[9]
  PIN ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 461.515 254.360 465.515 254.960 ;
    END
  END ready
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END resetn
  PIN valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 461.515 66.680 465.515 67.280 ;
    END
  END valid
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 459.540 465.205 ;
      LAYER met1 ;
        RECT 4.670 10.240 460.390 465.360 ;
      LAYER met2 ;
        RECT 4.690 4.280 460.370 465.305 ;
        RECT 4.690 4.000 115.730 4.280 ;
        RECT 116.570 4.000 348.490 4.280 ;
        RECT 349.330 4.000 460.370 4.280 ;
      LAYER met3 ;
        RECT 3.990 459.360 461.515 465.285 ;
        RECT 4.400 457.960 461.515 459.360 ;
        RECT 3.990 425.360 461.515 457.960 ;
        RECT 4.400 423.960 461.515 425.360 ;
        RECT 3.990 407.680 461.515 423.960 ;
        RECT 3.990 406.280 461.115 407.680 ;
        RECT 3.990 404.960 461.515 406.280 ;
        RECT 3.990 403.560 461.115 404.960 ;
        RECT 3.990 402.240 461.515 403.560 ;
        RECT 3.990 400.840 461.115 402.240 ;
        RECT 3.990 399.520 461.515 400.840 ;
        RECT 3.990 398.120 461.115 399.520 ;
        RECT 3.990 396.800 461.515 398.120 ;
        RECT 3.990 395.400 461.115 396.800 ;
        RECT 3.990 394.080 461.515 395.400 ;
        RECT 3.990 392.680 461.115 394.080 ;
        RECT 3.990 391.360 461.515 392.680 ;
        RECT 4.400 389.960 461.115 391.360 ;
        RECT 3.990 388.640 461.515 389.960 ;
        RECT 3.990 387.240 461.115 388.640 ;
        RECT 3.990 385.920 461.515 387.240 ;
        RECT 3.990 384.520 461.115 385.920 ;
        RECT 3.990 383.200 461.515 384.520 ;
        RECT 3.990 381.800 461.115 383.200 ;
        RECT 3.990 380.480 461.515 381.800 ;
        RECT 3.990 379.080 461.115 380.480 ;
        RECT 3.990 377.760 461.515 379.080 ;
        RECT 3.990 376.360 461.115 377.760 ;
        RECT 3.990 375.040 461.515 376.360 ;
        RECT 3.990 373.640 461.115 375.040 ;
        RECT 3.990 372.320 461.515 373.640 ;
        RECT 3.990 370.920 461.115 372.320 ;
        RECT 3.990 369.600 461.515 370.920 ;
        RECT 3.990 368.200 461.115 369.600 ;
        RECT 3.990 366.880 461.515 368.200 ;
        RECT 3.990 365.480 461.115 366.880 ;
        RECT 3.990 364.160 461.515 365.480 ;
        RECT 3.990 362.760 461.115 364.160 ;
        RECT 3.990 361.440 461.515 362.760 ;
        RECT 3.990 360.040 461.115 361.440 ;
        RECT 3.990 358.720 461.515 360.040 ;
        RECT 3.990 357.360 461.115 358.720 ;
        RECT 4.400 357.320 461.115 357.360 ;
        RECT 4.400 356.000 461.515 357.320 ;
        RECT 4.400 355.960 461.115 356.000 ;
        RECT 3.990 354.600 461.115 355.960 ;
        RECT 3.990 353.280 461.515 354.600 ;
        RECT 3.990 351.880 461.115 353.280 ;
        RECT 3.990 350.560 461.515 351.880 ;
        RECT 3.990 349.160 461.115 350.560 ;
        RECT 3.990 347.840 461.515 349.160 ;
        RECT 3.990 346.440 461.115 347.840 ;
        RECT 3.990 345.120 461.515 346.440 ;
        RECT 3.990 343.720 461.115 345.120 ;
        RECT 3.990 342.400 461.515 343.720 ;
        RECT 3.990 341.000 461.115 342.400 ;
        RECT 3.990 339.680 461.515 341.000 ;
        RECT 3.990 338.280 461.115 339.680 ;
        RECT 3.990 336.960 461.515 338.280 ;
        RECT 3.990 335.560 461.115 336.960 ;
        RECT 3.990 334.240 461.515 335.560 ;
        RECT 3.990 332.840 461.115 334.240 ;
        RECT 3.990 331.520 461.515 332.840 ;
        RECT 3.990 330.120 461.115 331.520 ;
        RECT 3.990 328.800 461.515 330.120 ;
        RECT 3.990 327.400 461.115 328.800 ;
        RECT 3.990 326.080 461.515 327.400 ;
        RECT 3.990 324.680 461.115 326.080 ;
        RECT 3.990 323.360 461.515 324.680 ;
        RECT 4.400 321.960 461.115 323.360 ;
        RECT 3.990 320.640 461.515 321.960 ;
        RECT 3.990 319.240 461.115 320.640 ;
        RECT 3.990 317.920 461.515 319.240 ;
        RECT 3.990 316.520 461.115 317.920 ;
        RECT 3.990 315.200 461.515 316.520 ;
        RECT 3.990 313.800 461.115 315.200 ;
        RECT 3.990 312.480 461.515 313.800 ;
        RECT 3.990 311.080 461.115 312.480 ;
        RECT 3.990 309.760 461.515 311.080 ;
        RECT 3.990 308.360 461.115 309.760 ;
        RECT 3.990 307.040 461.515 308.360 ;
        RECT 3.990 305.640 461.115 307.040 ;
        RECT 3.990 304.320 461.515 305.640 ;
        RECT 3.990 302.920 461.115 304.320 ;
        RECT 3.990 301.600 461.515 302.920 ;
        RECT 3.990 300.200 461.115 301.600 ;
        RECT 3.990 298.880 461.515 300.200 ;
        RECT 3.990 297.480 461.115 298.880 ;
        RECT 3.990 296.160 461.515 297.480 ;
        RECT 3.990 294.760 461.115 296.160 ;
        RECT 3.990 293.440 461.515 294.760 ;
        RECT 3.990 292.040 461.115 293.440 ;
        RECT 3.990 290.720 461.515 292.040 ;
        RECT 3.990 289.360 461.115 290.720 ;
        RECT 4.400 289.320 461.115 289.360 ;
        RECT 4.400 288.000 461.515 289.320 ;
        RECT 4.400 287.960 461.115 288.000 ;
        RECT 3.990 286.600 461.115 287.960 ;
        RECT 3.990 285.280 461.515 286.600 ;
        RECT 3.990 283.880 461.115 285.280 ;
        RECT 3.990 282.560 461.515 283.880 ;
        RECT 3.990 281.160 461.115 282.560 ;
        RECT 3.990 279.840 461.515 281.160 ;
        RECT 3.990 278.440 461.115 279.840 ;
        RECT 3.990 277.120 461.515 278.440 ;
        RECT 3.990 275.720 461.115 277.120 ;
        RECT 3.990 274.400 461.515 275.720 ;
        RECT 3.990 273.000 461.115 274.400 ;
        RECT 3.990 271.680 461.515 273.000 ;
        RECT 3.990 270.280 461.115 271.680 ;
        RECT 3.990 268.960 461.515 270.280 ;
        RECT 3.990 267.560 461.115 268.960 ;
        RECT 3.990 266.240 461.515 267.560 ;
        RECT 3.990 264.840 461.115 266.240 ;
        RECT 3.990 263.520 461.515 264.840 ;
        RECT 3.990 262.120 461.115 263.520 ;
        RECT 3.990 260.800 461.515 262.120 ;
        RECT 3.990 259.400 461.115 260.800 ;
        RECT 3.990 258.080 461.515 259.400 ;
        RECT 3.990 256.680 461.115 258.080 ;
        RECT 3.990 255.360 461.515 256.680 ;
        RECT 4.400 253.960 461.115 255.360 ;
        RECT 3.990 252.640 461.515 253.960 ;
        RECT 3.990 251.240 461.115 252.640 ;
        RECT 3.990 249.920 461.515 251.240 ;
        RECT 3.990 248.520 461.115 249.920 ;
        RECT 3.990 247.200 461.515 248.520 ;
        RECT 3.990 245.800 461.115 247.200 ;
        RECT 3.990 244.480 461.515 245.800 ;
        RECT 3.990 243.080 461.115 244.480 ;
        RECT 3.990 241.760 461.515 243.080 ;
        RECT 3.990 240.360 461.115 241.760 ;
        RECT 3.990 239.040 461.515 240.360 ;
        RECT 3.990 237.640 461.115 239.040 ;
        RECT 3.990 236.320 461.515 237.640 ;
        RECT 3.990 234.920 461.115 236.320 ;
        RECT 3.990 233.600 461.515 234.920 ;
        RECT 3.990 232.200 461.115 233.600 ;
        RECT 3.990 230.880 461.515 232.200 ;
        RECT 3.990 229.480 461.115 230.880 ;
        RECT 3.990 228.160 461.515 229.480 ;
        RECT 3.990 226.760 461.115 228.160 ;
        RECT 3.990 225.440 461.515 226.760 ;
        RECT 3.990 224.040 461.115 225.440 ;
        RECT 3.990 222.720 461.515 224.040 ;
        RECT 3.990 221.360 461.115 222.720 ;
        RECT 4.400 221.320 461.115 221.360 ;
        RECT 4.400 220.000 461.515 221.320 ;
        RECT 4.400 219.960 461.115 220.000 ;
        RECT 3.990 218.600 461.115 219.960 ;
        RECT 3.990 217.280 461.515 218.600 ;
        RECT 3.990 215.880 461.115 217.280 ;
        RECT 3.990 214.560 461.515 215.880 ;
        RECT 3.990 213.160 461.115 214.560 ;
        RECT 3.990 211.840 461.515 213.160 ;
        RECT 3.990 210.440 461.115 211.840 ;
        RECT 3.990 209.120 461.515 210.440 ;
        RECT 3.990 207.720 461.115 209.120 ;
        RECT 3.990 206.400 461.515 207.720 ;
        RECT 3.990 205.000 461.115 206.400 ;
        RECT 3.990 203.680 461.515 205.000 ;
        RECT 3.990 202.280 461.115 203.680 ;
        RECT 3.990 200.960 461.515 202.280 ;
        RECT 3.990 199.560 461.115 200.960 ;
        RECT 3.990 198.240 461.515 199.560 ;
        RECT 3.990 196.840 461.115 198.240 ;
        RECT 3.990 195.520 461.515 196.840 ;
        RECT 3.990 194.120 461.115 195.520 ;
        RECT 3.990 192.800 461.515 194.120 ;
        RECT 3.990 191.400 461.115 192.800 ;
        RECT 3.990 190.080 461.515 191.400 ;
        RECT 3.990 188.680 461.115 190.080 ;
        RECT 3.990 187.360 461.515 188.680 ;
        RECT 4.400 185.960 461.115 187.360 ;
        RECT 3.990 184.640 461.515 185.960 ;
        RECT 3.990 183.240 461.115 184.640 ;
        RECT 3.990 181.920 461.515 183.240 ;
        RECT 3.990 180.520 461.115 181.920 ;
        RECT 3.990 179.200 461.515 180.520 ;
        RECT 3.990 177.800 461.115 179.200 ;
        RECT 3.990 176.480 461.515 177.800 ;
        RECT 3.990 175.080 461.115 176.480 ;
        RECT 3.990 173.760 461.515 175.080 ;
        RECT 3.990 172.360 461.115 173.760 ;
        RECT 3.990 171.040 461.515 172.360 ;
        RECT 3.990 169.640 461.115 171.040 ;
        RECT 3.990 168.320 461.515 169.640 ;
        RECT 3.990 166.920 461.115 168.320 ;
        RECT 3.990 165.600 461.515 166.920 ;
        RECT 3.990 164.200 461.115 165.600 ;
        RECT 3.990 162.880 461.515 164.200 ;
        RECT 3.990 161.480 461.115 162.880 ;
        RECT 3.990 160.160 461.515 161.480 ;
        RECT 3.990 158.760 461.115 160.160 ;
        RECT 3.990 157.440 461.515 158.760 ;
        RECT 3.990 156.040 461.115 157.440 ;
        RECT 3.990 154.720 461.515 156.040 ;
        RECT 3.990 153.360 461.115 154.720 ;
        RECT 4.400 153.320 461.115 153.360 ;
        RECT 4.400 152.000 461.515 153.320 ;
        RECT 4.400 151.960 461.115 152.000 ;
        RECT 3.990 150.600 461.115 151.960 ;
        RECT 3.990 149.280 461.515 150.600 ;
        RECT 3.990 147.880 461.115 149.280 ;
        RECT 3.990 146.560 461.515 147.880 ;
        RECT 3.990 145.160 461.115 146.560 ;
        RECT 3.990 143.840 461.515 145.160 ;
        RECT 3.990 142.440 461.115 143.840 ;
        RECT 3.990 141.120 461.515 142.440 ;
        RECT 3.990 139.720 461.115 141.120 ;
        RECT 3.990 138.400 461.515 139.720 ;
        RECT 3.990 137.000 461.115 138.400 ;
        RECT 3.990 135.680 461.515 137.000 ;
        RECT 3.990 134.280 461.115 135.680 ;
        RECT 3.990 132.960 461.515 134.280 ;
        RECT 3.990 131.560 461.115 132.960 ;
        RECT 3.990 130.240 461.515 131.560 ;
        RECT 3.990 128.840 461.115 130.240 ;
        RECT 3.990 127.520 461.515 128.840 ;
        RECT 3.990 126.120 461.115 127.520 ;
        RECT 3.990 124.800 461.515 126.120 ;
        RECT 3.990 123.400 461.115 124.800 ;
        RECT 3.990 122.080 461.515 123.400 ;
        RECT 3.990 120.680 461.115 122.080 ;
        RECT 3.990 119.360 461.515 120.680 ;
        RECT 4.400 117.960 461.115 119.360 ;
        RECT 3.990 116.640 461.515 117.960 ;
        RECT 3.990 115.240 461.115 116.640 ;
        RECT 3.990 113.920 461.515 115.240 ;
        RECT 3.990 112.520 461.115 113.920 ;
        RECT 3.990 111.200 461.515 112.520 ;
        RECT 3.990 109.800 461.115 111.200 ;
        RECT 3.990 108.480 461.515 109.800 ;
        RECT 3.990 107.080 461.115 108.480 ;
        RECT 3.990 105.760 461.515 107.080 ;
        RECT 3.990 104.360 461.115 105.760 ;
        RECT 3.990 103.040 461.515 104.360 ;
        RECT 3.990 101.640 461.115 103.040 ;
        RECT 3.990 100.320 461.515 101.640 ;
        RECT 3.990 98.920 461.115 100.320 ;
        RECT 3.990 97.600 461.515 98.920 ;
        RECT 3.990 96.200 461.115 97.600 ;
        RECT 3.990 94.880 461.515 96.200 ;
        RECT 3.990 93.480 461.115 94.880 ;
        RECT 3.990 92.160 461.515 93.480 ;
        RECT 3.990 90.760 461.115 92.160 ;
        RECT 3.990 89.440 461.515 90.760 ;
        RECT 3.990 88.040 461.115 89.440 ;
        RECT 3.990 86.720 461.515 88.040 ;
        RECT 3.990 85.360 461.115 86.720 ;
        RECT 4.400 85.320 461.115 85.360 ;
        RECT 4.400 84.000 461.515 85.320 ;
        RECT 4.400 83.960 461.115 84.000 ;
        RECT 3.990 82.600 461.115 83.960 ;
        RECT 3.990 81.280 461.515 82.600 ;
        RECT 3.990 79.880 461.115 81.280 ;
        RECT 3.990 78.560 461.515 79.880 ;
        RECT 3.990 77.160 461.115 78.560 ;
        RECT 3.990 75.840 461.515 77.160 ;
        RECT 3.990 74.440 461.115 75.840 ;
        RECT 3.990 73.120 461.515 74.440 ;
        RECT 3.990 71.720 461.115 73.120 ;
        RECT 3.990 70.400 461.515 71.720 ;
        RECT 3.990 69.000 461.115 70.400 ;
        RECT 3.990 67.680 461.515 69.000 ;
        RECT 3.990 66.280 461.115 67.680 ;
        RECT 3.990 51.360 461.515 66.280 ;
        RECT 4.400 49.960 461.515 51.360 ;
        RECT 3.990 17.360 461.515 49.960 ;
        RECT 4.400 15.960 461.515 17.360 ;
        RECT 3.990 10.715 461.515 15.960 ;
      LAYER met4 ;
        RECT 317.695 85.855 327.840 345.265 ;
        RECT 330.240 85.855 332.745 345.265 ;
  END
END spimemio
END LIBRARY

