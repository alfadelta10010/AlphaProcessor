module spimemio (clk,
    flash_clk,
    flash_csb,
    flash_io0_di,
    flash_io0_do,
    flash_io0_oe,
    flash_io1_di,
    flash_io1_do,
    flash_io1_oe,
    flash_io2_di,
    flash_io2_do,
    flash_io2_oe,
    flash_io3_di,
    flash_io3_do,
    flash_io3_oe,
    ready,
    resetn,
    valid,
    addr,
    cfgreg_di,
    cfgreg_do,
    cfgreg_we,
    rdata);
 input clk;
 output flash_clk;
 output flash_csb;
 input flash_io0_di;
 output flash_io0_do;
 output flash_io0_oe;
 input flash_io1_di;
 output flash_io1_do;
 output flash_io1_oe;
 input flash_io2_di;
 output flash_io2_do;
 output flash_io2_oe;
 input flash_io3_di;
 output flash_io3_do;
 output flash_io3_oe;
 output ready;
 input resetn;
 input valid;
 input [23:0] addr;
 input [31:0] cfgreg_di;
 output [31:0] cfgreg_do;
 input [3:0] cfgreg_we;
 output [31:0] rdata;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire net129;
 wire net130;
 wire net131;
 wire clknet_0_clk;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire \buffer[0] ;
 wire \buffer[10] ;
 wire \buffer[11] ;
 wire \buffer[12] ;
 wire \buffer[13] ;
 wire \buffer[14] ;
 wire \buffer[15] ;
 wire \buffer[16] ;
 wire \buffer[17] ;
 wire \buffer[18] ;
 wire \buffer[19] ;
 wire \buffer[1] ;
 wire \buffer[20] ;
 wire \buffer[21] ;
 wire \buffer[22] ;
 wire \buffer[23] ;
 wire \buffer[2] ;
 wire \buffer[3] ;
 wire \buffer[4] ;
 wire \buffer[5] ;
 wire \buffer[6] ;
 wire \buffer[7] ;
 wire \buffer[8] ;
 wire \buffer[9] ;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net115;
 wire net116;
 wire config_clk;
 wire config_cont;
 wire config_csb;
 wire config_ddr;
 wire \config_do[0] ;
 wire \config_do[1] ;
 wire \config_do[2] ;
 wire \config_do[3] ;
 wire config_en;
 wire \config_oe[0] ;
 wire \config_oe[1] ;
 wire \config_oe[2] ;
 wire \config_oe[3] ;
 wire config_qspi;
 wire din_ddr;
 wire \rd_addr[0] ;
 wire \rd_addr[10] ;
 wire \rd_addr[11] ;
 wire \rd_addr[12] ;
 wire \rd_addr[13] ;
 wire \rd_addr[14] ;
 wire \rd_addr[15] ;
 wire \rd_addr[16] ;
 wire \rd_addr[17] ;
 wire \rd_addr[18] ;
 wire \rd_addr[19] ;
 wire \rd_addr[1] ;
 wire \rd_addr[20] ;
 wire \rd_addr[21] ;
 wire \rd_addr[22] ;
 wire \rd_addr[23] ;
 wire \rd_addr[2] ;
 wire \rd_addr[3] ;
 wire \rd_addr[4] ;
 wire \rd_addr[5] ;
 wire \rd_addr[6] ;
 wire \rd_addr[7] ;
 wire \rd_addr[8] ;
 wire \rd_addr[9] ;
 wire rd_inc;
 wire rd_valid;
 wire rd_wait;
 wire softreset;
 wire \state[0] ;
 wire \state[10] ;
 wire \state[11] ;
 wire \state[12] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire \state[6] ;
 wire \state[7] ;
 wire \state[8] ;
 wire \state[9] ;
 wire \xfer.count[0] ;
 wire \xfer.count[1] ;
 wire \xfer.count[2] ;
 wire \xfer.count[3] ;
 wire \xfer.din_data[0] ;
 wire \xfer.din_data[1] ;
 wire \xfer.din_data[2] ;
 wire \xfer.din_data[3] ;
 wire \xfer.din_data[4] ;
 wire \xfer.din_data[5] ;
 wire \xfer.din_data[6] ;
 wire \xfer.din_data[7] ;
 wire \xfer.din_qspi ;
 wire \xfer.din_rd ;
 wire \xfer.din_tag[0] ;
 wire \xfer.din_tag[1] ;
 wire \xfer.din_tag[2] ;
 wire \xfer.din_valid ;
 wire \xfer.dout_data[0] ;
 wire \xfer.dout_data[1] ;
 wire \xfer.dout_data[2] ;
 wire \xfer.dout_data[3] ;
 wire \xfer.dout_data[4] ;
 wire \xfer.dout_data[5] ;
 wire \xfer.dout_data[6] ;
 wire \xfer.dout_data[7] ;
 wire \xfer.dout_tag[0] ;
 wire \xfer.dout_tag[1] ;
 wire \xfer.dout_tag[2] ;
 wire \xfer.dummy_count[0] ;
 wire \xfer.dummy_count[1] ;
 wire \xfer.dummy_count[2] ;
 wire \xfer.dummy_count[3] ;
 wire \xfer.fetch ;
 wire \xfer.flash_clk ;
 wire \xfer.flash_csb ;
 wire \xfer.flash_io0_do ;
 wire \xfer.flash_io1_do ;
 wire \xfer.flash_io2_do ;
 wire \xfer.flash_io3_do ;
 wire \xfer.last_fetch ;
 wire \xfer.obuffer[0] ;
 wire \xfer.obuffer[1] ;
 wire \xfer.obuffer[2] ;
 wire \xfer.obuffer[3] ;
 wire \xfer.obuffer[4] ;
 wire \xfer.obuffer[5] ;
 wire \xfer.obuffer[6] ;
 wire \xfer.obuffer[7] ;
 wire \xfer.resetn ;
 wire \xfer.xfer_ddr ;
 wire \xfer.xfer_ddr_q ;
 wire \xfer.xfer_dspi ;
 wire \xfer.xfer_qspi ;
 wire \xfer.xfer_rd ;
 wire \xfer.xfer_tag[0] ;
 wire \xfer.xfer_tag[1] ;
 wire \xfer.xfer_tag[2] ;
 wire xfer_io0_90;
 wire xfer_io1_90;
 wire xfer_io2_90;
 wire xfer_io3_90;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sky130_fd_sc_hd__xor2_1 _0766_ (.A(\rd_addr[10] ),
    .B(net2),
    .X(_0314_));
 sky130_fd_sc_hd__xnor2_2 _0767_ (.A(\rd_addr[19] ),
    .B(net11),
    .Y(_0315_));
 sky130_fd_sc_hd__xnor2_2 _0768_ (.A(\rd_addr[23] ),
    .B(net16),
    .Y(_0316_));
 sky130_fd_sc_hd__nand2_1 _0769_ (.A(_0315_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__xor2_2 _0770_ (.A(\rd_addr[6] ),
    .B(net21),
    .X(_0318_));
 sky130_fd_sc_hd__xor2_2 _0771_ (.A(\rd_addr[11] ),
    .B(net3),
    .X(_0319_));
 sky130_fd_sc_hd__xor2_2 _0772_ (.A(\rd_addr[7] ),
    .B(net22),
    .X(_0320_));
 sky130_fd_sc_hd__xor2_4 _0773_ (.A(\rd_addr[9] ),
    .B(net24),
    .X(_0321_));
 sky130_fd_sc_hd__or4_1 _0774_ (.A(_0318_),
    .B(_0319_),
    .C(_0320_),
    .D(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__xor2_2 _0775_ (.A(\rd_addr[15] ),
    .B(net7),
    .X(_0323_));
 sky130_fd_sc_hd__xor2_2 _0776_ (.A(net17),
    .B(\rd_addr[2] ),
    .X(_0324_));
 sky130_fd_sc_hd__or2b_1 _0777_ (.A(net9),
    .B_N(\rd_addr[17] ),
    .X(_0325_));
 sky130_fd_sc_hd__or2b_1 _0778_ (.A(\rd_addr[17] ),
    .B_N(net9),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_1 _0779_ (.A(_0325_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__xnor2_2 _0780_ (.A(\rd_addr[14] ),
    .B(net6),
    .Y(_0328_));
 sky130_fd_sc_hd__or4b_1 _0781_ (.A(_0323_),
    .B(_0324_),
    .C(_0327_),
    .D_N(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__or4_1 _0782_ (.A(_0314_),
    .B(_0317_),
    .C(_0322_),
    .D(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__and2b_1 _0783_ (.A_N(net13),
    .B(\rd_addr[20] ),
    .X(_0331_));
 sky130_fd_sc_hd__inv_2 _0784_ (.A(net13),
    .Y(_0332_));
 sky130_fd_sc_hd__clkbuf_4 _0785_ (.A(\rd_addr[13] ),
    .X(_0333_));
 sky130_fd_sc_hd__inv_2 _0786_ (.A(net5),
    .Y(_0334_));
 sky130_fd_sc_hd__a2bb2o_1 _0787_ (.A1_N(\rd_addr[20] ),
    .A2_N(_0332_),
    .B1(_0333_),
    .B2(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__inv_2 _0788_ (.A(net18),
    .Y(_0336_));
 sky130_fd_sc_hd__inv_2 _0789_ (.A(\rd_addr[3] ),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_2 _0790_ (.A(\rd_addr[21] ),
    .Y(_0338_));
 sky130_fd_sc_hd__a22o_1 _0791_ (.A1(_0337_),
    .A2(net18),
    .B1(_0338_),
    .B2(net14),
    .X(_0339_));
 sky130_fd_sc_hd__and2b_1 _0792_ (.A_N(net23),
    .B(\rd_addr[8] ),
    .X(_0340_));
 sky130_fd_sc_hd__a211o_1 _0793_ (.A1(\rd_addr[3] ),
    .A2(_0336_),
    .B1(_0339_),
    .C1(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__nand2_1 _0794_ (.A(\rd_addr[0] ),
    .B(net1),
    .Y(_0342_));
 sky130_fd_sc_hd__or2_1 _0795_ (.A(\rd_addr[0] ),
    .B(net1),
    .X(_0343_));
 sky130_fd_sc_hd__xor2_1 _0796_ (.A(\rd_addr[1] ),
    .B(net12),
    .X(_0344_));
 sky130_fd_sc_hd__a21oi_4 _0797_ (.A1(_0342_),
    .A2(_0343_),
    .B1(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__or4b_1 _0798_ (.A(_0331_),
    .B(_0335_),
    .C(_0341_),
    .D_N(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__xor2_2 _0799_ (.A(\rd_addr[5] ),
    .B(net20),
    .X(_0347_));
 sky130_fd_sc_hd__xor2_2 _0800_ (.A(\rd_addr[12] ),
    .B(net4),
    .X(_0348_));
 sky130_fd_sc_hd__xnor2_2 _0801_ (.A(\rd_addr[22] ),
    .B(net15),
    .Y(_0349_));
 sky130_fd_sc_hd__xnor2_2 _0802_ (.A(\rd_addr[18] ),
    .B(net10),
    .Y(_0350_));
 sky130_fd_sc_hd__or4bb_1 _0803_ (.A(_0347_),
    .B(_0348_),
    .C_N(_0349_),
    .D_N(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__inv_2 _0804_ (.A(\rd_addr[4] ),
    .Y(_0352_));
 sky130_fd_sc_hd__and2b_1 _0805_ (.A_N(\rd_addr[8] ),
    .B(net23),
    .X(_0353_));
 sky130_fd_sc_hd__inv_2 _0806_ (.A(\rd_addr[13] ),
    .Y(_0354_));
 sky130_fd_sc_hd__inv_2 _0807_ (.A(net14),
    .Y(_0355_));
 sky130_fd_sc_hd__a22o_1 _0808_ (.A1(_0354_),
    .A2(net5),
    .B1(\rd_addr[21] ),
    .B2(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__a211o_1 _0809_ (.A1(_0352_),
    .A2(net19),
    .B1(_0353_),
    .C1(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__xor2_2 _0810_ (.A(\rd_addr[16] ),
    .B(net8),
    .X(_0358_));
 sky130_fd_sc_hd__o211a_1 _0811_ (.A1(_0352_),
    .A2(net19),
    .B1(net52),
    .C1(rd_valid),
    .X(_0359_));
 sky130_fd_sc_hd__or4b_1 _0812_ (.A(_0351_),
    .B(_0357_),
    .C(_0358_),
    .D_N(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__nor3_2 _0813_ (.A(_0330_),
    .B(_0346_),
    .C(_0360_),
    .Y(net113));
 sky130_fd_sc_hd__clkinv_2 _0814_ (.A(net51),
    .Y(_0361_));
 sky130_fd_sc_hd__or2_1 _0815_ (.A(_0361_),
    .B(softreset),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_4 _0816_ (.A(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__and2_1 _0817_ (.A(\rd_addr[16] ),
    .B(\rd_addr[17] ),
    .X(_0364_));
 sky130_fd_sc_hd__and2_1 _0818_ (.A(\rd_addr[14] ),
    .B(\rd_addr[15] ),
    .X(_0365_));
 sky130_fd_sc_hd__and4_1 _0819_ (.A(\rd_addr[2] ),
    .B(\rd_addr[3] ),
    .C(\rd_addr[4] ),
    .D(\rd_addr[5] ),
    .X(_0366_));
 sky130_fd_sc_hd__and2_1 _0820_ (.A(\rd_addr[6] ),
    .B(\rd_addr[7] ),
    .X(_0367_));
 sky130_fd_sc_hd__and2_1 _0821_ (.A(\rd_addr[8] ),
    .B(\rd_addr[9] ),
    .X(_0368_));
 sky130_fd_sc_hd__and3_1 _0822_ (.A(\rd_addr[10] ),
    .B(\rd_addr[11] ),
    .C(\rd_addr[12] ),
    .X(_0369_));
 sky130_fd_sc_hd__and4_1 _0823_ (.A(_0366_),
    .B(_0367_),
    .C(_0368_),
    .D(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_2 _0824_ (.A(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__and4_1 _0825_ (.A(_0333_),
    .B(_0364_),
    .C(_0365_),
    .D(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__buf_2 _0826_ (.A(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__a31o_1 _0827_ (.A1(\rd_addr[18] ),
    .A2(\rd_addr[19] ),
    .A3(_0373_),
    .B1(\rd_addr[20] ),
    .X(_0374_));
 sky130_fd_sc_hd__and3_1 _0828_ (.A(\rd_addr[18] ),
    .B(\rd_addr[19] ),
    .C(\rd_addr[20] ),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_4 _0829_ (.A(_0366_),
    .X(_0376_));
 sky130_fd_sc_hd__and4_1 _0830_ (.A(\rd_addr[10] ),
    .B(\rd_addr[11] ),
    .C(\rd_addr[12] ),
    .D(_0333_),
    .X(_0377_));
 sky130_fd_sc_hd__and4_1 _0831_ (.A(_0376_),
    .B(_0367_),
    .C(_0368_),
    .D(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__nand4_2 _0832_ (.A(_0375_),
    .B(_0364_),
    .C(_0365_),
    .D(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__and3_1 _0833_ (.A(net13),
    .B(_0374_),
    .C(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__a21oi_1 _0834_ (.A1(_0374_),
    .A2(_0379_),
    .B1(net13),
    .Y(_0381_));
 sky130_fd_sc_hd__and4_1 _0835_ (.A(\rd_addr[21] ),
    .B(\rd_addr[22] ),
    .C(_0375_),
    .D(_0373_),
    .X(_0382_));
 sky130_fd_sc_hd__and4_1 _0836_ (.A(_0333_),
    .B(\rd_addr[16] ),
    .C(_0365_),
    .D(_0371_),
    .X(_0383_));
 sky130_fd_sc_hd__and2_1 _0837_ (.A(_0327_),
    .B(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__nor2_1 _0838_ (.A(_0327_),
    .B(_0383_),
    .Y(_0385_));
 sky130_fd_sc_hd__o2bb2a_1 _0839_ (.A1_N(_0316_),
    .A2_N(_0382_),
    .B1(_0384_),
    .B2(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__and2_1 _0840_ (.A(\rd_addr[18] ),
    .B(_0373_),
    .X(_0387_));
 sky130_fd_sc_hd__xnor2_1 _0841_ (.A(_0333_),
    .B(_0371_),
    .Y(_0388_));
 sky130_fd_sc_hd__xnor2_1 _0842_ (.A(_0334_),
    .B(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__a21oi_1 _0843_ (.A1(\rd_addr[18] ),
    .A2(_0315_),
    .B1(_0350_),
    .Y(_0390_));
 sky130_fd_sc_hd__mux2_1 _0844_ (.A0(_0350_),
    .A1(_0390_),
    .S(_0373_),
    .X(_0391_));
 sky130_fd_sc_hd__and3_1 _0845_ (.A(_0333_),
    .B(\rd_addr[14] ),
    .C(_0371_),
    .X(_0392_));
 sky130_fd_sc_hd__xnor2_1 _0846_ (.A(_0323_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__o2111a_1 _0847_ (.A1(_0315_),
    .A2(_0387_),
    .B1(_0389_),
    .C1(_0391_),
    .D1(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__and3_1 _0848_ (.A(_0333_),
    .B(_0365_),
    .C(_0371_),
    .X(_0395_));
 sky130_fd_sc_hd__xnor2_1 _0849_ (.A(_0358_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__and2_1 _0850_ (.A(_0333_),
    .B(_0371_),
    .X(_0397_));
 sky130_fd_sc_hd__xor2_1 _0851_ (.A(_0328_),
    .B(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__and3_1 _0852_ (.A(\rd_addr[8] ),
    .B(_0366_),
    .C(_0367_),
    .X(_0399_));
 sky130_fd_sc_hd__a21oi_1 _0853_ (.A1(_0376_),
    .A2(_0367_),
    .B1(\rd_addr[8] ),
    .Y(_0400_));
 sky130_fd_sc_hd__o21ai_1 _0854_ (.A1(_0399_),
    .A2(_0400_),
    .B1(net23),
    .Y(_0401_));
 sky130_fd_sc_hd__and3_1 _0855_ (.A(_0376_),
    .B(_0367_),
    .C(_0368_),
    .X(_0402_));
 sky130_fd_sc_hd__xnor2_1 _0856_ (.A(_0314_),
    .B(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__and3_1 _0857_ (.A(\rd_addr[2] ),
    .B(\rd_addr[3] ),
    .C(\rd_addr[4] ),
    .X(_0404_));
 sky130_fd_sc_hd__a21oi_1 _0858_ (.A1(\rd_addr[2] ),
    .A2(\rd_addr[3] ),
    .B1(\rd_addr[4] ),
    .Y(_0405_));
 sky130_fd_sc_hd__o21ai_1 _0859_ (.A1(_0404_),
    .A2(_0405_),
    .B1(net19),
    .Y(_0406_));
 sky130_fd_sc_hd__or3_1 _0860_ (.A(net19),
    .B(_0404_),
    .C(_0405_),
    .X(_0407_));
 sky130_fd_sc_hd__and4_1 _0861_ (.A(_0324_),
    .B(_0345_),
    .C(_0406_),
    .D(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__and3_1 _0862_ (.A(\rd_addr[6] ),
    .B(_0320_),
    .C(_0376_),
    .X(_0409_));
 sky130_fd_sc_hd__a21oi_1 _0863_ (.A1(\rd_addr[6] ),
    .A2(_0376_),
    .B1(_0320_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand3_1 _0864_ (.A(\rd_addr[2] ),
    .B(\rd_addr[3] ),
    .C(\rd_addr[4] ),
    .Y(_0411_));
 sky130_fd_sc_hd__xor2_1 _0865_ (.A(\rd_addr[2] ),
    .B(\rd_addr[3] ),
    .X(_0412_));
 sky130_fd_sc_hd__o2bb2a_1 _0866_ (.A1_N(_0347_),
    .A2_N(_0411_),
    .B1(_0412_),
    .B2(_0336_),
    .X(_0413_));
 sky130_fd_sc_hd__o2bb2a_1 _0867_ (.A1_N(_0336_),
    .A2_N(_0412_),
    .B1(_0347_),
    .B2(_0411_),
    .X(_0414_));
 sky130_fd_sc_hd__xnor2_1 _0868_ (.A(_0318_),
    .B(_0376_),
    .Y(_0415_));
 sky130_fd_sc_hd__o2111a_1 _0869_ (.A1(_0409_),
    .A2(_0410_),
    .B1(_0413_),
    .C1(_0414_),
    .D1(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__and4_1 _0870_ (.A(_0401_),
    .B(_0403_),
    .C(_0408_),
    .D(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__and4_1 _0871_ (.A(\rd_addr[10] ),
    .B(_0366_),
    .C(_0367_),
    .D(_0368_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_2 _0872_ (.A(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__a21oi_1 _0873_ (.A1(\rd_addr[11] ),
    .A2(_0419_),
    .B1(_0348_),
    .Y(_0420_));
 sky130_fd_sc_hd__and3_1 _0874_ (.A(\rd_addr[11] ),
    .B(_0348_),
    .C(_0419_),
    .X(_0421_));
 sky130_fd_sc_hd__xnor2_1 _0875_ (.A(_0319_),
    .B(_0419_),
    .Y(_0422_));
 sky130_fd_sc_hd__or3_1 _0876_ (.A(net23),
    .B(_0399_),
    .C(_0400_),
    .X(_0423_));
 sky130_fd_sc_hd__xnor2_1 _0877_ (.A(_0321_),
    .B(_0399_),
    .Y(_0424_));
 sky130_fd_sc_hd__o2111a_1 _0878_ (.A1(_0420_),
    .A2(_0421_),
    .B1(_0422_),
    .C1(_0423_),
    .D1(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__and4_1 _0879_ (.A(_0396_),
    .B(_0398_),
    .C(_0417_),
    .D(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__o2111a_2 _0880_ (.A1(_0380_),
    .A2(_0381_),
    .B1(_0386_),
    .C1(_0394_),
    .D1(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__xnor2_1 _0881_ (.A(_0338_),
    .B(_0379_),
    .Y(_0428_));
 sky130_fd_sc_hd__xnor2_1 _0882_ (.A(_0355_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__and3_1 _0883_ (.A(\rd_addr[21] ),
    .B(_0375_),
    .C(_0373_),
    .X(_0430_));
 sky130_fd_sc_hd__xor2_1 _0884_ (.A(_0349_),
    .B(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__nand2_1 _0885_ (.A(\rd_addr[23] ),
    .B(_0382_),
    .Y(_0432_));
 sky130_fd_sc_hd__o2111a_1 _0886_ (.A1(_0316_),
    .A2(_0382_),
    .B1(_0429_),
    .C1(_0431_),
    .D1(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__inv_2 _0887_ (.A(net52),
    .Y(_0434_));
 sky130_fd_sc_hd__or3b_2 _0888_ (.A(_0434_),
    .B(net113),
    .C_N(rd_valid),
    .X(_0435_));
 sky130_fd_sc_hd__a21oi_4 _0889_ (.A1(_0427_),
    .A2(_0433_),
    .B1(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__nor2_4 _0890_ (.A(_0363_),
    .B(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__clkbuf_8 _0891_ (.A(\xfer.resetn ),
    .X(_0438_));
 sky130_fd_sc_hd__clkinv_2 _0892_ (.A(\xfer.din_valid ),
    .Y(_0439_));
 sky130_fd_sc_hd__or2_1 _0893_ (.A(\xfer.count[0] ),
    .B(\xfer.count[1] ),
    .X(_0440_));
 sky130_fd_sc_hd__or2b_1 _0894_ (.A(\xfer.xfer_qspi ),
    .B_N(\xfer.flash_clk ),
    .X(_0441_));
 sky130_fd_sc_hd__and2_1 _0895_ (.A(\xfer.count[0] ),
    .B(\xfer.xfer_dspi ),
    .X(_0442_));
 sky130_fd_sc_hd__and2b_1 _0896_ (.A_N(\xfer.xfer_dspi ),
    .B(\xfer.count[1] ),
    .X(_0443_));
 sky130_fd_sc_hd__a2111o_1 _0897_ (.A1(_0440_),
    .A2(_0441_),
    .B1(_0442_),
    .C1(_0443_),
    .D1(\xfer.count[3] ),
    .X(_0444_));
 sky130_fd_sc_hd__nor2_2 _0898_ (.A(\xfer.xfer_dspi ),
    .B(\xfer.xfer_qspi ),
    .Y(_0445_));
 sky130_fd_sc_hd__or4_4 _0899_ (.A(\xfer.dummy_count[3] ),
    .B(\xfer.dummy_count[2] ),
    .C(\xfer.dummy_count[1] ),
    .D(\xfer.dummy_count[0] ),
    .X(_0446_));
 sky130_fd_sc_hd__a21o_1 _0900_ (.A1(\xfer.xfer_ddr ),
    .A2(_0445_),
    .B1(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__inv_2 _0901_ (.A(\xfer.flash_clk ),
    .Y(_0448_));
 sky130_fd_sc_hd__clkinv_2 _0902_ (.A(\xfer.xfer_qspi ),
    .Y(_0449_));
 sky130_fd_sc_hd__nand2_1 _0903_ (.A(\xfer.xfer_ddr ),
    .B(\xfer.xfer_qspi ),
    .Y(_0450_));
 sky130_fd_sc_hd__buf_2 _0904_ (.A(\xfer.count[2] ),
    .X(_0451_));
 sky130_fd_sc_hd__o211a_1 _0905_ (.A1(_0448_),
    .A2(_0449_),
    .B1(_0450_),
    .C1(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__or3_2 _0906_ (.A(_0444_),
    .B(_0447_),
    .C(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__nor2_8 _0907_ (.A(_0439_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__nand2_4 _0908_ (.A(_0438_),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__buf_4 _0909_ (.A(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__a31o_1 _0910_ (.A1(\state[0] ),
    .A2(_0437_),
    .A3(_0456_),
    .B1(_0363_),
    .X(_0000_));
 sky130_fd_sc_hd__inv_2 _0911_ (.A(\xfer.resetn ),
    .Y(_0457_));
 sky130_fd_sc_hd__or2_2 _0912_ (.A(_0451_),
    .B(\xfer.count[3] ),
    .X(_0458_));
 sky130_fd_sc_hd__buf_4 _0913_ (.A(\xfer.flash_clk ),
    .X(_0459_));
 sky130_fd_sc_hd__or4_2 _0914_ (.A(\xfer.count[0] ),
    .B(\xfer.count[2] ),
    .C(\xfer.count[1] ),
    .D(\xfer.count[3] ),
    .X(_0460_));
 sky130_fd_sc_hd__nand2_1 _0915_ (.A(_0459_),
    .B(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__nor2_1 _0916_ (.A(\xfer.count[1] ),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__a21o_1 _0917_ (.A1(_0448_),
    .A2(\xfer.count[1] ),
    .B1(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__nand2_2 _0918_ (.A(\xfer.xfer_dspi ),
    .B(_0449_),
    .Y(_0464_));
 sky130_fd_sc_hd__clkinv_2 _0919_ (.A(\xfer.xfer_ddr ),
    .Y(_0465_));
 sky130_fd_sc_hd__nand2_2 _0920_ (.A(_0465_),
    .B(_0445_),
    .Y(_0466_));
 sky130_fd_sc_hd__a211o_1 _0921_ (.A1(\xfer.count[0] ),
    .A2(_0448_),
    .B1(\xfer.count[1] ),
    .C1(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__o31a_1 _0922_ (.A1(\xfer.count[0] ),
    .A2(_0463_),
    .A3(_0464_),
    .B1(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__nand2_1 _0923_ (.A(_0465_),
    .B(\xfer.xfer_qspi ),
    .Y(_0469_));
 sky130_fd_sc_hd__nor2_1 _0924_ (.A(\xfer.count[0] ),
    .B(\xfer.count[1] ),
    .Y(_0470_));
 sky130_fd_sc_hd__nand2_1 _0925_ (.A(_0451_),
    .B(\xfer.count[3] ),
    .Y(_0471_));
 sky130_fd_sc_hd__o21ai_1 _0926_ (.A1(_0470_),
    .A2(_0458_),
    .B1(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__mux2_1 _0927_ (.A0(\xfer.count[3] ),
    .A1(_0472_),
    .S(_0459_),
    .X(_0473_));
 sky130_fd_sc_hd__nand2_1 _0928_ (.A(_0448_),
    .B(_0451_),
    .Y(_0474_));
 sky130_fd_sc_hd__o21ai_1 _0929_ (.A1(_0451_),
    .A2(_0461_),
    .B1(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__o32a_1 _0930_ (.A1(_0469_),
    .A2(_0473_),
    .A3(_0475_),
    .B1(_0450_),
    .B2(\xfer.count[3] ),
    .X(_0476_));
 sky130_fd_sc_hd__o22a_1 _0931_ (.A1(_0458_),
    .A2(_0468_),
    .B1(_0476_),
    .B2(_0440_),
    .X(_0477_));
 sky130_fd_sc_hd__or4_4 _0932_ (.A(_0439_),
    .B(_0457_),
    .C(_0446_),
    .D(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__nor2_4 _0933_ (.A(_0361_),
    .B(softreset),
    .Y(_0479_));
 sky130_fd_sc_hd__and3b_1 _0934_ (.A_N(_0436_),
    .B(_0478_),
    .C(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__buf_2 _0935_ (.A(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__and2_1 _0936_ (.A(_0438_),
    .B(_0454_),
    .X(_0482_));
 sky130_fd_sc_hd__clkbuf_4 _0937_ (.A(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__and3b_1 _0938_ (.A_N(_0436_),
    .B(_0483_),
    .C(_0479_),
    .X(_0484_));
 sky130_fd_sc_hd__buf_2 _0939_ (.A(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__a22o_1 _0940_ (.A1(\state[5] ),
    .A2(_0481_),
    .B1(_0485_),
    .B2(\state[8] ),
    .X(_0008_));
 sky130_fd_sc_hd__or2_1 _0941_ (.A(config_qspi),
    .B(config_ddr),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_4 _0942_ (.A(\state[1] ),
    .X(_0487_));
 sky130_fd_sc_hd__a32o_1 _0943_ (.A1(\state[12] ),
    .A2(_0485_),
    .A3(_0486_),
    .B1(_0481_),
    .B2(_0487_),
    .X(_0004_));
 sky130_fd_sc_hd__or2_1 _0944_ (.A(\xfer.fetch ),
    .B(\xfer.xfer_ddr_q ),
    .X(_0488_));
 sky130_fd_sc_hd__or4_1 _0945_ (.A(_0444_),
    .B(_0447_),
    .C(_0452_),
    .D(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__nand3b_1 _0946_ (.A_N(\xfer.last_fetch ),
    .B(\xfer.xfer_ddr_q ),
    .C(\xfer.fetch ),
    .Y(_0490_));
 sky130_fd_sc_hd__a21oi_4 _0947_ (.A1(_0489_),
    .A2(_0490_),
    .B1(_0457_),
    .Y(_0491_));
 sky130_fd_sc_hd__a32o_1 _0948_ (.A1(\state[7] ),
    .A2(_0437_),
    .A3(_0491_),
    .B1(_0481_),
    .B2(\state[4] ),
    .X(_0007_));
 sky130_fd_sc_hd__and2_1 _0949_ (.A(_0434_),
    .B(rd_wait),
    .X(_0492_));
 sky130_fd_sc_hd__or2_1 _0950_ (.A(_0455_),
    .B(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__a22o_1 _0951_ (.A1(\state[11] ),
    .A2(_0483_),
    .B1(_0493_),
    .B2(\state[3] ),
    .X(_0494_));
 sky130_fd_sc_hd__and2_1 _0952_ (.A(_0437_),
    .B(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_1 _0953_ (.A(_0495_),
    .X(_0006_));
 sky130_fd_sc_hd__nand2_1 _0954_ (.A(\state[10] ),
    .B(_0491_),
    .Y(_0496_));
 sky130_fd_sc_hd__a211o_2 _0955_ (.A1(_0427_),
    .A2(_0433_),
    .B1(config_cont),
    .C1(_0435_),
    .X(_0497_));
 sky130_fd_sc_hd__o21a_1 _0956_ (.A1(_0436_),
    .A2(_0496_),
    .B1(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_4 _0957_ (.A(\state[2] ),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_4 _0958_ (.A(_0479_),
    .X(_0500_));
 sky130_fd_sc_hd__and4b_1 _0959_ (.A_N(_0436_),
    .B(_0456_),
    .C(_0499_),
    .D(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__o21bai_1 _0960_ (.A1(_0363_),
    .A2(_0498_),
    .B1_N(_0501_),
    .Y(_0005_));
 sky130_fd_sc_hd__a22o_1 _0961_ (.A1(\state[11] ),
    .A2(_0481_),
    .B1(_0485_),
    .B2(\state[5] ),
    .X(_0002_));
 sky130_fd_sc_hd__inv_2 _0962_ (.A(_0491_),
    .Y(_0502_));
 sky130_fd_sc_hd__a32o_1 _0963_ (.A1(\state[10] ),
    .A2(_0437_),
    .A3(_0502_),
    .B1(_0485_),
    .B2(\state[4] ),
    .X(_0001_));
 sky130_fd_sc_hd__clkbuf_4 _0964_ (.A(\state[9] ),
    .X(_0503_));
 sky130_fd_sc_hd__or4_1 _0965_ (.A(_0319_),
    .B(_0320_),
    .C(_0323_),
    .D(_0358_),
    .X(_0504_));
 sky130_fd_sc_hd__nor4_1 _0966_ (.A(_0318_),
    .B(_0347_),
    .C(_0348_),
    .D(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__a2111oi_1 _0967_ (.A1(_0338_),
    .A2(net14),
    .B1(_0331_),
    .C1(_0340_),
    .D1(_0353_),
    .Y(_0506_));
 sky130_fd_sc_hd__inv_2 _0968_ (.A(net2),
    .Y(_0507_));
 sky130_fd_sc_hd__o221a_1 _0969_ (.A1(\rd_addr[10] ),
    .A2(_0507_),
    .B1(\rd_addr[20] ),
    .B2(_0332_),
    .C1(_0326_),
    .X(_0508_));
 sky130_fd_sc_hd__o221a_1 _0970_ (.A1(\rd_addr[3] ),
    .A2(_0336_),
    .B1(_0338_),
    .B2(net14),
    .C1(_0325_),
    .X(_0509_));
 sky130_fd_sc_hd__and4_1 _0971_ (.A(_0345_),
    .B(_0506_),
    .C(_0508_),
    .D(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__xnor2_1 _0972_ (.A(\rd_addr[4] ),
    .B(net19),
    .Y(_0511_));
 sky130_fd_sc_hd__o2111a_1 _0973_ (.A1(_0333_),
    .A2(_0334_),
    .B1(_0511_),
    .C1(rd_valid),
    .D1(net52),
    .X(_0512_));
 sky130_fd_sc_hd__o221a_1 _0974_ (.A1(_0337_),
    .A2(net18),
    .B1(_0354_),
    .B2(net5),
    .C1(_0350_),
    .X(_0513_));
 sky130_fd_sc_hd__inv_2 _0975_ (.A(\rd_addr[10] ),
    .Y(_0514_));
 sky130_fd_sc_hd__o211a_1 _0976_ (.A1(_0514_),
    .A2(net2),
    .B1(_0328_),
    .C1(_0349_),
    .X(_0515_));
 sky130_fd_sc_hd__xor2_1 _0977_ (.A(\rd_addr[23] ),
    .B(net16),
    .X(_0516_));
 sky130_fd_sc_hd__nor4b_1 _0978_ (.A(_0516_),
    .B(_0321_),
    .C(_0324_),
    .D_N(_0315_),
    .Y(_0517_));
 sky130_fd_sc_hd__and4_1 _0979_ (.A(_0512_),
    .B(_0513_),
    .C(_0515_),
    .D(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__a31o_1 _0980_ (.A1(_0505_),
    .A2(_0510_),
    .A3(_0518_),
    .B1(_0434_),
    .X(_0519_));
 sky130_fd_sc_hd__and2_1 _0981_ (.A(\state[9] ),
    .B(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__o211a_1 _0982_ (.A1(_0436_),
    .A2(_0520_),
    .B1(_0497_),
    .C1(_0500_),
    .X(_0521_));
 sky130_fd_sc_hd__a221o_1 _0983_ (.A1(_0503_),
    .A2(_0481_),
    .B1(_0485_),
    .B2(_0499_),
    .C1(_0521_),
    .X(_0012_));
 sky130_fd_sc_hd__buf_4 _0984_ (.A(config_ddr),
    .X(_0522_));
 sky130_fd_sc_hd__nor2_1 _0985_ (.A(config_qspi),
    .B(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__and2b_1 _0986_ (.A_N(_0492_),
    .B(\state[3] ),
    .X(_0524_));
 sky130_fd_sc_hd__a211o_1 _0987_ (.A1(\state[12] ),
    .A2(_0523_),
    .B1(_0524_),
    .C1(_0487_),
    .X(_0525_));
 sky130_fd_sc_hd__a22o_1 _0988_ (.A1(\state[8] ),
    .A2(_0481_),
    .B1(_0485_),
    .B2(_0525_),
    .X(_0011_));
 sky130_fd_sc_hd__buf_4 _0989_ (.A(_0483_),
    .X(_0526_));
 sky130_fd_sc_hd__and4b_1 _0990_ (.A_N(_0436_),
    .B(_0502_),
    .C(\state[7] ),
    .D(_0500_),
    .X(_0527_));
 sky130_fd_sc_hd__a31o_1 _0991_ (.A1(\state[0] ),
    .A2(_0437_),
    .A3(_0526_),
    .B1(_0527_),
    .X(_0010_));
 sky130_fd_sc_hd__clkbuf_4 _0992_ (.A(\state[6] ),
    .X(_0528_));
 sky130_fd_sc_hd__inv_2 _0993_ (.A(_0503_),
    .Y(_0529_));
 sky130_fd_sc_hd__nor2_2 _0994_ (.A(_0529_),
    .B(_0519_),
    .Y(_0530_));
 sky130_fd_sc_hd__a22o_1 _0995_ (.A1(_0528_),
    .A2(_0481_),
    .B1(_0485_),
    .B2(_0530_),
    .X(_0009_));
 sky130_fd_sc_hd__a22o_1 _0996_ (.A1(\state[12] ),
    .A2(_0481_),
    .B1(_0485_),
    .B2(_0528_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _0997_ (.A0(config_csb),
    .A1(\xfer.flash_csb ),
    .S(config_en),
    .X(_0531_));
 sky130_fd_sc_hd__buf_6 _0998_ (.A(_0531_),
    .X(net72));
 sky130_fd_sc_hd__mux2_1 _0999_ (.A0(config_clk),
    .A1(_0459_),
    .S(config_en),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_8 _1000_ (.A(_0532_),
    .X(net71));
 sky130_fd_sc_hd__nor4_4 _1001_ (.A(\xfer.dummy_count[3] ),
    .B(\xfer.dummy_count[2] ),
    .C(\xfer.dummy_count[1] ),
    .D(\xfer.dummy_count[0] ),
    .Y(_0533_));
 sky130_fd_sc_hd__and2_2 _1002_ (.A(_0465_),
    .B(_0445_),
    .X(_0534_));
 sky130_fd_sc_hd__buf_4 _1003_ (.A(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__buf_4 _1004_ (.A(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__clkinv_2 _1005_ (.A(config_en),
    .Y(_0537_));
 sky130_fd_sc_hd__or2_1 _1006_ (.A(_0446_),
    .B(_0445_),
    .X(_0538_));
 sky130_fd_sc_hd__or3_1 _1007_ (.A(\xfer.xfer_rd ),
    .B(_0537_),
    .C(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__a21bo_1 _1008_ (.A1(\config_oe[0] ),
    .A2(_0537_),
    .B1_N(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__a31o_4 _1009_ (.A1(config_en),
    .A2(_0533_),
    .A3(_0536_),
    .B1(_0540_),
    .X(net74));
 sky130_fd_sc_hd__a21bo_4 _1010_ (.A1(\config_oe[1] ),
    .A2(_0537_),
    .B1_N(_0539_),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 _1011_ (.A(\xfer.xfer_qspi ),
    .X(_0541_));
 sky130_fd_sc_hd__buf_4 _1012_ (.A(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__and4b_1 _1013_ (.A_N(\xfer.xfer_rd ),
    .B(config_en),
    .C(_0533_),
    .D(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__a21o_4 _1014_ (.A1(\config_oe[2] ),
    .A2(_0537_),
    .B1(_0543_),
    .X(net78));
 sky130_fd_sc_hd__a21o_4 _1015_ (.A1(\config_oe[3] ),
    .A2(_0537_),
    .B1(_0543_),
    .X(net80));
 sky130_fd_sc_hd__a21oi_1 _1016_ (.A1(\xfer.xfer_ddr ),
    .A2(_0445_),
    .B1(_0446_),
    .Y(_0544_));
 sky130_fd_sc_hd__o221a_1 _1017_ (.A1(_0449_),
    .A2(\xfer.obuffer[4] ),
    .B1(_0464_),
    .B2(\xfer.obuffer[6] ),
    .C1(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__o21a_1 _1018_ (.A1(\xfer.obuffer[7] ),
    .A2(_0466_),
    .B1(_0545_),
    .X(\xfer.flash_io0_do ));
 sky130_fd_sc_hd__mux2_1 _1019_ (.A0(\xfer.flash_io0_do ),
    .A1(xfer_io0_90),
    .S(_0522_),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_4 _1020_ (.A0(\config_do[0] ),
    .A1(_0546_),
    .S(config_en),
    .X(_0547_));
 sky130_fd_sc_hd__clkbuf_1 _1021_ (.A(_0547_),
    .X(net73));
 sky130_fd_sc_hd__inv_2 _1022_ (.A(_0538_),
    .Y(_0548_));
 sky130_fd_sc_hd__o221a_1 _1023_ (.A1(_0449_),
    .A2(\xfer.obuffer[5] ),
    .B1(_0464_),
    .B2(\xfer.obuffer[7] ),
    .C1(_0548_),
    .X(\xfer.flash_io1_do ));
 sky130_fd_sc_hd__mux2_1 _1024_ (.A0(\xfer.flash_io1_do ),
    .A1(xfer_io1_90),
    .S(_0522_),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_2 _1025_ (.A0(\config_do[1] ),
    .A1(_0549_),
    .S(config_en),
    .X(_0550_));
 sky130_fd_sc_hd__clkbuf_2 _1026_ (.A(_0550_),
    .X(net75));
 sky130_fd_sc_hd__and3_1 _1027_ (.A(_0541_),
    .B(\xfer.obuffer[6] ),
    .C(_0533_),
    .X(_0551_));
 sky130_fd_sc_hd__clkbuf_1 _1028_ (.A(_0551_),
    .X(\xfer.flash_io2_do ));
 sky130_fd_sc_hd__mux2_1 _1029_ (.A0(\xfer.flash_io2_do ),
    .A1(xfer_io2_90),
    .S(_0522_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_4 _1030_ (.A0(\config_do[2] ),
    .A1(_0552_),
    .S(config_en),
    .X(_0553_));
 sky130_fd_sc_hd__clkbuf_1 _1031_ (.A(_0553_),
    .X(net77));
 sky130_fd_sc_hd__and3_1 _1032_ (.A(_0541_),
    .B(\xfer.obuffer[7] ),
    .C(_0533_),
    .X(_0554_));
 sky130_fd_sc_hd__clkbuf_1 _1033_ (.A(_0554_),
    .X(\xfer.flash_io3_do ));
 sky130_fd_sc_hd__mux2_1 _1034_ (.A0(\xfer.flash_io3_do ),
    .A1(xfer_io3_90),
    .S(_0522_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_4 _1035_ (.A0(\config_do[3] ),
    .A1(_0555_),
    .S(config_en),
    .X(_0556_));
 sky130_fd_sc_hd__clkbuf_1 _1036_ (.A(_0556_),
    .X(net79));
 sky130_fd_sc_hd__and2b_1 _1037_ (.A_N(\xfer.dout_tag[0] ),
    .B(_0491_),
    .X(_0557_));
 sky130_fd_sc_hd__and3b_1 _1038_ (.A_N(\xfer.dout_tag[2] ),
    .B(_0479_),
    .C(\xfer.dout_tag[1] ),
    .X(_0558_));
 sky130_fd_sc_hd__nand2_4 _1039_ (.A(_0557_),
    .B(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__mux2_1 _1040_ (.A0(\xfer.dout_data[0] ),
    .A1(\buffer[8] ),
    .S(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__clkbuf_1 _1041_ (.A(_0560_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _1042_ (.A0(\xfer.dout_data[1] ),
    .A1(\buffer[9] ),
    .S(_0559_),
    .X(_0561_));
 sky130_fd_sc_hd__clkbuf_1 _1043_ (.A(_0561_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _1044_ (.A0(\xfer.dout_data[2] ),
    .A1(\buffer[10] ),
    .S(_0559_),
    .X(_0562_));
 sky130_fd_sc_hd__clkbuf_1 _1045_ (.A(_0562_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _1046_ (.A0(\xfer.dout_data[3] ),
    .A1(\buffer[11] ),
    .S(_0559_),
    .X(_0563_));
 sky130_fd_sc_hd__clkbuf_1 _1047_ (.A(_0563_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _1048_ (.A0(\xfer.dout_data[4] ),
    .A1(\buffer[12] ),
    .S(_0559_),
    .X(_0564_));
 sky130_fd_sc_hd__clkbuf_1 _1049_ (.A(_0564_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _1050_ (.A0(\xfer.dout_data[5] ),
    .A1(\buffer[13] ),
    .S(_0559_),
    .X(_0565_));
 sky130_fd_sc_hd__clkbuf_1 _1051_ (.A(_0565_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _1052_ (.A0(\xfer.dout_data[6] ),
    .A1(\buffer[14] ),
    .S(_0559_),
    .X(_0566_));
 sky130_fd_sc_hd__clkbuf_1 _1053_ (.A(_0566_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _1054_ (.A0(\xfer.dout_data[7] ),
    .A1(\buffer[15] ),
    .S(_0559_),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_1 _1055_ (.A(_0567_),
    .X(_0024_));
 sky130_fd_sc_hd__nor2_2 _1056_ (.A(_0440_),
    .B(_0458_),
    .Y(_0568_));
 sky130_fd_sc_hd__nor2_4 _1057_ (.A(_0447_),
    .B(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__a211o_1 _1058_ (.A1(\xfer.xfer_ddr ),
    .A2(_0464_),
    .B1(_0568_),
    .C1(_0459_),
    .X(_0570_));
 sky130_fd_sc_hd__o211ai_4 _1059_ (.A1(_0454_),
    .A2(_0569_),
    .B1(_0570_),
    .C1(_0438_),
    .Y(_0571_));
 sky130_fd_sc_hd__a22o_1 _1060_ (.A1(\xfer.din_data[0] ),
    .A2(_0526_),
    .B1(_0571_),
    .B2(\xfer.obuffer[0] ),
    .X(_0025_));
 sky130_fd_sc_hd__and3_1 _1061_ (.A(\xfer.dout_tag[0] ),
    .B(_0491_),
    .C(_0558_),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_4 _1062_ (.A(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _1063_ (.A0(\buffer[16] ),
    .A1(\xfer.dout_data[0] ),
    .S(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__clkbuf_1 _1064_ (.A(_0574_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _1065_ (.A0(\buffer[17] ),
    .A1(\xfer.dout_data[1] ),
    .S(_0573_),
    .X(_0575_));
 sky130_fd_sc_hd__clkbuf_1 _1066_ (.A(_0575_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _1067_ (.A0(\buffer[18] ),
    .A1(\xfer.dout_data[2] ),
    .S(_0573_),
    .X(_0576_));
 sky130_fd_sc_hd__clkbuf_1 _1068_ (.A(_0576_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _1069_ (.A0(\buffer[19] ),
    .A1(\xfer.dout_data[3] ),
    .S(_0573_),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_1 _1070_ (.A(_0577_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _1071_ (.A0(\buffer[20] ),
    .A1(\xfer.dout_data[4] ),
    .S(_0573_),
    .X(_0578_));
 sky130_fd_sc_hd__clkbuf_1 _1072_ (.A(_0578_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _1073_ (.A0(\buffer[21] ),
    .A1(\xfer.dout_data[5] ),
    .S(_0573_),
    .X(_0579_));
 sky130_fd_sc_hd__clkbuf_1 _1074_ (.A(_0579_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _1075_ (.A0(\buffer[22] ),
    .A1(\xfer.dout_data[6] ),
    .S(_0573_),
    .X(_0580_));
 sky130_fd_sc_hd__clkbuf_1 _1076_ (.A(_0580_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _1077_ (.A0(\buffer[23] ),
    .A1(\xfer.dout_data[7] ),
    .S(_0573_),
    .X(_0581_));
 sky130_fd_sc_hd__clkbuf_1 _1078_ (.A(_0581_),
    .X(_0033_));
 sky130_fd_sc_hd__a21o_1 _1079_ (.A1(\xfer.obuffer[0] ),
    .A2(_0536_),
    .B1(_0482_),
    .X(_0582_));
 sky130_fd_sc_hd__o21a_1 _1080_ (.A1(\xfer.din_data[1] ),
    .A2(_0456_),
    .B1(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _1081_ (.A0(_0583_),
    .A1(\xfer.obuffer[1] ),
    .S(_0571_),
    .X(_0584_));
 sky130_fd_sc_hd__clkbuf_1 _1082_ (.A(_0584_),
    .X(_0034_));
 sky130_fd_sc_hd__nor2_4 _1083_ (.A(_0541_),
    .B(_0534_),
    .Y(_0585_));
 sky130_fd_sc_hd__a22o_1 _1084_ (.A1(\xfer.obuffer[1] ),
    .A2(_0535_),
    .B1(_0585_),
    .B2(\xfer.obuffer[0] ),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _1085_ (.A0(\xfer.din_data[2] ),
    .A1(_0586_),
    .S(_0456_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _1086_ (.A0(_0587_),
    .A1(\xfer.obuffer[2] ),
    .S(_0571_),
    .X(_0588_));
 sky130_fd_sc_hd__clkbuf_1 _1087_ (.A(_0588_),
    .X(_0035_));
 sky130_fd_sc_hd__a22o_1 _1088_ (.A1(\xfer.obuffer[2] ),
    .A2(_0535_),
    .B1(_0585_),
    .B2(\xfer.obuffer[1] ),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _1089_ (.A0(\xfer.din_data[3] ),
    .A1(_0589_),
    .S(_0456_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _1090_ (.A0(_0590_),
    .A1(\xfer.obuffer[3] ),
    .S(_0571_),
    .X(_0591_));
 sky130_fd_sc_hd__clkbuf_1 _1091_ (.A(_0591_),
    .X(_0036_));
 sky130_fd_sc_hd__buf_4 _1092_ (.A(_0585_),
    .X(_0592_));
 sky130_fd_sc_hd__a22o_1 _1093_ (.A1(_0541_),
    .A2(\xfer.obuffer[0] ),
    .B1(\xfer.obuffer[3] ),
    .B2(_0534_),
    .X(_0593_));
 sky130_fd_sc_hd__a21o_1 _1094_ (.A1(\xfer.obuffer[2] ),
    .A2(_0592_),
    .B1(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _1095_ (.A0(\xfer.din_data[4] ),
    .A1(_0594_),
    .S(_0455_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _1096_ (.A0(_0595_),
    .A1(\xfer.obuffer[4] ),
    .S(_0571_),
    .X(_0596_));
 sky130_fd_sc_hd__clkbuf_1 _1097_ (.A(_0596_),
    .X(_0037_));
 sky130_fd_sc_hd__a22o_1 _1098_ (.A1(_0541_),
    .A2(\xfer.obuffer[1] ),
    .B1(_0535_),
    .B2(\xfer.obuffer[4] ),
    .X(_0597_));
 sky130_fd_sc_hd__a21o_1 _1099_ (.A1(\xfer.obuffer[3] ),
    .A2(_0592_),
    .B1(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _1100_ (.A0(\xfer.din_data[5] ),
    .A1(_0598_),
    .S(_0455_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _1101_ (.A0(_0599_),
    .A1(\xfer.obuffer[5] ),
    .S(_0571_),
    .X(_0600_));
 sky130_fd_sc_hd__clkbuf_1 _1102_ (.A(_0600_),
    .X(_0038_));
 sky130_fd_sc_hd__a22o_1 _1103_ (.A1(_0541_),
    .A2(\xfer.obuffer[2] ),
    .B1(_0535_),
    .B2(\xfer.obuffer[5] ),
    .X(_0601_));
 sky130_fd_sc_hd__a21o_1 _1104_ (.A1(\xfer.obuffer[4] ),
    .A2(_0592_),
    .B1(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _1105_ (.A0(\xfer.din_data[6] ),
    .A1(_0602_),
    .S(_0455_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _1106_ (.A0(_0603_),
    .A1(\xfer.obuffer[6] ),
    .S(_0571_),
    .X(_0604_));
 sky130_fd_sc_hd__clkbuf_1 _1107_ (.A(_0604_),
    .X(_0039_));
 sky130_fd_sc_hd__a22o_1 _1108_ (.A1(_0541_),
    .A2(\xfer.obuffer[3] ),
    .B1(_0585_),
    .B2(\xfer.obuffer[5] ),
    .X(_0605_));
 sky130_fd_sc_hd__a211o_1 _1109_ (.A1(\xfer.obuffer[6] ),
    .A2(_0535_),
    .B1(_0482_),
    .C1(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__o21a_1 _1110_ (.A1(\xfer.din_data[7] ),
    .A2(_0456_),
    .B1(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _1111_ (.A0(_0607_),
    .A1(\xfer.obuffer[7] ),
    .S(_0571_),
    .X(_0608_));
 sky130_fd_sc_hd__clkbuf_1 _1112_ (.A(_0608_),
    .X(_0040_));
 sky130_fd_sc_hd__nor2_1 _1113_ (.A(_0446_),
    .B(_0460_),
    .Y(_0609_));
 sky130_fd_sc_hd__and3_1 _1114_ (.A(_0459_),
    .B(_0470_),
    .C(_0458_),
    .X(_0610_));
 sky130_fd_sc_hd__and2b_1 _1115_ (.A_N(_0451_),
    .B(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__or3_1 _1116_ (.A(_0451_),
    .B(\xfer.count[1] ),
    .C(_0461_),
    .X(_0612_));
 sky130_fd_sc_hd__nand2_1 _1117_ (.A(_0592_),
    .B(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__o21ai_1 _1118_ (.A1(_0466_),
    .A2(_0611_),
    .B1(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__and3_1 _1119_ (.A(\xfer.xfer_ddr ),
    .B(_0542_),
    .C(_0472_),
    .X(_0615_));
 sky130_fd_sc_hd__and4_1 _1120_ (.A(\xfer.xfer_ddr ),
    .B(_0533_),
    .C(_0445_),
    .D(_0460_),
    .X(_0616_));
 sky130_fd_sc_hd__nor3b_1 _1121_ (.A(_0612_),
    .B(\xfer.count[3] ),
    .C_N(_0585_),
    .Y(_0617_));
 sky130_fd_sc_hd__a311o_1 _1122_ (.A1(_0465_),
    .A2(_0541_),
    .A3(_0473_),
    .B1(_0616_),
    .C1(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__a211o_1 _1123_ (.A1(\xfer.count[3] ),
    .A2(_0614_),
    .B1(_0615_),
    .C1(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__o21a_1 _1124_ (.A1(_0446_),
    .A2(_0454_),
    .B1(_0438_),
    .X(_0620_));
 sky130_fd_sc_hd__a21o_1 _1125_ (.A1(_0438_),
    .A2(_0619_),
    .B1(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__o31a_1 _1126_ (.A1(\xfer.count[3] ),
    .A2(_0544_),
    .A3(_0609_),
    .B1(_0621_),
    .X(_0041_));
 sky130_fd_sc_hd__or3_1 _1127_ (.A(_0465_),
    .B(_0457_),
    .C(\xfer.fetch ),
    .X(_0622_));
 sky130_fd_sc_hd__clkbuf_1 _1128_ (.A(_0622_),
    .X(_0042_));
 sky130_fd_sc_hd__and4b_1 _1129_ (.A_N(\xfer.dout_tag[1] ),
    .B(\xfer.dout_tag[2] ),
    .C(_0479_),
    .D(_0557_),
    .X(_0623_));
 sky130_fd_sc_hd__buf_4 _1130_ (.A(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _1131_ (.A0(net81),
    .A1(\buffer[0] ),
    .S(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__clkbuf_1 _1132_ (.A(_0625_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _1133_ (.A0(net92),
    .A1(\buffer[1] ),
    .S(_0624_),
    .X(_0626_));
 sky130_fd_sc_hd__clkbuf_1 _1134_ (.A(_0626_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _1135_ (.A0(net103),
    .A1(\buffer[2] ),
    .S(_0624_),
    .X(_0627_));
 sky130_fd_sc_hd__clkbuf_1 _1136_ (.A(_0627_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _1137_ (.A0(net106),
    .A1(\buffer[3] ),
    .S(_0624_),
    .X(_0628_));
 sky130_fd_sc_hd__clkbuf_1 _1138_ (.A(_0628_),
    .X(_0046_));
 sky130_fd_sc_hd__clkbuf_8 _1139_ (.A(_0623_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _1140_ (.A0(net107),
    .A1(\buffer[4] ),
    .S(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__clkbuf_1 _1141_ (.A(_0630_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _1142_ (.A0(net108),
    .A1(\buffer[5] ),
    .S(_0629_),
    .X(_0631_));
 sky130_fd_sc_hd__clkbuf_1 _1143_ (.A(_0631_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _1144_ (.A0(net109),
    .A1(\buffer[6] ),
    .S(_0629_),
    .X(_0632_));
 sky130_fd_sc_hd__clkbuf_1 _1145_ (.A(_0632_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _1146_ (.A0(net110),
    .A1(\buffer[7] ),
    .S(_0629_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_1 _1147_ (.A(_0633_),
    .X(_0050_));
 sky130_fd_sc_hd__or4bb_1 _1148_ (.A(_0363_),
    .B(\xfer.dout_tag[1] ),
    .C_N(\xfer.dout_tag[2] ),
    .D_N(_0557_),
    .X(_0634_));
 sky130_fd_sc_hd__clkbuf_4 _1149_ (.A(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__buf_4 _1150_ (.A(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _1151_ (.A0(\buffer[8] ),
    .A1(net111),
    .S(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__clkbuf_1 _1152_ (.A(_0637_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _1153_ (.A0(\buffer[9] ),
    .A1(net112),
    .S(_0636_),
    .X(_0638_));
 sky130_fd_sc_hd__clkbuf_1 _1154_ (.A(_0638_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _1155_ (.A0(\buffer[10] ),
    .A1(net82),
    .S(_0636_),
    .X(_0639_));
 sky130_fd_sc_hd__clkbuf_1 _1156_ (.A(_0639_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _1157_ (.A0(\buffer[11] ),
    .A1(net83),
    .S(_0636_),
    .X(_0640_));
 sky130_fd_sc_hd__clkbuf_1 _1158_ (.A(_0640_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _1159_ (.A0(\buffer[12] ),
    .A1(net84),
    .S(_0636_),
    .X(_0641_));
 sky130_fd_sc_hd__clkbuf_1 _1160_ (.A(_0641_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _1161_ (.A0(\buffer[13] ),
    .A1(net85),
    .S(_0636_),
    .X(_0642_));
 sky130_fd_sc_hd__clkbuf_1 _1162_ (.A(_0642_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _1163_ (.A0(\buffer[14] ),
    .A1(net86),
    .S(_0636_),
    .X(_0643_));
 sky130_fd_sc_hd__clkbuf_1 _1164_ (.A(_0643_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _1165_ (.A0(\buffer[15] ),
    .A1(net87),
    .S(_0636_),
    .X(_0644_));
 sky130_fd_sc_hd__clkbuf_1 _1166_ (.A(_0644_),
    .X(_0058_));
 sky130_fd_sc_hd__buf_4 _1167_ (.A(_0635_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _1168_ (.A0(\buffer[16] ),
    .A1(net88),
    .S(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__clkbuf_1 _1169_ (.A(_0646_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _1170_ (.A0(\buffer[17] ),
    .A1(net89),
    .S(_0645_),
    .X(_0647_));
 sky130_fd_sc_hd__clkbuf_1 _1171_ (.A(_0647_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1172_ (.A0(\buffer[18] ),
    .A1(net90),
    .S(_0645_),
    .X(_0648_));
 sky130_fd_sc_hd__clkbuf_1 _1173_ (.A(_0648_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1174_ (.A0(\buffer[19] ),
    .A1(net91),
    .S(_0645_),
    .X(_0649_));
 sky130_fd_sc_hd__clkbuf_1 _1175_ (.A(_0649_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1176_ (.A0(\buffer[20] ),
    .A1(net93),
    .S(_0645_),
    .X(_0650_));
 sky130_fd_sc_hd__clkbuf_1 _1177_ (.A(_0650_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1178_ (.A0(\buffer[21] ),
    .A1(net94),
    .S(_0645_),
    .X(_0651_));
 sky130_fd_sc_hd__clkbuf_1 _1179_ (.A(_0651_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1180_ (.A0(\buffer[22] ),
    .A1(net95),
    .S(_0645_),
    .X(_0652_));
 sky130_fd_sc_hd__clkbuf_1 _1181_ (.A(_0652_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1182_ (.A0(\buffer[23] ),
    .A1(net96),
    .S(_0645_),
    .X(_0653_));
 sky130_fd_sc_hd__clkbuf_1 _1183_ (.A(_0653_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1184_ (.A0(\xfer.dout_data[0] ),
    .A1(net97),
    .S(_0645_),
    .X(_0654_));
 sky130_fd_sc_hd__clkbuf_1 _1185_ (.A(_0654_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1186_ (.A0(\xfer.dout_data[1] ),
    .A1(net98),
    .S(_0645_),
    .X(_0655_));
 sky130_fd_sc_hd__clkbuf_1 _1187_ (.A(_0655_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1188_ (.A0(\xfer.dout_data[2] ),
    .A1(net99),
    .S(_0635_),
    .X(_0656_));
 sky130_fd_sc_hd__clkbuf_1 _1189_ (.A(_0656_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1190_ (.A0(\xfer.dout_data[3] ),
    .A1(net100),
    .S(_0635_),
    .X(_0657_));
 sky130_fd_sc_hd__clkbuf_1 _1191_ (.A(_0657_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1192_ (.A0(\xfer.dout_data[4] ),
    .A1(net101),
    .S(_0635_),
    .X(_0658_));
 sky130_fd_sc_hd__clkbuf_1 _1193_ (.A(_0658_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1194_ (.A0(\xfer.dout_data[5] ),
    .A1(net102),
    .S(_0635_),
    .X(_0659_));
 sky130_fd_sc_hd__clkbuf_1 _1195_ (.A(_0659_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1196_ (.A0(\xfer.dout_data[6] ),
    .A1(net104),
    .S(_0635_),
    .X(_0660_));
 sky130_fd_sc_hd__clkbuf_1 _1197_ (.A(_0660_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1198_ (.A0(\xfer.dout_data[7] ),
    .A1(net105),
    .S(_0635_),
    .X(_0661_));
 sky130_fd_sc_hd__clkbuf_1 _1199_ (.A(_0661_),
    .X(_0074_));
 sky130_fd_sc_hd__inv_2 _1200_ (.A(\state[7] ),
    .Y(_0662_));
 sky130_fd_sc_hd__o211a_1 _1201_ (.A1(_0662_),
    .A2(_0502_),
    .B1(_0496_),
    .C1(_0437_),
    .X(_0075_));
 sky130_fd_sc_hd__or4_1 _1202_ (.A(\state[5] ),
    .B(\state[2] ),
    .C(\state[4] ),
    .D(\state[6] ),
    .X(_0663_));
 sky130_fd_sc_hd__or3_1 _1203_ (.A(\state[8] ),
    .B(\state[12] ),
    .C(\state[11] ),
    .X(_0664_));
 sky130_fd_sc_hd__or4_1 _1204_ (.A(\state[0] ),
    .B(\state[1] ),
    .C(_0663_),
    .D(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__or3b_1 _1205_ (.A(_0665_),
    .B(_0524_),
    .C_N(_0519_),
    .X(_0666_));
 sky130_fd_sc_hd__or3_1 _1206_ (.A(\state[3] ),
    .B(\state[9] ),
    .C(_0665_),
    .X(_0667_));
 sky130_fd_sc_hd__and4_1 _1207_ (.A(_0500_),
    .B(_0456_),
    .C(_0666_),
    .D(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__clkbuf_1 _1208_ (.A(_0668_),
    .X(_0076_));
 sky130_fd_sc_hd__nor2_4 _1209_ (.A(_0457_),
    .B(_0454_),
    .Y(_0669_));
 sky130_fd_sc_hd__a22o_1 _1210_ (.A1(\xfer.din_tag[0] ),
    .A2(_0526_),
    .B1(_0669_),
    .B2(\xfer.xfer_tag[0] ),
    .X(_0077_));
 sky130_fd_sc_hd__a22o_1 _1211_ (.A1(\xfer.din_tag[1] ),
    .A2(_0526_),
    .B1(_0669_),
    .B2(\xfer.xfer_tag[1] ),
    .X(_0078_));
 sky130_fd_sc_hd__a22o_1 _1212_ (.A1(\xfer.din_tag[2] ),
    .A2(_0526_),
    .B1(_0669_),
    .B2(\xfer.xfer_tag[2] ),
    .X(_0079_));
 sky130_fd_sc_hd__or2_2 _1213_ (.A(_0363_),
    .B(_0520_),
    .X(_0670_));
 sky130_fd_sc_hd__inv_2 _1214_ (.A(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__nor4_1 _1215_ (.A(_0487_),
    .B(\state[12] ),
    .C(\state[9] ),
    .D(_0663_),
    .Y(_0672_));
 sky130_fd_sc_hd__or2_2 _1216_ (.A(_0670_),
    .B(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__a21bo_2 _1217_ (.A1(\state[0] ),
    .A2(_0671_),
    .B1_N(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__and2_2 _1218_ (.A(\state[12] ),
    .B(_0455_),
    .X(_0675_));
 sky130_fd_sc_hd__a211o_1 _1219_ (.A1(net56),
    .A2(_0487_),
    .B1(\state[4] ),
    .C1(_0499_),
    .X(_0676_));
 sky130_fd_sc_hd__a22o_1 _1220_ (.A1(net8),
    .A2(_0503_),
    .B1(_0528_),
    .B2(net23),
    .X(_0677_));
 sky130_fd_sc_hd__or2_1 _1221_ (.A(_0676_),
    .B(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__and2_1 _1222_ (.A(_0487_),
    .B(_0455_),
    .X(_0679_));
 sky130_fd_sc_hd__a211o_1 _1223_ (.A1(net1),
    .A2(_0675_),
    .B1(_0678_),
    .C1(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__o22a_1 _1224_ (.A1(\xfer.din_data[0] ),
    .A2(_0674_),
    .B1(_0680_),
    .B2(_0673_),
    .X(_0080_));
 sky130_fd_sc_hd__a21boi_1 _1225_ (.A1(config_qspi),
    .A2(_0522_),
    .B1_N(_0499_),
    .Y(_0681_));
 sky130_fd_sc_hd__a221o_1 _1226_ (.A1(net9),
    .A2(_0503_),
    .B1(_0528_),
    .B2(net24),
    .C1(\state[4] ),
    .X(_0682_));
 sky130_fd_sc_hd__a211o_1 _1227_ (.A1(net12),
    .A2(_0675_),
    .B1(_0681_),
    .C1(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__a31o_1 _1228_ (.A1(net57),
    .A2(_0487_),
    .A3(_0483_),
    .B1(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__inv_2 _1229_ (.A(config_cont),
    .Y(_0685_));
 sky130_fd_sc_hd__a31o_1 _1230_ (.A1(_0685_),
    .A2(_0487_),
    .A3(_0455_),
    .B1(_0672_),
    .X(_0686_));
 sky130_fd_sc_hd__o32a_1 _1231_ (.A1(_0670_),
    .A2(_0684_),
    .A3(_0686_),
    .B1(_0674_),
    .B2(\xfer.din_data[1] ),
    .X(_0081_));
 sky130_fd_sc_hd__a22o_1 _1232_ (.A1(net58),
    .A2(_0487_),
    .B1(_0503_),
    .B2(net10),
    .X(_0687_));
 sky130_fd_sc_hd__a32o_1 _1233_ (.A1(config_qspi),
    .A2(_0522_),
    .A3(_0499_),
    .B1(_0528_),
    .B2(net2),
    .X(_0688_));
 sky130_fd_sc_hd__or2_1 _1234_ (.A(_0687_),
    .B(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__a211o_1 _1235_ (.A1(net17),
    .A2(_0675_),
    .B1(_0689_),
    .C1(_0679_),
    .X(_0690_));
 sky130_fd_sc_hd__o22a_1 _1236_ (.A1(\xfer.din_data[2] ),
    .A2(_0674_),
    .B1(_0690_),
    .B2(_0673_),
    .X(_0082_));
 sky130_fd_sc_hd__a221o_1 _1237_ (.A1(net3),
    .A2(_0528_),
    .B1(_0486_),
    .B2(_0499_),
    .C1(\state[4] ),
    .X(_0691_));
 sky130_fd_sc_hd__a221o_1 _1238_ (.A1(net11),
    .A2(_0503_),
    .B1(_0675_),
    .B2(net18),
    .C1(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__a31o_1 _1239_ (.A1(net59),
    .A2(_0487_),
    .A3(_0483_),
    .B1(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__o32a_1 _1240_ (.A1(_0670_),
    .A2(_0686_),
    .A3(_0693_),
    .B1(_0674_),
    .B2(\xfer.din_data[3] ),
    .X(_0083_));
 sky130_fd_sc_hd__and3b_1 _1241_ (.A_N(config_qspi),
    .B(_0522_),
    .C(_0499_),
    .X(_0694_));
 sky130_fd_sc_hd__a221o_1 _1242_ (.A1(net13),
    .A2(_0503_),
    .B1(_0528_),
    .B2(net4),
    .C1(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__a211o_1 _1243_ (.A1(net19),
    .A2(_0675_),
    .B1(_0686_),
    .C1(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _1244_ (.A0(\xfer.din_data[4] ),
    .A1(_0696_),
    .S(_0674_),
    .X(_0697_));
 sky130_fd_sc_hd__clkbuf_1 _1245_ (.A(_0697_),
    .X(_0084_));
 sky130_fd_sc_hd__a2111o_1 _1246_ (.A1(_0499_),
    .A2(_0486_),
    .B1(_0673_),
    .C1(\state[4] ),
    .D1(_0679_),
    .X(_0698_));
 sky130_fd_sc_hd__a22o_1 _1247_ (.A1(net14),
    .A2(_0503_),
    .B1(_0528_),
    .B2(net5),
    .X(_0699_));
 sky130_fd_sc_hd__a31o_1 _1248_ (.A1(net20),
    .A2(\state[12] ),
    .A3(_0456_),
    .B1(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__o22a_1 _1249_ (.A1(\xfer.din_data[5] ),
    .A2(_0674_),
    .B1(_0698_),
    .B2(_0700_),
    .X(_0085_));
 sky130_fd_sc_hd__a22o_1 _1250_ (.A1(config_qspi),
    .A2(_0499_),
    .B1(_0503_),
    .B2(net15),
    .X(_0701_));
 sky130_fd_sc_hd__a221o_1 _1251_ (.A1(net6),
    .A2(_0528_),
    .B1(_0675_),
    .B2(net21),
    .C1(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__or2_1 _1252_ (.A(_0686_),
    .B(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _1253_ (.A0(\xfer.din_data[6] ),
    .A1(_0703_),
    .S(_0674_),
    .X(_0704_));
 sky130_fd_sc_hd__clkbuf_1 _1254_ (.A(_0704_),
    .X(_0086_));
 sky130_fd_sc_hd__a22o_1 _1255_ (.A1(net16),
    .A2(_0503_),
    .B1(_0528_),
    .B2(net7),
    .X(_0705_));
 sky130_fd_sc_hd__a31o_1 _1256_ (.A1(net22),
    .A2(\state[12] ),
    .A3(_0456_),
    .B1(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__o22a_1 _1257_ (.A1(\xfer.din_data[7] ),
    .A2(_0674_),
    .B1(_0698_),
    .B2(_0706_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _1258_ (.A0(\xfer.din_qspi ),
    .A1(config_qspi),
    .S(_0530_),
    .X(_0707_));
 sky130_fd_sc_hd__and3_1 _1259_ (.A(_0500_),
    .B(_0497_),
    .C(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__clkbuf_1 _1260_ (.A(_0708_),
    .X(_0088_));
 sky130_fd_sc_hd__a31o_1 _1261_ (.A1(_0438_),
    .A2(_0487_),
    .A3(_0454_),
    .B1(\xfer.din_rd ),
    .X(_0709_));
 sky130_fd_sc_hd__and2_1 _1262_ (.A(_0437_),
    .B(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__clkbuf_1 _1263_ (.A(_0710_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _1264_ (.A0(din_ddr),
    .A1(_0522_),
    .S(_0530_),
    .X(_0711_));
 sky130_fd_sc_hd__and3_1 _1265_ (.A(_0500_),
    .B(_0497_),
    .C(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__clkbuf_1 _1266_ (.A(_0712_),
    .X(_0090_));
 sky130_fd_sc_hd__nor2_1 _1267_ (.A(\xfer.dout_tag[1] ),
    .B(\xfer.dout_tag[2] ),
    .Y(_0713_));
 sky130_fd_sc_hd__and4_1 _1268_ (.A(\xfer.dout_tag[0] ),
    .B(_0479_),
    .C(_0491_),
    .D(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__clkbuf_4 _1269_ (.A(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _1270_ (.A0(\buffer[0] ),
    .A1(\xfer.dout_data[0] ),
    .S(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__clkbuf_1 _1271_ (.A(_0716_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _1272_ (.A0(\buffer[1] ),
    .A1(\xfer.dout_data[1] ),
    .S(_0715_),
    .X(_0717_));
 sky130_fd_sc_hd__clkbuf_1 _1273_ (.A(_0717_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _1274_ (.A0(\buffer[2] ),
    .A1(\xfer.dout_data[2] ),
    .S(_0715_),
    .X(_0718_));
 sky130_fd_sc_hd__clkbuf_1 _1275_ (.A(_0718_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _1276_ (.A0(\buffer[3] ),
    .A1(\xfer.dout_data[3] ),
    .S(_0715_),
    .X(_0719_));
 sky130_fd_sc_hd__clkbuf_1 _1277_ (.A(_0719_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _1278_ (.A0(\buffer[4] ),
    .A1(\xfer.dout_data[4] ),
    .S(_0715_),
    .X(_0720_));
 sky130_fd_sc_hd__clkbuf_1 _1279_ (.A(_0720_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _1280_ (.A0(\buffer[5] ),
    .A1(\xfer.dout_data[5] ),
    .S(_0715_),
    .X(_0721_));
 sky130_fd_sc_hd__clkbuf_1 _1281_ (.A(_0721_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _1282_ (.A0(\buffer[6] ),
    .A1(\xfer.dout_data[6] ),
    .S(_0715_),
    .X(_0722_));
 sky130_fd_sc_hd__clkbuf_1 _1283_ (.A(_0722_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _1284_ (.A0(\buffer[7] ),
    .A1(\xfer.dout_data[7] ),
    .S(_0715_),
    .X(_0723_));
 sky130_fd_sc_hd__clkbuf_1 _1285_ (.A(_0723_),
    .X(_0098_));
 sky130_fd_sc_hd__nand2_1 _1286_ (.A(\xfer.dout_tag[2] ),
    .B(_0557_),
    .Y(_0724_));
 sky130_fd_sc_hd__nor2_1 _1287_ (.A(\xfer.dout_tag[1] ),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__o21a_1 _1288_ (.A1(rd_valid),
    .A2(_0725_),
    .B1(_0437_),
    .X(_0099_));
 sky130_fd_sc_hd__buf_4 _1289_ (.A(rd_inc),
    .X(_0726_));
 sky130_fd_sc_hd__o211a_1 _1290_ (.A1(_0434_),
    .A2(_0363_),
    .B1(_0636_),
    .C1(rd_wait),
    .X(_0727_));
 sky130_fd_sc_hd__a31o_1 _1291_ (.A1(_0726_),
    .A2(_0434_),
    .A3(_0624_),
    .B1(_0727_),
    .X(_0100_));
 sky130_fd_sc_hd__nor2_1 _1292_ (.A(_0499_),
    .B(_0436_),
    .Y(_0728_));
 sky130_fd_sc_hd__o22a_1 _1293_ (.A1(_0726_),
    .A2(_0624_),
    .B1(_0728_),
    .B2(_0363_),
    .X(_0101_));
 sky130_fd_sc_hd__inv_2 _1295__2 (.A(clknet_4_0_0_clk),
    .Y(net129));
 sky130_fd_sc_hd__inv_2 _1296__3 (.A(clknet_4_0_0_clk),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _1297__4 (.A(clknet_4_1_0_clk),
    .Y(net131));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__mux2_1 _1298_ (.A0(config_en),
    .A1(net37),
    .S(net46),
    .X(_0729_));
 sky130_fd_sc_hd__or2_1 _1299_ (.A(_0361_),
    .B(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__clkbuf_1 _1300_ (.A(_0730_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_2 _1301_ (.A(net51),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_1 _1302_ (.A0(_0522_),
    .A1(net35),
    .S(net45),
    .X(_0732_));
 sky130_fd_sc_hd__and2_1 _1303_ (.A(_0731_),
    .B(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__clkbuf_1 _1304_ (.A(_0733_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _1305_ (.A0(config_qspi),
    .A1(net34),
    .S(net45),
    .X(_0734_));
 sky130_fd_sc_hd__and2_1 _1306_ (.A(_0731_),
    .B(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__clkbuf_1 _1307_ (.A(_0735_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _1308_ (.A0(config_cont),
    .A1(net33),
    .S(net45),
    .X(_0736_));
 sky130_fd_sc_hd__and2_1 _1309_ (.A(_0731_),
    .B(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__clkbuf_1 _1310_ (.A(_0737_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1311_ (.A0(net56),
    .A1(net28),
    .S(net45),
    .X(_0738_));
 sky130_fd_sc_hd__and2_1 _1312_ (.A(_0731_),
    .B(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__clkbuf_1 _1313_ (.A(_0739_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _1314_ (.A0(net57),
    .A1(net29),
    .S(net45),
    .X(_0740_));
 sky130_fd_sc_hd__and2_1 _1315_ (.A(_0731_),
    .B(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__clkbuf_1 _1316_ (.A(_0741_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _1317_ (.A0(net58),
    .A1(net30),
    .S(net45),
    .X(_0742_));
 sky130_fd_sc_hd__and2_1 _1318_ (.A(_0731_),
    .B(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__clkbuf_1 _1319_ (.A(_0743_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _1320_ (.A0(net59),
    .A1(net31),
    .S(net45),
    .X(_0744_));
 sky130_fd_sc_hd__or2_1 _1321_ (.A(_0361_),
    .B(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__clkbuf_1 _1322_ (.A(_0745_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _1323_ (.A0(\config_oe[0] ),
    .A1(net41),
    .S(net44),
    .X(_0746_));
 sky130_fd_sc_hd__and2_1 _1324_ (.A(_0731_),
    .B(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__clkbuf_1 _1325_ (.A(_0747_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _1326_ (.A0(\config_oe[1] ),
    .A1(net42),
    .S(net44),
    .X(_0748_));
 sky130_fd_sc_hd__and2_1 _1327_ (.A(_0731_),
    .B(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__clkbuf_1 _1328_ (.A(_0749_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _1329_ (.A0(\config_oe[2] ),
    .A1(net26),
    .S(net44),
    .X(_0750_));
 sky130_fd_sc_hd__and2_1 _1330_ (.A(_0731_),
    .B(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__clkbuf_1 _1331_ (.A(_0751_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _1332_ (.A0(\config_oe[3] ),
    .A1(net27),
    .S(net44),
    .X(_0752_));
 sky130_fd_sc_hd__and2_1 _1333_ (.A(_0731_),
    .B(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__clkbuf_1 _1334_ (.A(_0753_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _1335_ (.A0(config_csb),
    .A1(net40),
    .S(net43),
    .X(_0754_));
 sky130_fd_sc_hd__and2_1 _1336_ (.A(net51),
    .B(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__clkbuf_1 _1337_ (.A(_0755_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _1338_ (.A0(config_clk),
    .A1(net39),
    .S(net43),
    .X(_0756_));
 sky130_fd_sc_hd__and2_1 _1339_ (.A(net51),
    .B(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__clkbuf_1 _1340_ (.A(_0757_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _1341_ (.A0(\config_do[0] ),
    .A1(net25),
    .S(net43),
    .X(_0758_));
 sky130_fd_sc_hd__and2_1 _1342_ (.A(net51),
    .B(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__clkbuf_1 _1343_ (.A(_0759_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _1344_ (.A0(\config_do[1] ),
    .A1(net32),
    .S(net43),
    .X(_0760_));
 sky130_fd_sc_hd__and2_1 _1345_ (.A(net51),
    .B(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__clkbuf_1 _1346_ (.A(_0761_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _1347_ (.A0(\config_do[2] ),
    .A1(net36),
    .S(net43),
    .X(_0762_));
 sky130_fd_sc_hd__and2_1 _1348_ (.A(net51),
    .B(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__clkbuf_1 _1349_ (.A(_0763_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _1350_ (.A0(\config_do[3] ),
    .A1(net38),
    .S(net43),
    .X(_0764_));
 sky130_fd_sc_hd__and2_1 _1351_ (.A(net51),
    .B(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__clkbuf_1 _1352_ (.A(_0765_),
    .X(_0119_));
 sky130_fd_sc_hd__or3_1 _1353_ (.A(net43),
    .B(net44),
    .C(net45),
    .X(_0170_));
 sky130_fd_sc_hd__or4_1 _1354_ (.A(_0537_),
    .B(net46),
    .C(_0361_),
    .D(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__clkbuf_1 _1355_ (.A(_0171_),
    .X(_0120_));
 sky130_fd_sc_hd__nand2_1 _1356_ (.A(_0438_),
    .B(_0453_),
    .Y(_0121_));
 sky130_fd_sc_hd__mux2_1 _1357_ (.A0(net47),
    .A1(net48),
    .S(_0536_),
    .X(_0172_));
 sky130_fd_sc_hd__a21o_1 _1358_ (.A1(\xfer.xfer_ddr ),
    .A2(_0464_),
    .B1(_0448_),
    .X(_0173_));
 sky130_fd_sc_hd__nand3_4 _1359_ (.A(_0438_),
    .B(_0569_),
    .C(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__mux2_1 _1360_ (.A0(_0172_),
    .A1(\xfer.dout_data[0] ),
    .S(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__clkbuf_1 _1361_ (.A(_0175_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _1362_ (.A0(net48),
    .A1(\xfer.dout_data[0] ),
    .S(_0536_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _1363_ (.A0(_0176_),
    .A1(\xfer.dout_data[1] ),
    .S(_0174_),
    .X(_0177_));
 sky130_fd_sc_hd__clkbuf_1 _1364_ (.A(_0177_),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_1 _1365_ (.A1(_0542_),
    .A2(net49),
    .B1(\xfer.dout_data[1] ),
    .B2(_0536_),
    .X(_0178_));
 sky130_fd_sc_hd__a21o_1 _1366_ (.A1(\xfer.dout_data[0] ),
    .A2(_0592_),
    .B1(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _1367_ (.A0(_0179_),
    .A1(\xfer.dout_data[2] ),
    .S(_0174_),
    .X(_0180_));
 sky130_fd_sc_hd__clkbuf_1 _1368_ (.A(_0180_),
    .X(_0124_));
 sky130_fd_sc_hd__a22o_1 _1369_ (.A1(_0542_),
    .A2(net50),
    .B1(\xfer.dout_data[2] ),
    .B2(_0536_),
    .X(_0181_));
 sky130_fd_sc_hd__a21o_1 _1370_ (.A1(\xfer.dout_data[1] ),
    .A2(_0592_),
    .B1(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _1371_ (.A0(_0182_),
    .A1(\xfer.dout_data[3] ),
    .S(_0174_),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_1 _1372_ (.A(_0183_),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _1373_ (.A1(_0542_),
    .A2(\xfer.dout_data[0] ),
    .B1(\xfer.dout_data[3] ),
    .B2(_0536_),
    .X(_0184_));
 sky130_fd_sc_hd__a21o_1 _1374_ (.A1(\xfer.dout_data[2] ),
    .A2(_0592_),
    .B1(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _1375_ (.A0(_0185_),
    .A1(\xfer.dout_data[4] ),
    .S(_0174_),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_1 _1376_ (.A(_0186_),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_1 _1377_ (.A1(_0542_),
    .A2(\xfer.dout_data[1] ),
    .B1(\xfer.dout_data[4] ),
    .B2(_0536_),
    .X(_0187_));
 sky130_fd_sc_hd__a21o_1 _1378_ (.A1(\xfer.dout_data[3] ),
    .A2(_0592_),
    .B1(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _1379_ (.A0(_0188_),
    .A1(\xfer.dout_data[5] ),
    .S(_0174_),
    .X(_0189_));
 sky130_fd_sc_hd__clkbuf_1 _1380_ (.A(_0189_),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_1 _1381_ (.A1(_0542_),
    .A2(\xfer.dout_data[2] ),
    .B1(\xfer.dout_data[5] ),
    .B2(_0535_),
    .X(_0190_));
 sky130_fd_sc_hd__a21o_1 _1382_ (.A1(\xfer.dout_data[4] ),
    .A2(_0592_),
    .B1(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _1383_ (.A0(_0191_),
    .A1(\xfer.dout_data[6] ),
    .S(_0174_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _1384_ (.A(_0192_),
    .X(_0128_));
 sky130_fd_sc_hd__a22o_1 _1385_ (.A1(_0542_),
    .A2(\xfer.dout_data[3] ),
    .B1(\xfer.dout_data[6] ),
    .B2(_0535_),
    .X(_0193_));
 sky130_fd_sc_hd__a21o_1 _1386_ (.A1(\xfer.dout_data[5] ),
    .A2(_0592_),
    .B1(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _1387_ (.A0(_0194_),
    .A1(\xfer.dout_data[7] ),
    .S(_0174_),
    .X(_0195_));
 sky130_fd_sc_hd__clkbuf_1 _1388_ (.A(_0195_),
    .X(_0129_));
 sky130_fd_sc_hd__a22o_1 _1389_ (.A1(\xfer.din_rd ),
    .A2(_0526_),
    .B1(_0669_),
    .B2(\xfer.xfer_rd ),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_1 _1390_ (.A1(\xfer.din_qspi ),
    .A2(_0526_),
    .B1(_0669_),
    .B2(_0542_),
    .X(_0131_));
 sky130_fd_sc_hd__xnor2_1 _1391_ (.A(_0459_),
    .B(\xfer.dummy_count[0] ),
    .Y(_0196_));
 sky130_fd_sc_hd__nor2_1 _1392_ (.A(_0526_),
    .B(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__and3_1 _1393_ (.A(\xfer.din_rd ),
    .B(\xfer.din_data[0] ),
    .C(_0483_),
    .X(_0198_));
 sky130_fd_sc_hd__o21a_1 _1394_ (.A1(_0197_),
    .A2(_0198_),
    .B1(_0620_),
    .X(_0132_));
 sky130_fd_sc_hd__o21ai_1 _1395_ (.A1(_0448_),
    .A2(\xfer.dummy_count[0] ),
    .B1(\xfer.dummy_count[1] ),
    .Y(_0199_));
 sky130_fd_sc_hd__or3_1 _1396_ (.A(_0448_),
    .B(\xfer.dummy_count[1] ),
    .C(\xfer.dummy_count[0] ),
    .X(_0200_));
 sky130_fd_sc_hd__a21oi_1 _1397_ (.A1(_0199_),
    .A2(_0200_),
    .B1(_0483_),
    .Y(_0201_));
 sky130_fd_sc_hd__and3_1 _1398_ (.A(\xfer.din_rd ),
    .B(\xfer.din_data[1] ),
    .C(_0483_),
    .X(_0202_));
 sky130_fd_sc_hd__o21a_1 _1399_ (.A1(_0201_),
    .A2(_0202_),
    .B1(_0620_),
    .X(_0133_));
 sky130_fd_sc_hd__nor2_1 _1400_ (.A(\xfer.dummy_count[2] ),
    .B(_0200_),
    .Y(_0203_));
 sky130_fd_sc_hd__and2_1 _1401_ (.A(\xfer.dummy_count[2] ),
    .B(_0200_),
    .X(_0204_));
 sky130_fd_sc_hd__o21a_1 _1402_ (.A1(_0203_),
    .A2(_0204_),
    .B1(_0456_),
    .X(_0205_));
 sky130_fd_sc_hd__and3_1 _1403_ (.A(\xfer.din_rd ),
    .B(\xfer.din_data[2] ),
    .C(_0483_),
    .X(_0206_));
 sky130_fd_sc_hd__o21a_1 _1404_ (.A1(_0205_),
    .A2(_0206_),
    .B1(_0620_),
    .X(_0134_));
 sky130_fd_sc_hd__xor2_1 _1405_ (.A(\xfer.dummy_count[3] ),
    .B(_0203_),
    .X(_0207_));
 sky130_fd_sc_hd__a32o_1 _1406_ (.A1(\xfer.din_rd ),
    .A2(\xfer.din_data[3] ),
    .A3(_0483_),
    .B1(_0478_),
    .B2(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__and2_1 _1407_ (.A(_0620_),
    .B(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__clkbuf_1 _1408_ (.A(_0209_),
    .X(_0135_));
 sky130_fd_sc_hd__inv_1 _1409_ (.A(\xfer.count[1] ),
    .Y(_0210_));
 sky130_fd_sc_hd__inv_2 _1410_ (.A(\xfer.count[0] ),
    .Y(_0211_));
 sky130_fd_sc_hd__a21o_1 _1411_ (.A1(_0211_),
    .A2(_0459_),
    .B1(_0466_),
    .X(_0212_));
 sky130_fd_sc_hd__o2111a_1 _1412_ (.A1(_0459_),
    .A2(_0535_),
    .B1(_0569_),
    .C1(_0212_),
    .D1(_0449_),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_1 _1413_ (.A1(_0462_),
    .A2(_0585_),
    .B1(_0610_),
    .B2(_0535_),
    .X(_0214_));
 sky130_fd_sc_hd__a2bb2o_1 _1414_ (.A1_N(_0210_),
    .A2_N(_0213_),
    .B1(_0569_),
    .B2(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__and3_1 _1415_ (.A(_0438_),
    .B(_0478_),
    .C(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__clkbuf_1 _1416_ (.A(_0216_),
    .X(_0136_));
 sky130_fd_sc_hd__nand2_1 _1417_ (.A(_0459_),
    .B(_0470_),
    .Y(_0217_));
 sky130_fd_sc_hd__a21o_1 _1418_ (.A1(_0451_),
    .A2(_0217_),
    .B1(_0611_),
    .X(_0218_));
 sky130_fd_sc_hd__nor2_1 _1419_ (.A(_0451_),
    .B(_0450_),
    .Y(_0219_));
 sky130_fd_sc_hd__a221o_1 _1420_ (.A1(_0534_),
    .A2(_0218_),
    .B1(_0219_),
    .B2(_0460_),
    .C1(_0585_),
    .X(_0220_));
 sky130_fd_sc_hd__a31o_1 _1421_ (.A1(_0465_),
    .A2(_0541_),
    .A3(_0475_),
    .B1(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__o31ai_1 _1422_ (.A1(_0542_),
    .A2(_0536_),
    .A3(_0462_),
    .B1(_0569_),
    .Y(_0222_));
 sky130_fd_sc_hd__a32o_1 _1423_ (.A1(_0569_),
    .A2(_0613_),
    .A3(_0221_),
    .B1(_0222_),
    .B2(_0451_),
    .X(_0223_));
 sky130_fd_sc_hd__and3_1 _1424_ (.A(_0438_),
    .B(_0478_),
    .C(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__clkbuf_1 _1425_ (.A(_0224_),
    .X(_0137_));
 sky130_fd_sc_hd__inv_2 _1426_ (.A(_0667_),
    .Y(_0225_));
 sky130_fd_sc_hd__a211o_1 _1427_ (.A1(\state[3] ),
    .A2(_0492_),
    .B1(_0520_),
    .C1(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__or2b_1 _1428_ (.A(\xfer.din_tag[0] ),
    .B_N(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__o311a_1 _1429_ (.A1(\state[8] ),
    .A2(\state[11] ),
    .A3(_0226_),
    .B1(_0227_),
    .C1(_0500_),
    .X(_0138_));
 sky130_fd_sc_hd__or2b_1 _1430_ (.A(\xfer.din_tag[1] ),
    .B_N(_0226_),
    .X(_0228_));
 sky130_fd_sc_hd__o311a_1 _1431_ (.A1(\state[5] ),
    .A2(\state[11] ),
    .A3(_0226_),
    .B1(_0228_),
    .C1(_0500_),
    .X(_0139_));
 sky130_fd_sc_hd__a32o_1 _1432_ (.A1(\xfer.din_tag[2] ),
    .A2(_0500_),
    .A3(_0226_),
    .B1(_0671_),
    .B2(_0524_),
    .X(_0140_));
 sky130_fd_sc_hd__a32o_1 _1433_ (.A1(\xfer.din_qspi ),
    .A2(din_ddr),
    .A3(_0526_),
    .B1(_0669_),
    .B2(\xfer.xfer_ddr ),
    .X(_0141_));
 sky130_fd_sc_hd__inv_2 _1434_ (.A(\xfer.din_qspi ),
    .Y(_0229_));
 sky130_fd_sc_hd__a32o_1 _1435_ (.A1(_0229_),
    .A2(din_ddr),
    .A3(_0526_),
    .B1(_0669_),
    .B2(\xfer.xfer_dspi ),
    .X(_0142_));
 sky130_fd_sc_hd__o21ai_1 _1436_ (.A1(\xfer.flash_csb ),
    .A2(_0609_),
    .B1(_0448_),
    .Y(_0230_));
 sky130_fd_sc_hd__o211a_1 _1437_ (.A1(_0448_),
    .A2(_0609_),
    .B1(_0669_),
    .C1(_0230_),
    .X(_0143_));
 sky130_fd_sc_hd__a21o_1 _1438_ (.A1(\xfer.flash_csb ),
    .A2(_0478_),
    .B1(_0457_),
    .X(_0144_));
 sky130_fd_sc_hd__inv_2 _1439_ (.A(rd_inc),
    .Y(_0231_));
 sky130_fd_sc_hd__buf_4 _1440_ (.A(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__and4bb_4 _1441_ (.A_N(_0724_),
    .B_N(\xfer.dout_tag[1] ),
    .C(_0232_),
    .D(_0479_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _1442_ (.A0(\rd_addr[0] ),
    .A1(net1),
    .S(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__clkbuf_1 _1443_ (.A(_0234_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(\rd_addr[1] ),
    .A1(net12),
    .S(_0233_),
    .X(_0235_));
 sky130_fd_sc_hd__clkbuf_1 _1445_ (.A(_0235_),
    .X(_0146_));
 sky130_fd_sc_hd__inv_1 _1446_ (.A(\rd_addr[2] ),
    .Y(_0236_));
 sky130_fd_sc_hd__buf_4 _1447_ (.A(rd_inc),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _1448_ (.A0(net17),
    .A1(_0236_),
    .S(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _1449_ (.A0(\rd_addr[2] ),
    .A1(_0238_),
    .S(_0629_),
    .X(_0239_));
 sky130_fd_sc_hd__clkbuf_1 _1450_ (.A(_0239_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _1451_ (.A0(net18),
    .A1(_0412_),
    .S(_0237_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _1452_ (.A0(\rd_addr[3] ),
    .A1(_0240_),
    .S(_0629_),
    .X(_0241_));
 sky130_fd_sc_hd__clkbuf_1 _1453_ (.A(_0241_),
    .X(_0148_));
 sky130_fd_sc_hd__nor2_1 _1454_ (.A(_0404_),
    .B(_0405_),
    .Y(_0242_));
 sky130_fd_sc_hd__mux2_1 _1455_ (.A0(net19),
    .A1(_0242_),
    .S(_0237_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _1456_ (.A0(\rd_addr[4] ),
    .A1(_0243_),
    .S(_0629_),
    .X(_0244_));
 sky130_fd_sc_hd__clkbuf_1 _1457_ (.A(_0244_),
    .X(_0149_));
 sky130_fd_sc_hd__nor2_1 _1458_ (.A(\rd_addr[5] ),
    .B(_0404_),
    .Y(_0245_));
 sky130_fd_sc_hd__o21ai_1 _1459_ (.A1(_0376_),
    .A2(_0245_),
    .B1(_0237_),
    .Y(_0246_));
 sky130_fd_sc_hd__o21a_1 _1460_ (.A1(_0726_),
    .A2(net20),
    .B1(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _1461_ (.A0(\rd_addr[5] ),
    .A1(_0247_),
    .S(_0629_),
    .X(_0248_));
 sky130_fd_sc_hd__clkbuf_1 _1462_ (.A(_0248_),
    .X(_0150_));
 sky130_fd_sc_hd__or3_4 _1463_ (.A(\xfer.dout_tag[1] ),
    .B(_0363_),
    .C(_0724_),
    .X(_0249_));
 sky130_fd_sc_hd__xnor2_1 _1464_ (.A(\rd_addr[6] ),
    .B(_0376_),
    .Y(_0250_));
 sky130_fd_sc_hd__nor2_1 _1465_ (.A(_0726_),
    .B(net21),
    .Y(_0251_));
 sky130_fd_sc_hd__a211o_1 _1466_ (.A1(_0726_),
    .A2(_0250_),
    .B1(_0251_),
    .C1(_0249_),
    .X(_0252_));
 sky130_fd_sc_hd__a21bo_1 _1467_ (.A1(\rd_addr[6] ),
    .A2(_0249_),
    .B1_N(_0252_),
    .X(_0151_));
 sky130_fd_sc_hd__nand2_1 _1468_ (.A(_0376_),
    .B(_0367_),
    .Y(_0253_));
 sky130_fd_sc_hd__a21o_1 _1469_ (.A1(\rd_addr[6] ),
    .A2(_0376_),
    .B1(\rd_addr[7] ),
    .X(_0254_));
 sky130_fd_sc_hd__and2_1 _1470_ (.A(_0232_),
    .B(net22),
    .X(_0255_));
 sky130_fd_sc_hd__a31o_1 _1471_ (.A1(_0726_),
    .A2(_0253_),
    .A3(_0254_),
    .B1(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _1472_ (.A0(\rd_addr[7] ),
    .A1(_0256_),
    .S(_0629_),
    .X(_0257_));
 sky130_fd_sc_hd__clkbuf_1 _1473_ (.A(_0257_),
    .X(_0152_));
 sky130_fd_sc_hd__or3_1 _1474_ (.A(_0231_),
    .B(_0399_),
    .C(_0400_),
    .X(_0258_));
 sky130_fd_sc_hd__a21bo_1 _1475_ (.A1(_0232_),
    .A2(net23),
    .B1_N(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _1476_ (.A0(\rd_addr[8] ),
    .A1(_0259_),
    .S(_0629_),
    .X(_0260_));
 sky130_fd_sc_hd__clkbuf_1 _1477_ (.A(_0260_),
    .X(_0153_));
 sky130_fd_sc_hd__inv_2 _1478_ (.A(_0402_),
    .Y(_0261_));
 sky130_fd_sc_hd__o211a_1 _1479_ (.A1(\rd_addr[9] ),
    .A2(_0399_),
    .B1(_0261_),
    .C1(_0726_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _1480_ (.A0(_0262_),
    .A1(\rd_addr[9] ),
    .S(_0249_),
    .X(_0263_));
 sky130_fd_sc_hd__a21o_1 _1481_ (.A1(net24),
    .A2(_0233_),
    .B1(_0263_),
    .X(_0154_));
 sky130_fd_sc_hd__nor2_1 _1482_ (.A(\rd_addr[10] ),
    .B(_0402_),
    .Y(_0264_));
 sky130_fd_sc_hd__nor2_1 _1483_ (.A(_0419_),
    .B(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__mux2_1 _1484_ (.A0(net2),
    .A1(_0265_),
    .S(_0237_),
    .X(_0266_));
 sky130_fd_sc_hd__buf_4 _1485_ (.A(_0623_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _1486_ (.A0(\rd_addr[10] ),
    .A1(_0266_),
    .S(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__clkbuf_1 _1487_ (.A(_0268_),
    .X(_0155_));
 sky130_fd_sc_hd__xor2_1 _1488_ (.A(\rd_addr[11] ),
    .B(_0419_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _1489_ (.A0(net3),
    .A1(_0269_),
    .S(_0237_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _1490_ (.A0(\rd_addr[11] ),
    .A1(_0270_),
    .S(_0267_),
    .X(_0271_));
 sky130_fd_sc_hd__clkbuf_1 _1491_ (.A(_0271_),
    .X(_0156_));
 sky130_fd_sc_hd__nor2_1 _1492_ (.A(_0232_),
    .B(_0371_),
    .Y(_0272_));
 sky130_fd_sc_hd__a21o_1 _1493_ (.A1(\rd_addr[11] ),
    .A2(_0419_),
    .B1(\rd_addr[12] ),
    .X(_0273_));
 sky130_fd_sc_hd__a22o_1 _1494_ (.A1(_0232_),
    .A2(net4),
    .B1(_0272_),
    .B2(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _1495_ (.A0(\rd_addr[12] ),
    .A1(_0274_),
    .S(_0267_),
    .X(_0275_));
 sky130_fd_sc_hd__clkbuf_1 _1496_ (.A(_0275_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _1497_ (.A0(_0334_),
    .A1(_0388_),
    .S(_0726_),
    .X(_0276_));
 sky130_fd_sc_hd__nand2_1 _1498_ (.A(_0624_),
    .B(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__o21a_1 _1499_ (.A1(_0333_),
    .A2(_0624_),
    .B1(_0277_),
    .X(_0158_));
 sky130_fd_sc_hd__nor2_1 _1500_ (.A(\rd_addr[14] ),
    .B(_0378_),
    .Y(_0278_));
 sky130_fd_sc_hd__nor2_1 _1501_ (.A(_0392_),
    .B(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__mux2_1 _1502_ (.A0(net6),
    .A1(_0279_),
    .S(_0237_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _1503_ (.A0(\rd_addr[14] ),
    .A1(_0280_),
    .S(_0267_),
    .X(_0281_));
 sky130_fd_sc_hd__clkbuf_1 _1504_ (.A(_0281_),
    .X(_0159_));
 sky130_fd_sc_hd__inv_2 _1505_ (.A(_0395_),
    .Y(_0282_));
 sky130_fd_sc_hd__o211a_1 _1506_ (.A1(\rd_addr[15] ),
    .A2(_0392_),
    .B1(_0282_),
    .C1(_0237_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _1507_ (.A0(_0283_),
    .A1(\rd_addr[15] ),
    .S(_0249_),
    .X(_0284_));
 sky130_fd_sc_hd__a21o_1 _1508_ (.A1(net7),
    .A2(_0233_),
    .B1(_0284_),
    .X(_0160_));
 sky130_fd_sc_hd__nor2_1 _1509_ (.A(\rd_addr[16] ),
    .B(_0395_),
    .Y(_0285_));
 sky130_fd_sc_hd__o21ai_1 _1510_ (.A1(_0285_),
    .A2(_0383_),
    .B1(_0237_),
    .Y(_0286_));
 sky130_fd_sc_hd__o21a_1 _1511_ (.A1(_0726_),
    .A2(net8),
    .B1(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _1512_ (.A0(\rd_addr[16] ),
    .A1(_0287_),
    .S(_0267_),
    .X(_0288_));
 sky130_fd_sc_hd__clkbuf_1 _1513_ (.A(_0288_),
    .X(_0161_));
 sky130_fd_sc_hd__o21ba_1 _1514_ (.A1(\rd_addr[17] ),
    .A2(_0383_),
    .B1_N(_0373_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _1515_ (.A0(net9),
    .A1(_0289_),
    .S(_0237_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _1516_ (.A0(\rd_addr[17] ),
    .A1(_0290_),
    .S(_0267_),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _1517_ (.A(_0291_),
    .X(_0162_));
 sky130_fd_sc_hd__xor2_1 _1518_ (.A(\rd_addr[18] ),
    .B(_0373_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _1519_ (.A0(net10),
    .A1(_0292_),
    .S(rd_inc),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _1520_ (.A0(\rd_addr[18] ),
    .A1(_0293_),
    .S(_0267_),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_1 _1521_ (.A(_0294_),
    .X(_0163_));
 sky130_fd_sc_hd__a31o_1 _1522_ (.A1(_0500_),
    .A2(_0387_),
    .A3(_0725_),
    .B1(\rd_addr[19] ),
    .X(_0295_));
 sky130_fd_sc_hd__a31o_1 _1523_ (.A1(\rd_addr[18] ),
    .A2(\rd_addr[19] ),
    .A3(_0373_),
    .B1(_0232_),
    .X(_0296_));
 sky130_fd_sc_hd__nand2_1 _1524_ (.A(_0624_),
    .B(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__a22o_1 _1525_ (.A1(net11),
    .A2(_0233_),
    .B1(_0295_),
    .B2(_0297_),
    .X(_0164_));
 sky130_fd_sc_hd__and3_1 _1526_ (.A(rd_inc),
    .B(_0374_),
    .C(_0379_),
    .X(_0298_));
 sky130_fd_sc_hd__a21o_1 _1527_ (.A1(_0232_),
    .A2(net13),
    .B1(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _1528_ (.A0(\rd_addr[20] ),
    .A1(_0299_),
    .S(_0267_),
    .X(_0300_));
 sky130_fd_sc_hd__clkbuf_1 _1529_ (.A(_0300_),
    .X(_0165_));
 sky130_fd_sc_hd__nor2_1 _1530_ (.A(_0232_),
    .B(_0428_),
    .Y(_0301_));
 sky130_fd_sc_hd__a21o_1 _1531_ (.A1(_0232_),
    .A2(net14),
    .B1(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _1532_ (.A0(\rd_addr[21] ),
    .A1(_0302_),
    .S(_0267_),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_1 _1533_ (.A(_0303_),
    .X(_0166_));
 sky130_fd_sc_hd__nor2_1 _1534_ (.A(\rd_addr[22] ),
    .B(_0430_),
    .Y(_0304_));
 sky130_fd_sc_hd__nor2_1 _1535_ (.A(_0382_),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__mux2_1 _1536_ (.A0(net15),
    .A1(_0305_),
    .S(rd_inc),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _1537_ (.A0(\rd_addr[22] ),
    .A1(_0306_),
    .S(_0267_),
    .X(_0307_));
 sky130_fd_sc_hd__clkbuf_1 _1538_ (.A(_0307_),
    .X(_0167_));
 sky130_fd_sc_hd__and2_1 _1539_ (.A(_0232_),
    .B(net16),
    .X(_0308_));
 sky130_fd_sc_hd__or2_1 _1540_ (.A(\rd_addr[23] ),
    .B(_0382_),
    .X(_0309_));
 sky130_fd_sc_hd__a31o_1 _1541_ (.A1(_0726_),
    .A2(_0432_),
    .A3(_0309_),
    .B1(_0636_),
    .X(_0310_));
 sky130_fd_sc_hd__o22a_1 _1542_ (.A1(\rd_addr[23] ),
    .A2(_0624_),
    .B1(_0308_),
    .B2(_0310_),
    .X(_0168_));
 sky130_fd_sc_hd__or4_1 _1543_ (.A(_0211_),
    .B(_0446_),
    .C(_0466_),
    .D(_0461_),
    .X(_0311_));
 sky130_fd_sc_hd__a41o_1 _1544_ (.A1(_0459_),
    .A2(_0533_),
    .A3(_0536_),
    .A4(_0460_),
    .B1(\xfer.count[0] ),
    .X(_0312_));
 sky130_fd_sc_hd__and3_1 _1545_ (.A(_0669_),
    .B(_0311_),
    .C(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_1 _1546_ (.A(_0313_),
    .X(_0169_));
 sky130_fd_sc_hd__dfxtp_1 _1547_ (.CLK(clknet_4_11_0_clk),
    .D(_0017_),
    .Q(\buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1548_ (.CLK(clknet_4_11_0_clk),
    .D(_0018_),
    .Q(\buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1549_ (.CLK(clknet_4_11_0_clk),
    .D(_0019_),
    .Q(\buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1550_ (.CLK(clknet_4_14_0_clk),
    .D(_0020_),
    .Q(\buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1551_ (.CLK(clknet_4_14_0_clk),
    .D(_0021_),
    .Q(\buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1552_ (.CLK(clknet_4_11_0_clk),
    .D(_0022_),
    .Q(\buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1553_ (.CLK(clknet_4_14_0_clk),
    .D(_0023_),
    .Q(\buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1554_ (.CLK(clknet_4_11_0_clk),
    .D(_0024_),
    .Q(\buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1555_ (.CLK(clknet_4_3_0_clk),
    .D(_0025_),
    .Q(\xfer.obuffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1556_ (.CLK(clknet_4_15_0_clk),
    .D(_0026_),
    .Q(\buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1557_ (.CLK(clknet_4_15_0_clk),
    .D(_0027_),
    .Q(\buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1558_ (.CLK(clknet_4_15_0_clk),
    .D(_0028_),
    .Q(\buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1559_ (.CLK(clknet_4_14_0_clk),
    .D(_0029_),
    .Q(\buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1560_ (.CLK(clknet_4_15_0_clk),
    .D(_0030_),
    .Q(\buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1561_ (.CLK(clknet_4_15_0_clk),
    .D(_0031_),
    .Q(\buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1562_ (.CLK(clknet_4_15_0_clk),
    .D(_0032_),
    .Q(\buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1563_ (.CLK(clknet_4_14_0_clk),
    .D(_0033_),
    .Q(\buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1564_ (.CLK(clknet_4_2_0_clk),
    .D(_0034_),
    .Q(\xfer.obuffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1565_ (.CLK(clknet_4_0_0_clk),
    .D(_0035_),
    .Q(\xfer.obuffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1566_ (.CLK(clknet_4_0_0_clk),
    .D(_0036_),
    .Q(\xfer.obuffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1567_ (.CLK(clknet_4_0_0_clk),
    .D(_0037_),
    .Q(\xfer.obuffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1568_ (.CLK(clknet_4_1_0_clk),
    .D(_0038_),
    .Q(\xfer.obuffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1569_ (.CLK(clknet_4_0_0_clk),
    .D(_0039_),
    .Q(\xfer.obuffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1570_ (.CLK(clknet_4_1_0_clk),
    .D(_0040_),
    .Q(\xfer.obuffer[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1571_ (.CLK(clknet_4_4_0_clk),
    .D(_0041_),
    .Q(\xfer.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1572_ (.CLK(clknet_4_4_0_clk),
    .D(_0042_),
    .Q(\xfer.last_fetch ));
 sky130_fd_sc_hd__dfxtp_1 _1573_ (.CLK(clknet_4_13_0_clk),
    .D(_0043_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _1574_ (.CLK(clknet_4_13_0_clk),
    .D(_0044_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_1 _1575_ (.CLK(clknet_4_13_0_clk),
    .D(_0045_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_1 _1576_ (.CLK(clknet_4_12_0_clk),
    .D(_0046_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_1 _1577_ (.CLK(clknet_4_13_0_clk),
    .D(_0047_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_1 _1578_ (.CLK(clknet_4_13_0_clk),
    .D(_0048_),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_1 _1579_ (.CLK(clknet_4_13_0_clk),
    .D(_0049_),
    .Q(net109));
 sky130_fd_sc_hd__dfxtp_1 _1580_ (.CLK(clknet_4_11_0_clk),
    .D(_0050_),
    .Q(net110));
 sky130_fd_sc_hd__dfxtp_1 _1581_ (.CLK(clknet_4_11_0_clk),
    .D(_0051_),
    .Q(net111));
 sky130_fd_sc_hd__dfxtp_1 _1582_ (.CLK(clknet_4_12_0_clk),
    .D(_0052_),
    .Q(net112));
 sky130_fd_sc_hd__dfxtp_1 _1583_ (.CLK(clknet_4_11_0_clk),
    .D(_0053_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _1584_ (.CLK(clknet_4_14_0_clk),
    .D(_0054_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_1 _1585_ (.CLK(clknet_4_14_0_clk),
    .D(_0055_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_1 _1586_ (.CLK(clknet_4_11_0_clk),
    .D(_0056_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_1 _1587_ (.CLK(clknet_4_14_0_clk),
    .D(_0057_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_1 _1588_ (.CLK(clknet_4_14_0_clk),
    .D(_0058_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_1 _1589_ (.CLK(clknet_4_15_0_clk),
    .D(_0059_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _1590_ (.CLK(clknet_4_15_0_clk),
    .D(_0060_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_1 _1591_ (.CLK(clknet_4_15_0_clk),
    .D(_0061_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_1 _1592_ (.CLK(clknet_4_14_0_clk),
    .D(_0062_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_1 _1593_ (.CLK(clknet_4_15_0_clk),
    .D(_0063_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_1 _1594_ (.CLK(clknet_4_15_0_clk),
    .D(_0064_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_1 _1595_ (.CLK(clknet_4_15_0_clk),
    .D(_0065_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_1 _1596_ (.CLK(clknet_4_14_0_clk),
    .D(_0066_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _1597_ (.CLK(clknet_4_15_0_clk),
    .D(_0067_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_1 _1598_ (.CLK(clknet_4_15_0_clk),
    .D(_0068_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _1599_ (.CLK(clknet_4_15_0_clk),
    .D(_0069_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _1600_ (.CLK(clknet_4_14_0_clk),
    .D(_0070_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_1 _1601_ (.CLK(clknet_4_15_0_clk),
    .D(_0071_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _1602_ (.CLK(clknet_4_15_0_clk),
    .D(_0072_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_1 _1603_ (.CLK(clknet_4_15_0_clk),
    .D(_0073_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_1 _1604_ (.CLK(clknet_4_14_0_clk),
    .D(_0074_),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_1 _1605_ (.CLK(clknet_4_5_0_clk),
    .D(_0075_),
    .Q(\xfer.resetn ));
 sky130_fd_sc_hd__dfxtp_1 _1606_ (.CLK(clknet_4_4_0_clk),
    .D(_0076_),
    .Q(\xfer.din_valid ));
 sky130_fd_sc_hd__dfxtp_1 _1607_ (.CLK(clknet_4_12_0_clk),
    .D(_0077_),
    .Q(\xfer.xfer_tag[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1608_ (.CLK(clknet_4_3_0_clk),
    .D(_0078_),
    .Q(\xfer.xfer_tag[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1609_ (.CLK(clknet_4_6_0_clk),
    .D(_0079_),
    .Q(\xfer.xfer_tag[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1610_ (.CLK(clknet_4_3_0_clk),
    .D(_0080_),
    .Q(\xfer.din_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1611_ (.CLK(clknet_4_3_0_clk),
    .D(_0081_),
    .Q(\xfer.din_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1612_ (.CLK(clknet_4_3_0_clk),
    .D(_0082_),
    .Q(\xfer.din_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1613_ (.CLK(clknet_4_3_0_clk),
    .D(_0083_),
    .Q(\xfer.din_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1614_ (.CLK(clknet_4_2_0_clk),
    .D(_0084_),
    .Q(\xfer.din_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1615_ (.CLK(clknet_4_3_0_clk),
    .D(_0085_),
    .Q(\xfer.din_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1616_ (.CLK(clknet_4_2_0_clk),
    .D(_0086_),
    .Q(\xfer.din_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1617_ (.CLK(clknet_4_3_0_clk),
    .D(_0087_),
    .Q(\xfer.din_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1618_ (.CLK(clknet_4_5_0_clk),
    .D(_0088_),
    .Q(\xfer.din_qspi ));
 sky130_fd_sc_hd__dfxtp_1 _1619_ (.CLK(clknet_4_6_0_clk),
    .D(_0089_),
    .Q(\xfer.din_rd ));
 sky130_fd_sc_hd__dfxtp_1 _1620_ (.CLK(clknet_4_4_0_clk),
    .D(_0090_),
    .Q(din_ddr));
 sky130_fd_sc_hd__dfxtp_1 _1621_ (.CLK(clknet_4_13_0_clk),
    .D(_0091_),
    .Q(\buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1622_ (.CLK(clknet_4_13_0_clk),
    .D(_0092_),
    .Q(\buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1623_ (.CLK(clknet_4_12_0_clk),
    .D(_0093_),
    .Q(\buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1624_ (.CLK(clknet_4_12_0_clk),
    .D(_0094_),
    .Q(\buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1625_ (.CLK(clknet_4_13_0_clk),
    .D(_0095_),
    .Q(\buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1626_ (.CLK(clknet_4_12_0_clk),
    .D(_0096_),
    .Q(\buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1627_ (.CLK(clknet_4_13_0_clk),
    .D(_0097_),
    .Q(\buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1628_ (.CLK(clknet_4_11_0_clk),
    .D(_0098_),
    .Q(\buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1629_ (.CLK(clknet_4_9_0_clk),
    .D(_0099_),
    .Q(rd_valid));
 sky130_fd_sc_hd__dfxtp_1 _1630_ (.CLK(clknet_4_9_0_clk),
    .D(_0100_),
    .Q(rd_wait));
 sky130_fd_sc_hd__dfxtp_2 _1631_ (.CLK(clknet_4_12_0_clk),
    .D(_0101_),
    .Q(rd_inc));
 sky130_fd_sc_hd__dfxtp_1 _1632_ (.CLK(net128),
    .D(\xfer.flash_io0_do ),
    .Q(xfer_io0_90));
 sky130_fd_sc_hd__dfxtp_1 _1633_ (.CLK(net129),
    .D(\xfer.flash_io1_do ),
    .Q(xfer_io1_90));
 sky130_fd_sc_hd__dfxtp_1 _1634_ (.CLK(net130),
    .D(\xfer.flash_io2_do ),
    .Q(xfer_io2_90));
 sky130_fd_sc_hd__dfxtp_1 _1635_ (.CLK(net131),
    .D(\xfer.flash_io3_do ),
    .Q(xfer_io3_90));
 sky130_fd_sc_hd__dfxtp_4 _1636_ (.CLK(clknet_4_5_0_clk),
    .D(_0102_),
    .Q(config_en));
 sky130_fd_sc_hd__dfxtp_1 _1637_ (.CLK(clknet_4_7_0_clk),
    .D(_0103_),
    .Q(config_ddr));
 sky130_fd_sc_hd__dfxtp_2 _1638_ (.CLK(clknet_4_7_0_clk),
    .D(_0104_),
    .Q(config_qspi));
 sky130_fd_sc_hd__dfxtp_2 _1639_ (.CLK(clknet_4_7_0_clk),
    .D(_0105_),
    .Q(config_cont));
 sky130_fd_sc_hd__dfxtp_1 _1640_ (.CLK(clknet_4_5_0_clk),
    .D(_0106_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _1641_ (.CLK(clknet_4_5_0_clk),
    .D(_0107_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _1642_ (.CLK(clknet_4_7_0_clk),
    .D(_0108_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _1643_ (.CLK(clknet_4_7_0_clk),
    .D(_0109_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _1644_ (.CLK(clknet_4_5_0_clk),
    .D(_0110_),
    .Q(\config_oe[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1645_ (.CLK(clknet_4_5_0_clk),
    .D(_0111_),
    .Q(\config_oe[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1646_ (.CLK(clknet_4_5_0_clk),
    .D(_0112_),
    .Q(\config_oe[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1647_ (.CLK(clknet_4_5_0_clk),
    .D(_0113_),
    .Q(\config_oe[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1648_ (.CLK(clknet_4_5_0_clk),
    .D(_0114_),
    .Q(config_csb));
 sky130_fd_sc_hd__dfxtp_1 _1649_ (.CLK(clknet_4_5_0_clk),
    .D(_0115_),
    .Q(config_clk));
 sky130_fd_sc_hd__dfxtp_1 _1650_ (.CLK(clknet_4_5_0_clk),
    .D(_0116_),
    .Q(\config_do[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1651_ (.CLK(clknet_4_5_0_clk),
    .D(_0117_),
    .Q(\config_do[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1652_ (.CLK(clknet_4_5_0_clk),
    .D(_0118_),
    .Q(\config_do[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1653_ (.CLK(clknet_4_5_0_clk),
    .D(_0119_),
    .Q(\config_do[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1654_ (.CLK(clknet_4_3_0_clk),
    .D(_0000_),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1655_ (.CLK(clknet_4_7_0_clk),
    .D(_0004_),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1656_ (.CLK(clknet_4_6_0_clk),
    .D(_0005_),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1657_ (.CLK(clknet_4_3_0_clk),
    .D(_0006_),
    .Q(\state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1658_ (.CLK(clknet_4_7_0_clk),
    .D(_0007_),
    .Q(\state[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1659_ (.CLK(clknet_4_7_0_clk),
    .D(_0008_),
    .Q(\state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1660_ (.CLK(clknet_4_6_0_clk),
    .D(_0009_),
    .Q(\state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1661_ (.CLK(clknet_4_6_0_clk),
    .D(_0010_),
    .Q(\state[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1662_ (.CLK(clknet_4_7_0_clk),
    .D(_0011_),
    .Q(\state[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1663_ (.CLK(clknet_4_6_0_clk),
    .D(_0012_),
    .Q(\state[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1664_ (.CLK(clknet_4_7_0_clk),
    .D(_0001_),
    .Q(\state[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1665_ (.CLK(clknet_4_6_0_clk),
    .D(_0002_),
    .Q(\state[11] ));
 sky130_fd_sc_hd__dfxtp_2 _1666_ (.CLK(clknet_4_7_0_clk),
    .D(_0003_),
    .Q(\state[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1667_ (.CLK(clknet_4_5_0_clk),
    .D(_0120_),
    .Q(softreset));
 sky130_fd_sc_hd__dfxtp_1 _1668_ (.CLK(clknet_4_4_0_clk),
    .D(\xfer.xfer_ddr ),
    .Q(\xfer.xfer_ddr_q ));
 sky130_fd_sc_hd__dfxtp_1 _1669_ (.CLK(clknet_4_4_0_clk),
    .D(_0121_),
    .Q(\xfer.fetch ));
 sky130_fd_sc_hd__dfxtp_2 _1670_ (.CLK(clknet_4_10_0_clk),
    .D(_0122_),
    .Q(\xfer.dout_data[0] ));
 sky130_fd_sc_hd__dfxtp_4 _1671_ (.CLK(clknet_4_10_0_clk),
    .D(_0123_),
    .Q(\xfer.dout_data[1] ));
 sky130_fd_sc_hd__dfxtp_4 _1672_ (.CLK(clknet_4_10_0_clk),
    .D(_0124_),
    .Q(\xfer.dout_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1673_ (.CLK(clknet_4_10_0_clk),
    .D(_0125_),
    .Q(\xfer.dout_data[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1674_ (.CLK(clknet_4_10_0_clk),
    .D(_0126_),
    .Q(\xfer.dout_data[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1675_ (.CLK(clknet_4_10_0_clk),
    .D(_0127_),
    .Q(\xfer.dout_data[5] ));
 sky130_fd_sc_hd__dfxtp_2 _1676_ (.CLK(clknet_4_10_0_clk),
    .D(_0128_),
    .Q(\xfer.dout_data[6] ));
 sky130_fd_sc_hd__dfxtp_2 _1677_ (.CLK(clknet_4_10_0_clk),
    .D(_0129_),
    .Q(\xfer.dout_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1678_ (.CLK(clknet_4_12_0_clk),
    .D(\xfer.xfer_tag[0] ),
    .Q(\xfer.dout_tag[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1679_ (.CLK(clknet_4_9_0_clk),
    .D(\xfer.xfer_tag[1] ),
    .Q(\xfer.dout_tag[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1680_ (.CLK(clknet_4_12_0_clk),
    .D(\xfer.xfer_tag[2] ),
    .Q(\xfer.dout_tag[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1681_ (.CLK(clknet_4_4_0_clk),
    .D(_0130_),
    .Q(\xfer.xfer_rd ));
 sky130_fd_sc_hd__dfxtp_2 _1682_ (.CLK(clknet_4_4_0_clk),
    .D(_0131_),
    .Q(\xfer.xfer_qspi ));
 sky130_fd_sc_hd__dfxtp_2 _1683_ (.CLK(clknet_4_4_0_clk),
    .D(_0132_),
    .Q(\xfer.dummy_count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1684_ (.CLK(clknet_4_4_0_clk),
    .D(_0133_),
    .Q(\xfer.dummy_count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1685_ (.CLK(clknet_4_1_0_clk),
    .D(_0134_),
    .Q(\xfer.dummy_count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1686_ (.CLK(clknet_4_1_0_clk),
    .D(_0135_),
    .Q(\xfer.dummy_count[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1687_ (.CLK(clknet_4_0_0_clk),
    .D(_0136_),
    .Q(\xfer.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1688_ (.CLK(clknet_4_1_0_clk),
    .D(_0137_),
    .Q(\xfer.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1689_ (.CLK(clknet_4_6_0_clk),
    .D(_0138_),
    .Q(\xfer.din_tag[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1690_ (.CLK(clknet_4_3_0_clk),
    .D(_0139_),
    .Q(\xfer.din_tag[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1691_ (.CLK(clknet_4_6_0_clk),
    .D(_0140_),
    .Q(\xfer.din_tag[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1692_ (.CLK(clknet_4_4_0_clk),
    .D(_0141_),
    .Q(\xfer.xfer_ddr ));
 sky130_fd_sc_hd__dfxtp_2 _1693_ (.CLK(clknet_4_4_0_clk),
    .D(_0142_),
    .Q(\xfer.xfer_dspi ));
 sky130_fd_sc_hd__dfxtp_1 _1694_ (.CLK(clknet_4_4_0_clk),
    .D(_0143_),
    .Q(\xfer.flash_clk ));
 sky130_fd_sc_hd__dfxtp_1 _1695_ (.CLK(clknet_4_4_0_clk),
    .D(_0144_),
    .Q(\xfer.flash_csb ));
 sky130_fd_sc_hd__dfxtp_1 _1696_ (.CLK(clknet_4_13_0_clk),
    .D(_0145_),
    .Q(\rd_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1697_ (.CLK(clknet_4_13_0_clk),
    .D(_0146_),
    .Q(\rd_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1698_ (.CLK(clknet_4_2_0_clk),
    .D(_0147_),
    .Q(\rd_addr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1699_ (.CLK(clknet_4_2_0_clk),
    .D(_0148_),
    .Q(\rd_addr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1700_ (.CLK(clknet_4_2_0_clk),
    .D(_0149_),
    .Q(\rd_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1701_ (.CLK(clknet_4_2_0_clk),
    .D(_0150_),
    .Q(\rd_addr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _1702_ (.CLK(clknet_4_2_0_clk),
    .D(_0151_),
    .Q(\rd_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1703_ (.CLK(clknet_4_2_0_clk),
    .D(_0152_),
    .Q(\rd_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1704_ (.CLK(clknet_4_8_0_clk),
    .D(_0153_),
    .Q(\rd_addr[8] ));
 sky130_fd_sc_hd__dfxtp_2 _1705_ (.CLK(clknet_4_8_0_clk),
    .D(_0154_),
    .Q(\rd_addr[9] ));
 sky130_fd_sc_hd__dfxtp_2 _1706_ (.CLK(clknet_4_8_0_clk),
    .D(_0155_),
    .Q(\rd_addr[10] ));
 sky130_fd_sc_hd__dfxtp_2 _1707_ (.CLK(clknet_4_8_0_clk),
    .D(_0156_),
    .Q(\rd_addr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1708_ (.CLK(clknet_4_8_0_clk),
    .D(_0157_),
    .Q(\rd_addr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1709_ (.CLK(clknet_4_9_0_clk),
    .D(_0158_),
    .Q(\rd_addr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1710_ (.CLK(clknet_4_8_0_clk),
    .D(_0159_),
    .Q(\rd_addr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1711_ (.CLK(clknet_4_8_0_clk),
    .D(_0160_),
    .Q(\rd_addr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1712_ (.CLK(clknet_4_8_0_clk),
    .D(_0161_),
    .Q(\rd_addr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1713_ (.CLK(clknet_4_8_0_clk),
    .D(_0162_),
    .Q(\rd_addr[17] ));
 sky130_fd_sc_hd__dfxtp_2 _1714_ (.CLK(clknet_4_12_0_clk),
    .D(_0163_),
    .Q(\rd_addr[18] ));
 sky130_fd_sc_hd__dfxtp_2 _1715_ (.CLK(clknet_4_9_0_clk),
    .D(_0164_),
    .Q(\rd_addr[19] ));
 sky130_fd_sc_hd__dfxtp_2 _1716_ (.CLK(clknet_4_9_0_clk),
    .D(_0165_),
    .Q(\rd_addr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1717_ (.CLK(clknet_4_10_0_clk),
    .D(_0166_),
    .Q(\rd_addr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1718_ (.CLK(clknet_4_10_0_clk),
    .D(_0167_),
    .Q(\rd_addr[22] ));
 sky130_fd_sc_hd__dfxtp_2 _1719_ (.CLK(clknet_4_9_0_clk),
    .D(_0168_),
    .Q(\rd_addr[23] ));
 sky130_fd_sc_hd__dfxtp_2 _1720_ (.CLK(clknet_4_4_0_clk),
    .D(_0169_),
    .Q(\xfer.count[0] ));
 sky130_fd_sc_hd__conb_1 spimemio_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 spimemio_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 spimemio_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 spimemio_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 spimemio_119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 spimemio_120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 spimemio_121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 spimemio_122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 spimemio_123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 spimemio_124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 spimemio_125 (.LO(net125));
 sky130_fd_sc_hd__conb_1 spimemio_126 (.LO(net126));
 sky130_fd_sc_hd__conb_1 spimemio_127 (.LO(net127));
 sky130_fd_sc_hd__inv_2 _1294__1 (.A(clknet_4_0_0_clk),
    .Y(net128));
 sky130_fd_sc_hd__clkbuf_1 _1735_ (.A(net47),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 _1736_ (.A(net48),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 _1737_ (.A(net49),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _1738_ (.A(net50),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _1739_ (.A(net71),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _1740_ (.A(net72),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _1741_ (.A(net74),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _1742_ (.A(net76),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _1743_ (.A(net78),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 _1744_ (.A(net80),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 _1745_ (.A(config_cont),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _1746_ (.A(config_qspi),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _1747_ (.A(config_ddr),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _1748_ (.A(config_en),
    .X(net65));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3290 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(addr[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(addr[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(addr[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(addr[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(addr[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(addr[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(addr[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(addr[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(addr[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(addr[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(addr[19]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(addr[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(addr[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(addr[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(addr[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(addr[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(addr[2]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(addr[3]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(addr[4]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(addr[5]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(addr[6]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(addr[7]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(addr[8]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(addr[9]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(cfgreg_di[0]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(cfgreg_di[10]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(cfgreg_di[11]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(cfgreg_di[16]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(cfgreg_di[17]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(cfgreg_di[18]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(cfgreg_di[19]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(cfgreg_di[1]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(cfgreg_di[20]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(cfgreg_di[21]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(cfgreg_di[22]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(cfgreg_di[2]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(cfgreg_di[31]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(cfgreg_di[3]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(cfgreg_di[4]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(cfgreg_di[5]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(cfgreg_di[8]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(cfgreg_di[9]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(cfgreg_we[0]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(cfgreg_we[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(cfgreg_we[2]),
    .X(net45));
 sky130_fd_sc_hd__dlymetal6s2s_1 input46 (.A(cfgreg_we[3]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_8 input47 (.A(flash_io0_di),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_8 input48 (.A(flash_io1_di),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_8 input49 (.A(flash_io2_di),
    .X(net49));
 sky130_fd_sc_hd__buf_4 input50 (.A(flash_io3_di),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 input51 (.A(resetn),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(valid),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net53),
    .X(cfgreg_do[0]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net54),
    .X(cfgreg_do[10]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .X(cfgreg_do[11]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(cfgreg_do[16]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(cfgreg_do[17]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(cfgreg_do[18]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(cfgreg_do[19]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(cfgreg_do[1]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(cfgreg_do[20]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .X(cfgreg_do[21]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net63),
    .X(cfgreg_do[22]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net64),
    .X(cfgreg_do[2]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net65),
    .X(cfgreg_do[31]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(cfgreg_do[3]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(cfgreg_do[4]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(cfgreg_do[5]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .X(cfgreg_do[8]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(cfgreg_do[9]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .X(flash_clk));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .X(flash_csb));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .X(flash_io0_do));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net74),
    .X(flash_io0_oe));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .X(flash_io1_do));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net76),
    .X(flash_io1_oe));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net77),
    .X(flash_io2_do));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net78),
    .X(flash_io2_oe));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net79),
    .X(flash_io3_do));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net80),
    .X(flash_io3_oe));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net81),
    .X(rdata[0]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net82),
    .X(rdata[10]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net83),
    .X(rdata[11]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net84),
    .X(rdata[12]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net85),
    .X(rdata[13]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net86),
    .X(rdata[14]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net87),
    .X(rdata[15]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net88),
    .X(rdata[16]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net89),
    .X(rdata[17]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net90),
    .X(rdata[18]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net91),
    .X(rdata[19]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net92),
    .X(rdata[1]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net93),
    .X(rdata[20]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net94),
    .X(rdata[21]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net95),
    .X(rdata[22]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net96),
    .X(rdata[23]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net97),
    .X(rdata[24]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net98),
    .X(rdata[25]));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net99),
    .X(rdata[26]));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net100),
    .X(rdata[27]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net101),
    .X(rdata[28]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net102),
    .X(rdata[29]));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net103),
    .X(rdata[2]));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net104),
    .X(rdata[30]));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net105),
    .X(rdata[31]));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net106),
    .X(rdata[3]));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net107),
    .X(rdata[4]));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net108),
    .X(rdata[5]));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net109),
    .X(rdata[6]));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net110),
    .X(rdata[7]));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net111),
    .X(rdata[8]));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net112),
    .X(rdata[9]));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net113),
    .X(ready));
 sky130_fd_sc_hd__conb_1 spimemio_114 (.LO(net114));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 assign cfgreg_do[12] = net116;
 assign cfgreg_do[13] = net117;
 assign cfgreg_do[14] = net118;
 assign cfgreg_do[15] = net119;
 assign cfgreg_do[23] = net120;
 assign cfgreg_do[24] = net121;
 assign cfgreg_do[25] = net122;
 assign cfgreg_do[26] = net123;
 assign cfgreg_do[27] = net124;
 assign cfgreg_do[28] = net125;
 assign cfgreg_do[29] = net126;
 assign cfgreg_do[30] = net127;
 assign cfgreg_do[6] = net114;
 assign cfgreg_do[7] = net115;
endmodule
