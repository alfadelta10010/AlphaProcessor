VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alphasoc_mem
  CLASS BLOCK ;
  FOREIGN alphasoc_mem ;
  ORIGIN 0.000 0.000 ;
  SIZE 882.575 BY 893.295 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 881.520 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 881.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 881.520 ;
    END
  END VPWR
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 49.770 889.295 50.050 893.295 ;
    END
  END addr[0]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 889.295 146.650 893.295 ;
    END
  END addr[10]
  PIN addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 889.295 156.310 893.295 ;
    END
  END addr[11]
  PIN addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 889.295 165.970 893.295 ;
    END
  END addr[12]
  PIN addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 889.295 175.630 893.295 ;
    END
  END addr[13]
  PIN addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 889.295 185.290 893.295 ;
    END
  END addr[14]
  PIN addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 889.295 194.950 893.295 ;
    END
  END addr[15]
  PIN addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 889.295 204.610 893.295 ;
    END
  END addr[16]
  PIN addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 889.295 214.270 893.295 ;
    END
  END addr[17]
  PIN addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 889.295 223.930 893.295 ;
    END
  END addr[18]
  PIN addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 889.295 233.590 893.295 ;
    END
  END addr[19]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 59.430 889.295 59.710 893.295 ;
    END
  END addr[1]
  PIN addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 889.295 243.250 893.295 ;
    END
  END addr[20]
  PIN addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 889.295 252.910 893.295 ;
    END
  END addr[21]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 69.090 889.295 69.370 893.295 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 78.750 889.295 79.030 893.295 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 88.410 889.295 88.690 893.295 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 98.070 889.295 98.350 893.295 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 107.730 889.295 108.010 893.295 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 117.390 889.295 117.670 893.295 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 889.295 127.330 893.295 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 889.295 136.990 893.295 ;
    END
  END addr[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END clk
  PIN rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 571.410 889.295 571.690 893.295 ;
    END
  END rdata[0]
  PIN rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 668.010 889.295 668.290 893.295 ;
    END
  END rdata[10]
  PIN rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 677.670 889.295 677.950 893.295 ;
    END
  END rdata[11]
  PIN rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 687.330 889.295 687.610 893.295 ;
    END
  END rdata[12]
  PIN rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 696.990 889.295 697.270 893.295 ;
    END
  END rdata[13]
  PIN rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 706.650 889.295 706.930 893.295 ;
    END
  END rdata[14]
  PIN rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 716.310 889.295 716.590 893.295 ;
    END
  END rdata[15]
  PIN rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 725.970 889.295 726.250 893.295 ;
    END
  END rdata[16]
  PIN rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 735.630 889.295 735.910 893.295 ;
    END
  END rdata[17]
  PIN rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 745.290 889.295 745.570 893.295 ;
    END
  END rdata[18]
  PIN rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 754.950 889.295 755.230 893.295 ;
    END
  END rdata[19]
  PIN rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 581.070 889.295 581.350 893.295 ;
    END
  END rdata[1]
  PIN rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 764.610 889.295 764.890 893.295 ;
    END
  END rdata[20]
  PIN rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 774.270 889.295 774.550 893.295 ;
    END
  END rdata[21]
  PIN rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 783.930 889.295 784.210 893.295 ;
    END
  END rdata[22]
  PIN rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 793.590 889.295 793.870 893.295 ;
    END
  END rdata[23]
  PIN rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 803.250 889.295 803.530 893.295 ;
    END
  END rdata[24]
  PIN rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 812.910 889.295 813.190 893.295 ;
    END
  END rdata[25]
  PIN rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 822.570 889.295 822.850 893.295 ;
    END
  END rdata[26]
  PIN rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 832.230 889.295 832.510 893.295 ;
    END
  END rdata[27]
  PIN rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 841.890 889.295 842.170 893.295 ;
    END
  END rdata[28]
  PIN rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 851.550 889.295 851.830 893.295 ;
    END
  END rdata[29]
  PIN rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 590.730 889.295 591.010 893.295 ;
    END
  END rdata[2]
  PIN rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 861.210 889.295 861.490 893.295 ;
    END
  END rdata[30]
  PIN rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 870.870 889.295 871.150 893.295 ;
    END
  END rdata[31]
  PIN rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 600.390 889.295 600.670 893.295 ;
    END
  END rdata[3]
  PIN rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 610.050 889.295 610.330 893.295 ;
    END
  END rdata[4]
  PIN rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 619.710 889.295 619.990 893.295 ;
    END
  END rdata[5]
  PIN rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 629.370 889.295 629.650 893.295 ;
    END
  END rdata[6]
  PIN rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 639.030 889.295 639.310 893.295 ;
    END
  END rdata[7]
  PIN rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 648.690 889.295 648.970 893.295 ;
    END
  END rdata[8]
  PIN rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 658.350 889.295 658.630 893.295 ;
    END
  END rdata[9]
  PIN wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 262.290 889.295 262.570 893.295 ;
    END
  END wdata[0]
  PIN wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 358.890 889.295 359.170 893.295 ;
    END
  END wdata[10]
  PIN wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 368.550 889.295 368.830 893.295 ;
    END
  END wdata[11]
  PIN wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 378.210 889.295 378.490 893.295 ;
    END
  END wdata[12]
  PIN wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 387.870 889.295 388.150 893.295 ;
    END
  END wdata[13]
  PIN wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 397.530 889.295 397.810 893.295 ;
    END
  END wdata[14]
  PIN wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 407.190 889.295 407.470 893.295 ;
    END
  END wdata[15]
  PIN wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 416.850 889.295 417.130 893.295 ;
    END
  END wdata[16]
  PIN wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 426.510 889.295 426.790 893.295 ;
    END
  END wdata[17]
  PIN wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 436.170 889.295 436.450 893.295 ;
    END
  END wdata[18]
  PIN wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 445.830 889.295 446.110 893.295 ;
    END
  END wdata[19]
  PIN wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 271.950 889.295 272.230 893.295 ;
    END
  END wdata[1]
  PIN wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 455.490 889.295 455.770 893.295 ;
    END
  END wdata[20]
  PIN wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 465.150 889.295 465.430 893.295 ;
    END
  END wdata[21]
  PIN wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 474.810 889.295 475.090 893.295 ;
    END
  END wdata[22]
  PIN wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 484.470 889.295 484.750 893.295 ;
    END
  END wdata[23]
  PIN wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 494.130 889.295 494.410 893.295 ;
    END
  END wdata[24]
  PIN wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 503.790 889.295 504.070 893.295 ;
    END
  END wdata[25]
  PIN wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 513.450 889.295 513.730 893.295 ;
    END
  END wdata[26]
  PIN wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 523.110 889.295 523.390 893.295 ;
    END
  END wdata[27]
  PIN wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 532.770 889.295 533.050 893.295 ;
    END
  END wdata[28]
  PIN wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 542.430 889.295 542.710 893.295 ;
    END
  END wdata[29]
  PIN wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 281.610 889.295 281.890 893.295 ;
    END
  END wdata[2]
  PIN wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 552.090 889.295 552.370 893.295 ;
    END
  END wdata[30]
  PIN wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 561.750 889.295 562.030 893.295 ;
    END
  END wdata[31]
  PIN wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 291.270 889.295 291.550 893.295 ;
    END
  END wdata[3]
  PIN wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 300.930 889.295 301.210 893.295 ;
    END
  END wdata[4]
  PIN wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 310.590 889.295 310.870 893.295 ;
    END
  END wdata[5]
  PIN wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 320.250 889.295 320.530 893.295 ;
    END
  END wdata[6]
  PIN wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 329.910 889.295 330.190 893.295 ;
    END
  END wdata[7]
  PIN wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 339.570 889.295 339.850 893.295 ;
    END
  END wdata[8]
  PIN wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 349.230 889.295 349.510 893.295 ;
    END
  END wdata[9]
  PIN wen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 11.130 889.295 11.410 893.295 ;
    END
  END wen[0]
  PIN wen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 20.790 889.295 21.070 893.295 ;
    END
  END wen[1]
  PIN wen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 30.450 889.295 30.730 893.295 ;
    END
  END wen[2]
  PIN wen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 40.110 889.295 40.390 893.295 ;
    END
  END wen[3]
  OBS
      LAYER nwell ;
        RECT 5.330 877.145 876.950 879.975 ;
        RECT 5.330 871.705 876.950 874.535 ;
        RECT 5.330 866.265 876.950 869.095 ;
        RECT 5.330 860.825 876.950 863.655 ;
        RECT 5.330 855.385 876.950 858.215 ;
        RECT 5.330 849.945 876.950 852.775 ;
        RECT 5.330 844.505 876.950 847.335 ;
        RECT 5.330 839.065 876.950 841.895 ;
        RECT 5.330 833.625 876.950 836.455 ;
        RECT 5.330 828.185 876.950 831.015 ;
        RECT 5.330 822.745 876.950 825.575 ;
        RECT 5.330 817.305 876.950 820.135 ;
        RECT 5.330 811.865 876.950 814.695 ;
        RECT 5.330 806.425 876.950 809.255 ;
        RECT 5.330 800.985 876.950 803.815 ;
        RECT 5.330 795.545 876.950 798.375 ;
        RECT 5.330 790.105 876.950 792.935 ;
        RECT 5.330 784.665 876.950 787.495 ;
        RECT 5.330 779.225 876.950 782.055 ;
        RECT 5.330 773.785 876.950 776.615 ;
        RECT 5.330 768.345 876.950 771.175 ;
        RECT 5.330 762.905 876.950 765.735 ;
        RECT 5.330 757.465 876.950 760.295 ;
        RECT 5.330 752.025 876.950 754.855 ;
        RECT 5.330 746.585 876.950 749.415 ;
        RECT 5.330 741.145 876.950 743.975 ;
        RECT 5.330 735.705 876.950 738.535 ;
        RECT 5.330 730.265 876.950 733.095 ;
        RECT 5.330 724.825 876.950 727.655 ;
        RECT 5.330 719.385 876.950 722.215 ;
        RECT 5.330 713.945 876.950 716.775 ;
        RECT 5.330 708.505 876.950 711.335 ;
        RECT 5.330 703.065 876.950 705.895 ;
        RECT 5.330 697.625 876.950 700.455 ;
        RECT 5.330 692.185 876.950 695.015 ;
        RECT 5.330 686.745 876.950 689.575 ;
        RECT 5.330 681.305 876.950 684.135 ;
        RECT 5.330 675.865 876.950 678.695 ;
        RECT 5.330 670.425 876.950 673.255 ;
        RECT 5.330 664.985 876.950 667.815 ;
        RECT 5.330 659.545 876.950 662.375 ;
        RECT 5.330 654.105 876.950 656.935 ;
        RECT 5.330 648.665 876.950 651.495 ;
        RECT 5.330 643.225 876.950 646.055 ;
        RECT 5.330 637.785 876.950 640.615 ;
        RECT 5.330 632.345 876.950 635.175 ;
        RECT 5.330 626.905 876.950 629.735 ;
        RECT 5.330 621.465 876.950 624.295 ;
        RECT 5.330 616.025 876.950 618.855 ;
        RECT 5.330 610.585 876.950 613.415 ;
        RECT 5.330 605.145 876.950 607.975 ;
        RECT 5.330 599.705 876.950 602.535 ;
        RECT 5.330 594.265 876.950 597.095 ;
        RECT 5.330 588.825 876.950 591.655 ;
        RECT 5.330 583.385 876.950 586.215 ;
        RECT 5.330 577.945 876.950 580.775 ;
        RECT 5.330 572.505 876.950 575.335 ;
        RECT 5.330 567.065 876.950 569.895 ;
        RECT 5.330 561.625 876.950 564.455 ;
        RECT 5.330 556.185 876.950 559.015 ;
        RECT 5.330 550.745 876.950 553.575 ;
        RECT 5.330 545.305 876.950 548.135 ;
        RECT 5.330 539.865 876.950 542.695 ;
        RECT 5.330 534.425 876.950 537.255 ;
        RECT 5.330 528.985 876.950 531.815 ;
        RECT 5.330 523.545 876.950 526.375 ;
        RECT 5.330 518.105 876.950 520.935 ;
        RECT 5.330 512.665 876.950 515.495 ;
        RECT 5.330 507.225 876.950 510.055 ;
        RECT 5.330 501.785 876.950 504.615 ;
        RECT 5.330 496.345 876.950 499.175 ;
        RECT 5.330 490.905 876.950 493.735 ;
        RECT 5.330 485.465 876.950 488.295 ;
        RECT 5.330 480.025 876.950 482.855 ;
        RECT 5.330 474.585 876.950 477.415 ;
        RECT 5.330 469.145 876.950 471.975 ;
        RECT 5.330 463.705 876.950 466.535 ;
        RECT 5.330 458.265 876.950 461.095 ;
        RECT 5.330 452.825 876.950 455.655 ;
        RECT 5.330 447.385 876.950 450.215 ;
        RECT 5.330 441.945 876.950 444.775 ;
        RECT 5.330 436.505 876.950 439.335 ;
        RECT 5.330 431.065 876.950 433.895 ;
        RECT 5.330 425.625 876.950 428.455 ;
        RECT 5.330 420.185 876.950 423.015 ;
        RECT 5.330 414.745 876.950 417.575 ;
        RECT 5.330 409.305 876.950 412.135 ;
        RECT 5.330 403.865 876.950 406.695 ;
        RECT 5.330 398.425 876.950 401.255 ;
        RECT 5.330 392.985 876.950 395.815 ;
        RECT 5.330 387.545 876.950 390.375 ;
        RECT 5.330 382.105 876.950 384.935 ;
        RECT 5.330 376.665 876.950 379.495 ;
        RECT 5.330 371.225 876.950 374.055 ;
        RECT 5.330 365.785 876.950 368.615 ;
        RECT 5.330 360.345 876.950 363.175 ;
        RECT 5.330 354.905 876.950 357.735 ;
        RECT 5.330 349.465 876.950 352.295 ;
        RECT 5.330 344.025 876.950 346.855 ;
        RECT 5.330 338.585 876.950 341.415 ;
        RECT 5.330 333.145 876.950 335.975 ;
        RECT 5.330 327.705 876.950 330.535 ;
        RECT 5.330 322.265 876.950 325.095 ;
        RECT 5.330 316.825 876.950 319.655 ;
        RECT 5.330 311.385 876.950 314.215 ;
        RECT 5.330 305.945 876.950 308.775 ;
        RECT 5.330 300.505 876.950 303.335 ;
        RECT 5.330 295.065 876.950 297.895 ;
        RECT 5.330 289.625 876.950 292.455 ;
        RECT 5.330 284.185 876.950 287.015 ;
        RECT 5.330 278.745 876.950 281.575 ;
        RECT 5.330 273.305 876.950 276.135 ;
        RECT 5.330 267.865 876.950 270.695 ;
        RECT 5.330 262.425 876.950 265.255 ;
        RECT 5.330 256.985 876.950 259.815 ;
        RECT 5.330 251.545 876.950 254.375 ;
        RECT 5.330 246.105 876.950 248.935 ;
        RECT 5.330 240.665 876.950 243.495 ;
        RECT 5.330 235.225 876.950 238.055 ;
        RECT 5.330 229.785 876.950 232.615 ;
        RECT 5.330 224.345 876.950 227.175 ;
        RECT 5.330 218.905 876.950 221.735 ;
        RECT 5.330 213.465 876.950 216.295 ;
        RECT 5.330 208.025 876.950 210.855 ;
        RECT 5.330 202.585 876.950 205.415 ;
        RECT 5.330 197.145 876.950 199.975 ;
        RECT 5.330 191.705 876.950 194.535 ;
        RECT 5.330 186.265 876.950 189.095 ;
        RECT 5.330 180.825 876.950 183.655 ;
        RECT 5.330 175.385 876.950 178.215 ;
        RECT 5.330 169.945 876.950 172.775 ;
        RECT 5.330 164.505 876.950 167.335 ;
        RECT 5.330 159.065 876.950 161.895 ;
        RECT 5.330 153.625 876.950 156.455 ;
        RECT 5.330 148.185 876.950 151.015 ;
        RECT 5.330 142.745 876.950 145.575 ;
        RECT 5.330 137.305 876.950 140.135 ;
        RECT 5.330 131.865 876.950 134.695 ;
        RECT 5.330 126.425 876.950 129.255 ;
        RECT 5.330 120.985 876.950 123.815 ;
        RECT 5.330 115.545 876.950 118.375 ;
        RECT 5.330 110.105 876.950 112.935 ;
        RECT 5.330 104.665 876.950 107.495 ;
        RECT 5.330 99.225 876.950 102.055 ;
        RECT 5.330 93.785 876.950 96.615 ;
        RECT 5.330 88.345 876.950 91.175 ;
        RECT 5.330 82.905 876.950 85.735 ;
        RECT 5.330 77.465 876.950 80.295 ;
        RECT 5.330 72.025 876.950 74.855 ;
        RECT 5.330 66.585 876.950 69.415 ;
        RECT 5.330 61.145 876.950 63.975 ;
        RECT 5.330 55.705 876.950 58.535 ;
        RECT 5.330 50.265 876.950 53.095 ;
        RECT 5.330 44.825 876.950 47.655 ;
        RECT 5.330 39.385 876.950 42.215 ;
        RECT 5.330 33.945 876.950 36.775 ;
        RECT 5.330 28.505 876.950 31.335 ;
        RECT 5.330 23.065 876.950 25.895 ;
        RECT 5.330 17.625 876.950 20.455 ;
        RECT 5.330 12.185 876.950 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 876.760 881.365 ;
      LAYER met1 ;
        RECT 5.520 10.640 877.060 883.280 ;
      LAYER met2 ;
        RECT 7.000 889.015 10.850 889.850 ;
        RECT 11.690 889.015 20.510 889.850 ;
        RECT 21.350 889.015 30.170 889.850 ;
        RECT 31.010 889.015 39.830 889.850 ;
        RECT 40.670 889.015 49.490 889.850 ;
        RECT 50.330 889.015 59.150 889.850 ;
        RECT 59.990 889.015 68.810 889.850 ;
        RECT 69.650 889.015 78.470 889.850 ;
        RECT 79.310 889.015 88.130 889.850 ;
        RECT 88.970 889.015 97.790 889.850 ;
        RECT 98.630 889.015 107.450 889.850 ;
        RECT 108.290 889.015 117.110 889.850 ;
        RECT 117.950 889.015 126.770 889.850 ;
        RECT 127.610 889.015 136.430 889.850 ;
        RECT 137.270 889.015 146.090 889.850 ;
        RECT 146.930 889.015 155.750 889.850 ;
        RECT 156.590 889.015 165.410 889.850 ;
        RECT 166.250 889.015 175.070 889.850 ;
        RECT 175.910 889.015 184.730 889.850 ;
        RECT 185.570 889.015 194.390 889.850 ;
        RECT 195.230 889.015 204.050 889.850 ;
        RECT 204.890 889.015 213.710 889.850 ;
        RECT 214.550 889.015 223.370 889.850 ;
        RECT 224.210 889.015 233.030 889.850 ;
        RECT 233.870 889.015 242.690 889.850 ;
        RECT 243.530 889.015 252.350 889.850 ;
        RECT 253.190 889.015 262.010 889.850 ;
        RECT 262.850 889.015 271.670 889.850 ;
        RECT 272.510 889.015 281.330 889.850 ;
        RECT 282.170 889.015 290.990 889.850 ;
        RECT 291.830 889.015 300.650 889.850 ;
        RECT 301.490 889.015 310.310 889.850 ;
        RECT 311.150 889.015 319.970 889.850 ;
        RECT 320.810 889.015 329.630 889.850 ;
        RECT 330.470 889.015 339.290 889.850 ;
        RECT 340.130 889.015 348.950 889.850 ;
        RECT 349.790 889.015 358.610 889.850 ;
        RECT 359.450 889.015 368.270 889.850 ;
        RECT 369.110 889.015 377.930 889.850 ;
        RECT 378.770 889.015 387.590 889.850 ;
        RECT 388.430 889.015 397.250 889.850 ;
        RECT 398.090 889.015 406.910 889.850 ;
        RECT 407.750 889.015 416.570 889.850 ;
        RECT 417.410 889.015 426.230 889.850 ;
        RECT 427.070 889.015 435.890 889.850 ;
        RECT 436.730 889.015 445.550 889.850 ;
        RECT 446.390 889.015 455.210 889.850 ;
        RECT 456.050 889.015 464.870 889.850 ;
        RECT 465.710 889.015 474.530 889.850 ;
        RECT 475.370 889.015 484.190 889.850 ;
        RECT 485.030 889.015 493.850 889.850 ;
        RECT 494.690 889.015 503.510 889.850 ;
        RECT 504.350 889.015 513.170 889.850 ;
        RECT 514.010 889.015 522.830 889.850 ;
        RECT 523.670 889.015 532.490 889.850 ;
        RECT 533.330 889.015 542.150 889.850 ;
        RECT 542.990 889.015 551.810 889.850 ;
        RECT 552.650 889.015 561.470 889.850 ;
        RECT 562.310 889.015 571.130 889.850 ;
        RECT 571.970 889.015 580.790 889.850 ;
        RECT 581.630 889.015 590.450 889.850 ;
        RECT 591.290 889.015 600.110 889.850 ;
        RECT 600.950 889.015 609.770 889.850 ;
        RECT 610.610 889.015 619.430 889.850 ;
        RECT 620.270 889.015 629.090 889.850 ;
        RECT 629.930 889.015 638.750 889.850 ;
        RECT 639.590 889.015 648.410 889.850 ;
        RECT 649.250 889.015 658.070 889.850 ;
        RECT 658.910 889.015 667.730 889.850 ;
        RECT 668.570 889.015 677.390 889.850 ;
        RECT 678.230 889.015 687.050 889.850 ;
        RECT 687.890 889.015 696.710 889.850 ;
        RECT 697.550 889.015 706.370 889.850 ;
        RECT 707.210 889.015 716.030 889.850 ;
        RECT 716.870 889.015 725.690 889.850 ;
        RECT 726.530 889.015 735.350 889.850 ;
        RECT 736.190 889.015 745.010 889.850 ;
        RECT 745.850 889.015 754.670 889.850 ;
        RECT 755.510 889.015 764.330 889.850 ;
        RECT 765.170 889.015 773.990 889.850 ;
        RECT 774.830 889.015 783.650 889.850 ;
        RECT 784.490 889.015 793.310 889.850 ;
        RECT 794.150 889.015 802.970 889.850 ;
        RECT 803.810 889.015 812.630 889.850 ;
        RECT 813.470 889.015 822.290 889.850 ;
        RECT 823.130 889.015 831.950 889.850 ;
        RECT 832.790 889.015 841.610 889.850 ;
        RECT 842.450 889.015 851.270 889.850 ;
        RECT 852.110 889.015 860.930 889.850 ;
        RECT 861.770 889.015 870.590 889.850 ;
        RECT 871.430 889.015 875.280 889.850 ;
        RECT 7.000 4.280 875.280 889.015 ;
        RECT 7.000 4.000 440.490 4.280 ;
        RECT 441.330 4.000 875.280 4.280 ;
      LAYER met3 ;
        RECT 13.865 10.715 872.555 881.445 ;
      LAYER met4 ;
        RECT 31.575 19.895 97.440 880.425 ;
        RECT 99.840 19.895 174.240 880.425 ;
        RECT 176.640 19.895 251.040 880.425 ;
        RECT 253.440 19.895 327.840 880.425 ;
        RECT 330.240 19.895 404.640 880.425 ;
        RECT 407.040 19.895 481.440 880.425 ;
        RECT 483.840 19.895 558.240 880.425 ;
        RECT 560.640 19.895 635.040 880.425 ;
        RECT 637.440 19.895 711.840 880.425 ;
        RECT 714.240 19.895 788.640 880.425 ;
        RECT 791.040 19.895 837.825 880.425 ;
      LAYER met5 ;
        RECT 135.820 354.500 752.900 611.100 ;
  END
END alphasoc_mem
END LIBRARY

