magic
tech sky130A
magscale 1 2
timestamp 1701616863
<< nwell >>
rect 1066 175429 175390 175995
rect 1066 174341 175390 174907
rect 1066 173253 175390 173819
rect 1066 172165 175390 172731
rect 1066 171077 175390 171643
rect 1066 169989 175390 170555
rect 1066 168901 175390 169467
rect 1066 167813 175390 168379
rect 1066 166725 175390 167291
rect 1066 165637 175390 166203
rect 1066 164549 175390 165115
rect 1066 163461 175390 164027
rect 1066 162373 175390 162939
rect 1066 161285 175390 161851
rect 1066 160197 175390 160763
rect 1066 159109 175390 159675
rect 1066 158021 175390 158587
rect 1066 156933 175390 157499
rect 1066 155845 175390 156411
rect 1066 154757 175390 155323
rect 1066 153669 175390 154235
rect 1066 152581 175390 153147
rect 1066 151493 175390 152059
rect 1066 150405 175390 150971
rect 1066 149317 175390 149883
rect 1066 148229 175390 148795
rect 1066 147141 175390 147707
rect 1066 146053 175390 146619
rect 1066 144965 175390 145531
rect 1066 143877 175390 144443
rect 1066 142789 175390 143355
rect 1066 141701 175390 142267
rect 1066 140613 175390 141179
rect 1066 139525 175390 140091
rect 1066 138437 175390 139003
rect 1066 137349 175390 137915
rect 1066 136261 175390 136827
rect 1066 135173 175390 135739
rect 1066 134085 175390 134651
rect 1066 132997 175390 133563
rect 1066 131909 175390 132475
rect 1066 130821 175390 131387
rect 1066 129733 175390 130299
rect 1066 128645 175390 129211
rect 1066 127557 175390 128123
rect 1066 126469 175390 127035
rect 1066 125381 175390 125947
rect 1066 124293 175390 124859
rect 1066 123205 175390 123771
rect 1066 122117 175390 122683
rect 1066 121029 175390 121595
rect 1066 119941 175390 120507
rect 1066 118853 175390 119419
rect 1066 117765 175390 118331
rect 1066 116677 175390 117243
rect 1066 115589 175390 116155
rect 1066 114501 175390 115067
rect 1066 113413 175390 113979
rect 1066 112325 175390 112891
rect 1066 111237 175390 111803
rect 1066 110149 175390 110715
rect 1066 109061 175390 109627
rect 1066 107973 175390 108539
rect 1066 106885 175390 107451
rect 1066 105797 175390 106363
rect 1066 104709 175390 105275
rect 1066 103621 175390 104187
rect 1066 102533 175390 103099
rect 1066 101445 175390 102011
rect 1066 100357 175390 100923
rect 1066 99269 175390 99835
rect 1066 98181 175390 98747
rect 1066 97093 175390 97659
rect 1066 96005 175390 96571
rect 1066 94917 175390 95483
rect 1066 93829 175390 94395
rect 1066 92741 175390 93307
rect 1066 91653 175390 92219
rect 1066 90565 175390 91131
rect 1066 89477 175390 90043
rect 1066 88389 175390 88955
rect 1066 87301 175390 87867
rect 1066 86213 175390 86779
rect 1066 85125 175390 85691
rect 1066 84037 175390 84603
rect 1066 82949 175390 83515
rect 1066 81861 175390 82427
rect 1066 80773 175390 81339
rect 1066 79685 175390 80251
rect 1066 78597 175390 79163
rect 1066 77509 175390 78075
rect 1066 76421 175390 76987
rect 1066 75333 175390 75899
rect 1066 74245 175390 74811
rect 1066 73157 175390 73723
rect 1066 72069 175390 72635
rect 1066 70981 175390 71547
rect 1066 69893 175390 70459
rect 1066 68805 175390 69371
rect 1066 67717 175390 68283
rect 1066 66629 175390 67195
rect 1066 65541 175390 66107
rect 1066 64453 175390 65019
rect 1066 63365 175390 63931
rect 1066 62277 175390 62843
rect 1066 61189 175390 61755
rect 1066 60101 175390 60667
rect 1066 59013 175390 59579
rect 1066 57925 175390 58491
rect 1066 56837 175390 57403
rect 1066 55749 175390 56315
rect 1066 54661 175390 55227
rect 1066 53573 175390 54139
rect 1066 52485 175390 53051
rect 1066 51397 175390 51963
rect 1066 50309 175390 50875
rect 1066 49221 175390 49787
rect 1066 48133 175390 48699
rect 1066 47045 175390 47611
rect 1066 45957 175390 46523
rect 1066 44869 175390 45435
rect 1066 43781 175390 44347
rect 1066 42693 175390 43259
rect 1066 41605 175390 42171
rect 1066 40517 175390 41083
rect 1066 39429 175390 39995
rect 1066 38341 175390 38907
rect 1066 37253 175390 37819
rect 1066 36165 175390 36731
rect 1066 35077 175390 35643
rect 1066 33989 175390 34555
rect 1066 32901 175390 33467
rect 1066 31813 175390 32379
rect 1066 30725 175390 31291
rect 1066 29637 175390 30203
rect 1066 28549 175390 29115
rect 1066 27461 175390 28027
rect 1066 26373 175390 26939
rect 1066 25285 175390 25851
rect 1066 24197 175390 24763
rect 1066 23109 175390 23675
rect 1066 22021 175390 22587
rect 1066 20933 175390 21499
rect 1066 19845 175390 20411
rect 1066 18757 175390 19323
rect 1066 17669 175390 18235
rect 1066 16581 175390 17147
rect 1066 15493 175390 16059
rect 1066 14405 175390 14971
rect 1066 13317 175390 13883
rect 1066 12229 175390 12795
rect 1066 11141 175390 11707
rect 1066 10053 175390 10619
rect 1066 8965 175390 9531
rect 1066 7877 175390 8443
rect 1066 6789 175390 7355
rect 1066 5701 175390 6267
rect 1066 4613 175390 5179
rect 1066 3525 175390 4091
rect 1066 2437 175390 3003
<< obsli1 >>
rect 1104 2159 175352 176273
<< obsm1 >>
rect 1104 2128 175412 176656
<< metal2 >>
rect 2226 177859 2282 178659
rect 4158 177859 4214 178659
rect 6090 177859 6146 178659
rect 8022 177859 8078 178659
rect 9954 177859 10010 178659
rect 11886 177859 11942 178659
rect 13818 177859 13874 178659
rect 15750 177859 15806 178659
rect 17682 177859 17738 178659
rect 19614 177859 19670 178659
rect 21546 177859 21602 178659
rect 23478 177859 23534 178659
rect 25410 177859 25466 178659
rect 27342 177859 27398 178659
rect 29274 177859 29330 178659
rect 31206 177859 31262 178659
rect 33138 177859 33194 178659
rect 35070 177859 35126 178659
rect 37002 177859 37058 178659
rect 38934 177859 38990 178659
rect 40866 177859 40922 178659
rect 42798 177859 42854 178659
rect 44730 177859 44786 178659
rect 46662 177859 46718 178659
rect 48594 177859 48650 178659
rect 50526 177859 50582 178659
rect 52458 177859 52514 178659
rect 54390 177859 54446 178659
rect 56322 177859 56378 178659
rect 58254 177859 58310 178659
rect 60186 177859 60242 178659
rect 62118 177859 62174 178659
rect 64050 177859 64106 178659
rect 65982 177859 66038 178659
rect 67914 177859 67970 178659
rect 69846 177859 69902 178659
rect 71778 177859 71834 178659
rect 73710 177859 73766 178659
rect 75642 177859 75698 178659
rect 77574 177859 77630 178659
rect 79506 177859 79562 178659
rect 81438 177859 81494 178659
rect 83370 177859 83426 178659
rect 85302 177859 85358 178659
rect 87234 177859 87290 178659
rect 89166 177859 89222 178659
rect 91098 177859 91154 178659
rect 93030 177859 93086 178659
rect 94962 177859 95018 178659
rect 96894 177859 96950 178659
rect 98826 177859 98882 178659
rect 100758 177859 100814 178659
rect 102690 177859 102746 178659
rect 104622 177859 104678 178659
rect 106554 177859 106610 178659
rect 108486 177859 108542 178659
rect 110418 177859 110474 178659
rect 112350 177859 112406 178659
rect 114282 177859 114338 178659
rect 116214 177859 116270 178659
rect 118146 177859 118202 178659
rect 120078 177859 120134 178659
rect 122010 177859 122066 178659
rect 123942 177859 123998 178659
rect 125874 177859 125930 178659
rect 127806 177859 127862 178659
rect 129738 177859 129794 178659
rect 131670 177859 131726 178659
rect 133602 177859 133658 178659
rect 135534 177859 135590 178659
rect 137466 177859 137522 178659
rect 139398 177859 139454 178659
rect 141330 177859 141386 178659
rect 143262 177859 143318 178659
rect 145194 177859 145250 178659
rect 147126 177859 147182 178659
rect 149058 177859 149114 178659
rect 150990 177859 151046 178659
rect 152922 177859 152978 178659
rect 154854 177859 154910 178659
rect 156786 177859 156842 178659
rect 158718 177859 158774 178659
rect 160650 177859 160706 178659
rect 162582 177859 162638 178659
rect 164514 177859 164570 178659
rect 166446 177859 166502 178659
rect 168378 177859 168434 178659
rect 170310 177859 170366 178659
rect 172242 177859 172298 178659
rect 174174 177859 174230 178659
rect 88154 0 88210 800
<< obsm2 >>
rect 1400 177803 2170 177970
rect 2338 177803 4102 177970
rect 4270 177803 6034 177970
rect 6202 177803 7966 177970
rect 8134 177803 9898 177970
rect 10066 177803 11830 177970
rect 11998 177803 13762 177970
rect 13930 177803 15694 177970
rect 15862 177803 17626 177970
rect 17794 177803 19558 177970
rect 19726 177803 21490 177970
rect 21658 177803 23422 177970
rect 23590 177803 25354 177970
rect 25522 177803 27286 177970
rect 27454 177803 29218 177970
rect 29386 177803 31150 177970
rect 31318 177803 33082 177970
rect 33250 177803 35014 177970
rect 35182 177803 36946 177970
rect 37114 177803 38878 177970
rect 39046 177803 40810 177970
rect 40978 177803 42742 177970
rect 42910 177803 44674 177970
rect 44842 177803 46606 177970
rect 46774 177803 48538 177970
rect 48706 177803 50470 177970
rect 50638 177803 52402 177970
rect 52570 177803 54334 177970
rect 54502 177803 56266 177970
rect 56434 177803 58198 177970
rect 58366 177803 60130 177970
rect 60298 177803 62062 177970
rect 62230 177803 63994 177970
rect 64162 177803 65926 177970
rect 66094 177803 67858 177970
rect 68026 177803 69790 177970
rect 69958 177803 71722 177970
rect 71890 177803 73654 177970
rect 73822 177803 75586 177970
rect 75754 177803 77518 177970
rect 77686 177803 79450 177970
rect 79618 177803 81382 177970
rect 81550 177803 83314 177970
rect 83482 177803 85246 177970
rect 85414 177803 87178 177970
rect 87346 177803 89110 177970
rect 89278 177803 91042 177970
rect 91210 177803 92974 177970
rect 93142 177803 94906 177970
rect 95074 177803 96838 177970
rect 97006 177803 98770 177970
rect 98938 177803 100702 177970
rect 100870 177803 102634 177970
rect 102802 177803 104566 177970
rect 104734 177803 106498 177970
rect 106666 177803 108430 177970
rect 108598 177803 110362 177970
rect 110530 177803 112294 177970
rect 112462 177803 114226 177970
rect 114394 177803 116158 177970
rect 116326 177803 118090 177970
rect 118258 177803 120022 177970
rect 120190 177803 121954 177970
rect 122122 177803 123886 177970
rect 124054 177803 125818 177970
rect 125986 177803 127750 177970
rect 127918 177803 129682 177970
rect 129850 177803 131614 177970
rect 131782 177803 133546 177970
rect 133714 177803 135478 177970
rect 135646 177803 137410 177970
rect 137578 177803 139342 177970
rect 139510 177803 141274 177970
rect 141442 177803 143206 177970
rect 143374 177803 145138 177970
rect 145306 177803 147070 177970
rect 147238 177803 149002 177970
rect 149170 177803 150934 177970
rect 151102 177803 152866 177970
rect 153034 177803 154798 177970
rect 154966 177803 156730 177970
rect 156898 177803 158662 177970
rect 158830 177803 160594 177970
rect 160762 177803 162526 177970
rect 162694 177803 164458 177970
rect 164626 177803 166390 177970
rect 166558 177803 168322 177970
rect 168490 177803 170254 177970
rect 170422 177803 172186 177970
rect 172354 177803 174118 177970
rect 174286 177803 175056 177970
rect 1400 856 175056 177803
rect 1400 800 88098 856
rect 88266 800 175056 856
<< obsm3 >>
rect 2773 2143 174511 176289
<< metal4 >>
rect 4208 2128 4528 176304
rect 19568 2128 19888 176304
rect 34928 2128 35248 176304
rect 50288 2128 50608 176304
rect 65648 2128 65968 176304
rect 81008 2128 81328 176304
rect 96368 2128 96688 176304
rect 111728 2128 112048 176304
rect 127088 2128 127408 176304
rect 142448 2128 142768 176304
rect 157808 2128 158128 176304
rect 173168 2128 173488 176304
<< obsm4 >>
rect 6315 3979 19488 176085
rect 19968 3979 34848 176085
rect 35328 3979 50208 176085
rect 50688 3979 65568 176085
rect 66048 3979 80928 176085
rect 81408 3979 96288 176085
rect 96768 3979 111648 176085
rect 112128 3979 127008 176085
rect 127488 3979 142368 176085
rect 142848 3979 157728 176085
rect 158208 3979 167565 176085
<< obsm5 >>
rect 27164 70900 150580 122220
<< labels >>
rlabel metal4 s 19568 2128 19888 176304 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 176304 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 176304 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 176304 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 176304 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 176304 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 176304 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 176304 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 176304 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 176304 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 176304 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 176304 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 9954 177859 10010 178659 6 addr[0]
port 3 nsew signal input
rlabel metal2 s 29274 177859 29330 178659 6 addr[10]
port 4 nsew signal input
rlabel metal2 s 31206 177859 31262 178659 6 addr[11]
port 5 nsew signal input
rlabel metal2 s 33138 177859 33194 178659 6 addr[12]
port 6 nsew signal input
rlabel metal2 s 35070 177859 35126 178659 6 addr[13]
port 7 nsew signal input
rlabel metal2 s 37002 177859 37058 178659 6 addr[14]
port 8 nsew signal input
rlabel metal2 s 38934 177859 38990 178659 6 addr[15]
port 9 nsew signal input
rlabel metal2 s 40866 177859 40922 178659 6 addr[16]
port 10 nsew signal input
rlabel metal2 s 42798 177859 42854 178659 6 addr[17]
port 11 nsew signal input
rlabel metal2 s 44730 177859 44786 178659 6 addr[18]
port 12 nsew signal input
rlabel metal2 s 46662 177859 46718 178659 6 addr[19]
port 13 nsew signal input
rlabel metal2 s 11886 177859 11942 178659 6 addr[1]
port 14 nsew signal input
rlabel metal2 s 48594 177859 48650 178659 6 addr[20]
port 15 nsew signal input
rlabel metal2 s 50526 177859 50582 178659 6 addr[21]
port 16 nsew signal input
rlabel metal2 s 13818 177859 13874 178659 6 addr[2]
port 17 nsew signal input
rlabel metal2 s 15750 177859 15806 178659 6 addr[3]
port 18 nsew signal input
rlabel metal2 s 17682 177859 17738 178659 6 addr[4]
port 19 nsew signal input
rlabel metal2 s 19614 177859 19670 178659 6 addr[5]
port 20 nsew signal input
rlabel metal2 s 21546 177859 21602 178659 6 addr[6]
port 21 nsew signal input
rlabel metal2 s 23478 177859 23534 178659 6 addr[7]
port 22 nsew signal input
rlabel metal2 s 25410 177859 25466 178659 6 addr[8]
port 23 nsew signal input
rlabel metal2 s 27342 177859 27398 178659 6 addr[9]
port 24 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 clk
port 25 nsew signal input
rlabel metal2 s 114282 177859 114338 178659 6 rdata[0]
port 26 nsew signal output
rlabel metal2 s 133602 177859 133658 178659 6 rdata[10]
port 27 nsew signal output
rlabel metal2 s 135534 177859 135590 178659 6 rdata[11]
port 28 nsew signal output
rlabel metal2 s 137466 177859 137522 178659 6 rdata[12]
port 29 nsew signal output
rlabel metal2 s 139398 177859 139454 178659 6 rdata[13]
port 30 nsew signal output
rlabel metal2 s 141330 177859 141386 178659 6 rdata[14]
port 31 nsew signal output
rlabel metal2 s 143262 177859 143318 178659 6 rdata[15]
port 32 nsew signal output
rlabel metal2 s 145194 177859 145250 178659 6 rdata[16]
port 33 nsew signal output
rlabel metal2 s 147126 177859 147182 178659 6 rdata[17]
port 34 nsew signal output
rlabel metal2 s 149058 177859 149114 178659 6 rdata[18]
port 35 nsew signal output
rlabel metal2 s 150990 177859 151046 178659 6 rdata[19]
port 36 nsew signal output
rlabel metal2 s 116214 177859 116270 178659 6 rdata[1]
port 37 nsew signal output
rlabel metal2 s 152922 177859 152978 178659 6 rdata[20]
port 38 nsew signal output
rlabel metal2 s 154854 177859 154910 178659 6 rdata[21]
port 39 nsew signal output
rlabel metal2 s 156786 177859 156842 178659 6 rdata[22]
port 40 nsew signal output
rlabel metal2 s 158718 177859 158774 178659 6 rdata[23]
port 41 nsew signal output
rlabel metal2 s 160650 177859 160706 178659 6 rdata[24]
port 42 nsew signal output
rlabel metal2 s 162582 177859 162638 178659 6 rdata[25]
port 43 nsew signal output
rlabel metal2 s 164514 177859 164570 178659 6 rdata[26]
port 44 nsew signal output
rlabel metal2 s 166446 177859 166502 178659 6 rdata[27]
port 45 nsew signal output
rlabel metal2 s 168378 177859 168434 178659 6 rdata[28]
port 46 nsew signal output
rlabel metal2 s 170310 177859 170366 178659 6 rdata[29]
port 47 nsew signal output
rlabel metal2 s 118146 177859 118202 178659 6 rdata[2]
port 48 nsew signal output
rlabel metal2 s 172242 177859 172298 178659 6 rdata[30]
port 49 nsew signal output
rlabel metal2 s 174174 177859 174230 178659 6 rdata[31]
port 50 nsew signal output
rlabel metal2 s 120078 177859 120134 178659 6 rdata[3]
port 51 nsew signal output
rlabel metal2 s 122010 177859 122066 178659 6 rdata[4]
port 52 nsew signal output
rlabel metal2 s 123942 177859 123998 178659 6 rdata[5]
port 53 nsew signal output
rlabel metal2 s 125874 177859 125930 178659 6 rdata[6]
port 54 nsew signal output
rlabel metal2 s 127806 177859 127862 178659 6 rdata[7]
port 55 nsew signal output
rlabel metal2 s 129738 177859 129794 178659 6 rdata[8]
port 56 nsew signal output
rlabel metal2 s 131670 177859 131726 178659 6 rdata[9]
port 57 nsew signal output
rlabel metal2 s 52458 177859 52514 178659 6 wdata[0]
port 58 nsew signal input
rlabel metal2 s 71778 177859 71834 178659 6 wdata[10]
port 59 nsew signal input
rlabel metal2 s 73710 177859 73766 178659 6 wdata[11]
port 60 nsew signal input
rlabel metal2 s 75642 177859 75698 178659 6 wdata[12]
port 61 nsew signal input
rlabel metal2 s 77574 177859 77630 178659 6 wdata[13]
port 62 nsew signal input
rlabel metal2 s 79506 177859 79562 178659 6 wdata[14]
port 63 nsew signal input
rlabel metal2 s 81438 177859 81494 178659 6 wdata[15]
port 64 nsew signal input
rlabel metal2 s 83370 177859 83426 178659 6 wdata[16]
port 65 nsew signal input
rlabel metal2 s 85302 177859 85358 178659 6 wdata[17]
port 66 nsew signal input
rlabel metal2 s 87234 177859 87290 178659 6 wdata[18]
port 67 nsew signal input
rlabel metal2 s 89166 177859 89222 178659 6 wdata[19]
port 68 nsew signal input
rlabel metal2 s 54390 177859 54446 178659 6 wdata[1]
port 69 nsew signal input
rlabel metal2 s 91098 177859 91154 178659 6 wdata[20]
port 70 nsew signal input
rlabel metal2 s 93030 177859 93086 178659 6 wdata[21]
port 71 nsew signal input
rlabel metal2 s 94962 177859 95018 178659 6 wdata[22]
port 72 nsew signal input
rlabel metal2 s 96894 177859 96950 178659 6 wdata[23]
port 73 nsew signal input
rlabel metal2 s 98826 177859 98882 178659 6 wdata[24]
port 74 nsew signal input
rlabel metal2 s 100758 177859 100814 178659 6 wdata[25]
port 75 nsew signal input
rlabel metal2 s 102690 177859 102746 178659 6 wdata[26]
port 76 nsew signal input
rlabel metal2 s 104622 177859 104678 178659 6 wdata[27]
port 77 nsew signal input
rlabel metal2 s 106554 177859 106610 178659 6 wdata[28]
port 78 nsew signal input
rlabel metal2 s 108486 177859 108542 178659 6 wdata[29]
port 79 nsew signal input
rlabel metal2 s 56322 177859 56378 178659 6 wdata[2]
port 80 nsew signal input
rlabel metal2 s 110418 177859 110474 178659 6 wdata[30]
port 81 nsew signal input
rlabel metal2 s 112350 177859 112406 178659 6 wdata[31]
port 82 nsew signal input
rlabel metal2 s 58254 177859 58310 178659 6 wdata[3]
port 83 nsew signal input
rlabel metal2 s 60186 177859 60242 178659 6 wdata[4]
port 84 nsew signal input
rlabel metal2 s 62118 177859 62174 178659 6 wdata[5]
port 85 nsew signal input
rlabel metal2 s 64050 177859 64106 178659 6 wdata[6]
port 86 nsew signal input
rlabel metal2 s 65982 177859 66038 178659 6 wdata[7]
port 87 nsew signal input
rlabel metal2 s 67914 177859 67970 178659 6 wdata[8]
port 88 nsew signal input
rlabel metal2 s 69846 177859 69902 178659 6 wdata[9]
port 89 nsew signal input
rlabel metal2 s 2226 177859 2282 178659 6 wen[0]
port 90 nsew signal input
rlabel metal2 s 4158 177859 4214 178659 6 wen[1]
port 91 nsew signal input
rlabel metal2 s 6090 177859 6146 178659 6 wen[2]
port 92 nsew signal input
rlabel metal2 s 8022 177859 8078 178659 6 wen[3]
port 93 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 176515 178659
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 83613758
string GDS_FILE /openlane/designs/alphasoc_mem/runs/RUN_2023.12.03_14.26.22/results/signoff/alphasoc_mem.magic.gds
string GDS_START 351350
<< end >>

