* NGSPICE file created from alphacore.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

.subckt alphacore VGND VPWR clk cpi_insn[0] cpi_insn[10] cpi_insn[11] cpi_insn[12]
+ cpi_insn[13] cpi_insn[14] cpi_insn[1] cpi_insn[20] cpi_insn[21] cpi_insn[22] cpi_insn[23]
+ cpi_insn[24] cpi_insn[25] cpi_insn[26] cpi_insn[27] cpi_insn[28] cpi_insn[29] cpi_insn[2]
+ cpi_insn[30] cpi_insn[31] cpi_insn[3] cpi_insn[4] cpi_insn[5] cpi_insn[6] cpi_insn[7]
+ cpi_insn[8] cpi_insn[9] cpi_rs1[0] cpi_rs1[10] cpi_rs1[11] cpi_rs1[12] cpi_rs1[13]
+ cpi_rs1[14] cpi_rs1[15] cpi_rs1[16] cpi_rs1[17] cpi_rs1[18] cpi_rs1[19] cpi_rs1[1]
+ cpi_rs1[20] cpi_rs1[21] cpi_rs1[22] cpi_rs1[23] cpi_rs1[24] cpi_rs1[25] cpi_rs1[26]
+ cpi_rs1[27] cpi_rs1[28] cpi_rs1[29] cpi_rs1[2] cpi_rs1[30] cpi_rs1[31] cpi_rs1[3]
+ cpi_rs1[4] cpi_rs1[5] cpi_rs1[6] cpi_rs1[7] cpi_rs1[8] cpi_rs1[9] cpi_rs2[0] cpi_rs2[10]
+ cpi_rs2[11] cpi_rs2[12] cpi_rs2[13] cpi_rs2[14] cpi_rs2[15] cpi_rs2[16] cpi_rs2[17]
+ cpi_rs2[18] cpi_rs2[19] cpi_rs2[1] cpi_rs2[20] cpi_rs2[21] cpi_rs2[22] cpi_rs2[23]
+ cpi_rs2[24] cpi_rs2[25] cpi_rs2[26] cpi_rs2[27] cpi_rs2[28] cpi_rs2[29] cpi_rs2[2]
+ cpi_rs2[30] cpi_rs2[31] cpi_rs2[3] cpi_rs2[4] cpi_rs2[5] cpi_rs2[6] cpi_rs2[7] cpi_rs2[8]
+ cpi_rs2[9] cpi_valid cpi_wait eoi[0] eoi[10] eoi[11] eoi[12] eoi[13] eoi[14] eoi[15]
+ eoi[16] eoi[17] eoi[18] eoi[19] eoi[1] eoi[20] eoi[21] eoi[22] eoi[23] eoi[24] eoi[25]
+ eoi[26] eoi[27] eoi[28] eoi[29] eoi[2] eoi[30] eoi[31] eoi[3] eoi[4] eoi[5] eoi[6]
+ eoi[7] eoi[8] eoi[9] irq[0] irq[10] irq[11] irq[12] irq[13] irq[14] irq[15] irq[16]
+ irq[17] irq[18] irq[19] irq[1] irq[20] irq[21] irq[22] irq[23] irq[24] irq[25] irq[26]
+ irq[27] irq[28] irq[29] irq[2] irq[30] irq[31] irq[3] irq[4] irq[5] irq[6] irq[7]
+ irq[8] irq[9] mem_addr[10] mem_addr[11] mem_addr[12] mem_addr[13] mem_addr[14] mem_addr[15]
+ mem_addr[16] mem_addr[17] mem_addr[18] mem_addr[19] mem_addr[1] mem_addr[20] mem_addr[21]
+ mem_addr[22] mem_addr[23] mem_addr[24] mem_addr[25] mem_addr[26] mem_addr[27] mem_addr[28]
+ mem_addr[29] mem_addr[2] mem_addr[30] mem_addr[31] mem_addr[3] mem_addr[4] mem_addr[5]
+ mem_addr[6] mem_addr[7] mem_addr[8] mem_addr[9] mem_instr mem_la_addr[0] mem_la_addr[10]
+ mem_la_addr[11] mem_la_addr[12] mem_la_addr[13] mem_la_addr[14] mem_la_addr[15]
+ mem_la_addr[16] mem_la_addr[17] mem_la_addr[18] mem_la_addr[19] mem_la_addr[1] mem_la_addr[20]
+ mem_la_addr[21] mem_la_addr[22] mem_la_addr[23] mem_la_addr[24] mem_la_addr[25]
+ mem_la_addr[26] mem_la_addr[27] mem_la_addr[28] mem_la_addr[29] mem_la_addr[2] mem_la_addr[30]
+ mem_la_addr[31] mem_la_addr[3] mem_la_addr[4] mem_la_addr[5] mem_la_addr[6] mem_la_addr[7]
+ mem_la_addr[8] mem_la_addr[9] mem_la_read mem_la_wdata[0] mem_la_wdata[10] mem_la_wdata[11]
+ mem_la_wdata[12] mem_la_wdata[13] mem_la_wdata[14] mem_la_wdata[15] mem_la_wdata[16]
+ mem_la_wdata[17] mem_la_wdata[18] mem_la_wdata[19] mem_la_wdata[1] mem_la_wdata[20]
+ mem_la_wdata[21] mem_la_wdata[22] mem_la_wdata[23] mem_la_wdata[24] mem_la_wdata[25]
+ mem_la_wdata[26] mem_la_wdata[27] mem_la_wdata[28] mem_la_wdata[29] mem_la_wdata[2]
+ mem_la_wdata[30] mem_la_wdata[31] mem_la_wdata[3] mem_la_wdata[4] mem_la_wdata[5]
+ mem_la_wdata[6] mem_la_wdata[7] mem_la_wdata[8] mem_la_wdata[9] mem_la_write mem_la_wstrb[0]
+ mem_la_wstrb[1] mem_la_wstrb[2] mem_la_wstrb[3] mem_rdata[0] mem_rdata[10] mem_rdata[11]
+ mem_rdata[12] mem_rdata[13] mem_rdata[14] mem_rdata[15] mem_rdata[16] mem_rdata[17]
+ mem_rdata[18] mem_rdata[19] mem_rdata[1] mem_rdata[20] mem_rdata[21] mem_rdata[22]
+ mem_rdata[23] mem_rdata[24] mem_rdata[25] mem_rdata[26] mem_rdata[27] mem_rdata[28]
+ mem_rdata[29] mem_rdata[2] mem_rdata[30] mem_rdata[31] mem_rdata[3] mem_rdata[4]
+ mem_rdata[5] mem_rdata[6] mem_rdata[7] mem_rdata[8] mem_rdata[9] mem_ready mem_valid
+ mem_wdata[0] mem_wdata[10] mem_wdata[11] mem_wdata[12] mem_wdata[13] mem_wdata[14]
+ mem_wdata[15] mem_wdata[16] mem_wdata[17] mem_wdata[18] mem_wdata[19] mem_wdata[1]
+ mem_wdata[20] mem_wdata[21] mem_wdata[22] mem_wdata[23] mem_wdata[24] mem_wdata[25]
+ mem_wdata[26] mem_wdata[27] mem_wdata[28] mem_wdata[29] mem_wdata[2] mem_wdata[30]
+ mem_wdata[31] mem_wdata[3] mem_wdata[4] mem_wdata[5] mem_wdata[6] mem_wdata[7] mem_wdata[8]
+ mem_wdata[9] mem_wstrb[0] mem_wstrb[1] mem_wstrb[2] mem_wstrb[3] resetn trace_data[0]
+ trace_data[18] trace_data[19] trace_data[1] trace_data[20] trace_data[21] trace_data[22]
+ trace_data[23] trace_data[24] trace_data[25] trace_data[26] trace_data[27] trace_data[28]
+ trace_data[29] trace_data[2] trace_data[3] trace_data[4] trace_data[5] trace_data[6]
+ trace_data[7] trace_data[8] trace_data[9] trace_valid trap cpi_insn[17] cpi_insn[16]
+ cpi_insn[15] trace_data[10] trace_data[30] mem_addr[0] trace_data[17] trace_data[16]
+ trace_data[15] cpi_insn[19] trace_data[14] cpi_insn[18] trace_data[35] trace_data[13]
+ trace_data[34] trace_data[12] trace_data[33] trace_data[11] trace_data[32] trace_data[31]
XANTENNA__10669__A1 _04566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09523__A2 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09671_ cpuregs.regs\[0\]\[8\] cpuregs.regs\[1\]\[8\] cpuregs.regs\[2\]\[8\] cpuregs.regs\[3\]\[8\]
+ _04072_ _04074_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__mux4_1
XANTENNA__15057__B1 _03692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11834__S _06359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13615__A _03575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08622_ _03271_ _03392_ _03395_ _03396_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_143_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09812__B decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08709__A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14804__B1 _01723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11618__B1 _06065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08553_ irq_mask\[20\] irq_pending\[20\] VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_59_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08428__B _03213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11094__A1 _05219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08484_ _03260_ _03265_ _03266_ _03267_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__or4_1
XFILLER_0_119_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15455__S1 _02000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16021__A2 _02711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08791__A_N net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15780__A1 _06186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08444__A _03206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09105_ _03862_ _03863_ _03864_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__o21a_1
XANTENNA__15976__S _03635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09036_ mem_16bit_buffer\[6\] _03797_ _03727_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__mux2_2
XFILLER_0_103_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_68_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15277__A _02066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09275__A _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10452__S0 _04085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09938_ _04646_ _04650_ _04100_ _04658_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_70_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10214__A _04206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15724__B _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08948__S1 _03662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09869_ _04296_ _04577_ _04582_ _04591_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_29_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11900_ _06399_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15143__S0 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12880_ _06343_ cpuregs.regs\[6\]\[31\] _06905_ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__mux2_1
XANTENNA__08619__A irq_mask\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11831_ _06361_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _07952_ _08206_ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__nor2_1
X_11762_ reg_out\[27\] alu_out_q\[27\] _06069_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13501_ _07274_ _07318_ _07358_ _07232_ VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__a31o_1
XANTENNA__16012__A2 mem_rdata_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10832__A1 _05288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10713_ _03526_ _05410_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15446__S1 _01980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14481_ _08137_ _08144_ _07937_ VGND VGND VPWR VPWR _08145_ sky130_fd_sc_hd__mux2_1
XANTENNA__12575__S _06774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11693_ _06247_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__buf_2
XFILLER_0_82_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15220__B1 _02017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _02834_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__clkbuf_1
X_13432_ _04251_ _05259_ VGND VGND VPWR VPWR _07294_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10644_ _04466_ _04532_ _04566_ _04602_ _05264_ _05232_ VGND VGND VPWR VPWR _05346_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14574__A2 _07948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10045__C1 _04070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12585__A1 _06588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16151_ _02793_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__clkbuf_1
X_10575_ _05267_ _05270_ _05273_ _05276_ _05277_ _05278_ VGND VGND VPWR VPWR _05279_
+ sky130_fd_sc_hd__mux4_2
X_13363_ _04036_ decoded_imm\[0\] _07227_ _07228_ VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__and4_1
XFILLER_0_63_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09450__A1 _04052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15102_ _01959_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__buf_8
XANTENNA__10060__A2 _04021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12314_ _06635_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__clkbuf_1
X_16082_ compressed_instr _05974_ _06016_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13294_ _07174_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output179_A net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15033_ _05037_ _01885_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__nor2_1
X_12245_ cpuregs.regs\[24\]\[30\] _06596_ _06533_ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10899__A1 _05288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12176_ _06156_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11560__A2 _03322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08961__B1 _03675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11127_ _03434_ _05799_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__xor2_1
XANTENNA__15915__A _02610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16510__S _02979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16984_ clknet_leaf_169_clk _00158_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11058_ _03456_ _03582_ _03587_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__o21ai_1
X_15935_ mem_rdata_q\[0\] mem_rdata_q\[1\] VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__nand2_1
XANTENNA__15634__B _03237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11312__A2 _05929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13435__A _03524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10009_ _04231_ _04727_ _04082_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__a21oi_1
X_15866_ instr_blt _02618_ _02622_ _02623_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08529__A is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14817_ count_cycle\[40\] count_cycle\[41\] _01762_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__and3_1
X_17605_ clknet_leaf_2_clk _00774_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_18585_ clknet_leaf_10_clk _01650_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_15797_ instr_lb _03291_ _02582_ latched_is_lb VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__a22o_1
XANTENNA__09808__A3 _04531_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17536_ clknet_leaf_172_clk _00705_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14748_ count_cycle\[19\] _01715_ _01717_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10823__A1 _05219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12485__S _06726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17467_ clknet_leaf_109_clk _00636_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14679_ _03294_ _07971_ _08033_ VGND VGND VPWR VPWR _08326_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12025__A0 _06132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16418_ _02939_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14565__A2 _07950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17398_ clknet_leaf_98_clk _00567_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16349_ _06955_ cpuregs.regs\[16\]\[6\] _02896_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__mux2_1
XANTENNA__10587__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15514__A1 decoded_imm\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18019_ clknet_leaf_104_clk _00026_ VGND VGND VPWR VPWR irq_pending\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10733__S _05363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08711__B net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11000__A1 _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08952__B1 _03692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15817__A2 _06016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10034__A _04673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09723_ _04168_ _04447_ _04449_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__a21o_1
XANTENNA__11564__S _06086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09654_ _04051_ _04382_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09034__S _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08605_ _03277_ cpu_state\[0\] VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09585_ _04313_ _04314_ _04223_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08536_ reg_sh\[1\] reg_sh\[0\] VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__or2_2
XANTENNA__13461__C1 _07221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08467_ _03240_ _03250_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__nor2_1
XANTENNA__12395__S _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16702__A0 _06968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10360_ _05056_ _05060_ _04227_ _05068_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__a211o_4
XANTENNA__10673__S0 _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12319__A1 _06598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09019_ _03780_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__clkbuf_4
X_10291_ _04223_ _05001_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__or2_1
XANTENNA__08621__B _03387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12030_ _06468_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15269__B1 _01963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_151_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15735__A _02476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13981_ _07753_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14492__A1 _07934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15720_ _04702_ _02479_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__nand2_1
XANTENNA__13255__A _07153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12932_ _06975_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09594__S1 _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_166_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15651_ _03301_ _04187_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__and2_1
X_12863_ _06931_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_103_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _08254_ _08255_ VGND VGND VPWR VPWR _08256_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_1_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ clknet_leaf_138_clk _01435_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11814_ _06352_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__clkbuf_1
X_15582_ net119 _01905_ _02412_ _02413_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15992__A1 _06016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12794_ _06894_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__clkbuf_1
X_17321_ clknet_leaf_132_clk _00495_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15419__S1 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _07986_ _08185_ _07995_ VGND VGND VPWR VPWR _08193_ sky130_fd_sc_hd__a21o_1
X_11745_ reg_out\[25\] alu_out_q\[25\] _06069_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14086__A _03239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12007__A0 _06328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17252_ clknet_leaf_143_clk _00426_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10281__A2 _04012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15744__A1 _04909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14464_ decoded_imm_j\[13\] _07934_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11676_ _06232_ cpuregs.regs\[10\]\[17\] _06176_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16203_ _03218_ _02822_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13415_ _04198_ _05258_ VGND VGND VPWR VPWR _07278_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10627_ _05265_ _05268_ _05240_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__mux2_1
X_17183_ clknet_leaf_179_clk _00357_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14395_ _07921_ _08048_ VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16134_ _02784_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__clkbuf_1
X_13346_ _04037_ decoded_imm\[0\] _03311_ VGND VGND VPWR VPWR _07213_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_118_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10558_ net74 _04744_ _05229_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11649__S _06176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16065_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__buf_2
XANTENNA__09627__B decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13277_ _06963_ cpuregs.regs\[5\]\[10\] _07165_ VGND VGND VPWR VPWR _07166_ sky130_fd_sc_hd__mux2_1
X_10489_ _05192_ _05193_ _04223_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15016_ _04776_ _01885_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__nor2_1
X_12228_ _06585_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10416__S0 _04579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15645__A _03239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15355__S0 _01970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12159_ cpuregs.regs\[24\]\[2\] _06538_ _06534_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__mux2_1
XANTENNA__09065__D _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16967_ clknet_leaf_145_clk _00141_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__14483__A1 _08012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15918_ mem_rdata_q\[29\] mem_rdata_q\[31\] VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__nor2_1
X_16898_ clknet_leaf_29_clk _00043_ VGND VGND VPWR VPWR mem_rdata_q\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18637_ clknet_leaf_140_clk _01697_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_15849_ _03402_ _06006_ _03788_ _02609_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__o22a_1
XFILLER_0_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09370_ instr_rdcycleh VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__clkbuf_4
X_18568_ clknet_leaf_151_clk _01633_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15811__C _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12797__A1 _06584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17519_ clknet_leaf_145_clk _00688_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09662__A1 _04156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18499_ clknet_leaf_148_clk _01564_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13104__S _07068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10272__A2 _04049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12943__S _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16415__S _02932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10024__A2 _04014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput220 net220 VGND VGND VPWR VPWR mem_la_addr[6] sky130_fd_sc_hd__buf_1
XANTENNA__12244__A _06335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput231 net231 VGND VGND VPWR VPWR mem_la_wdata[15] sky130_fd_sc_hd__buf_1
Xoutput242 net242 VGND VGND VPWR VPWR mem_la_wdata[25] sky130_fd_sc_hd__clkbuf_1
Xoutput253 net253 VGND VGND VPWR VPWR mem_la_wdata[6] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput264 net264 VGND VGND VPWR VPWR mem_wdata[10] sky130_fd_sc_hd__clkbuf_1
Xoutput275 net275 VGND VGND VPWR VPWR mem_wdata[20] sky130_fd_sc_hd__clkbuf_1
XANTENNA__13774__S _05227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput286 net286 VGND VGND VPWR VPWR mem_wdata[30] sky130_fd_sc_hd__clkbuf_1
Xoutput297 net297 VGND VGND VPWR VPWR mem_wstrb[2] sky130_fd_sc_hd__buf_1
XFILLER_0_10_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09553__A _04283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15671__B1 _03240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09706_ cpuregs.regs\[4\]\[9\] cpuregs.regs\[5\]\[9\] cpuregs.regs\[6\]\[9\] cpuregs.regs\[7\]\[9\]
+ _04291_ _04292_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__mux4_1
XANTENNA__12485__A0 _06184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09637_ _04364_ _04365_ _04321_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09568_ cpuregs.regs\[28\]\[5\] cpuregs.regs\[29\]\[5\] cpuregs.regs\[30\]\[5\] cpuregs.regs\[31\]\[5\]
+ _04275_ _04278_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_65_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08519_ _03291_ _03283_ _03287_ instr_sh VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__a22o_1
XANTENNA__13985__B1 _06054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10638__S _05323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09499_ _04052_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__buf_6
XFILLER_0_154_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11323__A reg_next_pc\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11530_ _06071_ reg_next_pc\[2\] _03326_ _06072_ _06101_ VGND VGND VPWR VPWR _06102_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11461_ irq_mask\[19\] _06042_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__or2_1
XANTENNA__12853__S _06917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14634__A _07998_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13200_ _06955_ cpuregs.regs\[8\]\[6\] _07118_ VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10412_ _03384_ _05116_ _05117_ _05118_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__and4_1
X_14180_ _07890_ _07815_ _07891_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__and3b_1
X_11392_ _05998_ _05999_ _06001_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13131_ _07088_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__clkbuf_1
X_10343_ _05048_ _05051_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14162__B1 _07877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10274_ reg_pc\[25\] decoded_imm\[25\] VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__and2_1
X_13062_ _06953_ cpuregs.regs\[7\]\[5\] _07046_ VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__mux2_1
Xalphacore_304 VGND VGND VPWR VPWR alphacore_304/HI cpi_insn[2] sky130_fd_sc_hd__conb_1
Xalphacore_315 VGND VGND VPWR VPWR alphacore_315/HI cpi_insn[13] sky130_fd_sc_hd__conb_1
Xalphacore_326 VGND VGND VPWR VPWR alphacore_326/HI cpi_insn[24] sky130_fd_sc_hd__conb_1
XANTENNA__08916__B1 _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_337 VGND VGND VPWR VPWR alphacore_337/HI mem_la_addr[0] sky130_fd_sc_hd__conb_1
X_12013_ _06080_ _06385_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__nand2_4
X_17870_ clknet_leaf_88_clk _01039_ VGND VGND VPWR VPWR count_cycle\[15\] sky130_fd_sc_hd__dfxtp_1
Xalphacore_348 VGND VGND VPWR VPWR alphacore_348/HI trace_data[9] sky130_fd_sc_hd__conb_1
Xalphacore_359 VGND VGND VPWR VPWR alphacore_359/HI trace_data[20] sky130_fd_sc_hd__conb_1
XFILLER_0_100_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16821_ _06536_ cpuregs.regs\[14\]\[1\] _03152_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15662__B1 _02484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12476__A0 _06150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16752_ _03117_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__clkbuf_1
X_13964_ _03325_ _07727_ _07728_ net149 VGND VGND VPWR VPWR _07742_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_85_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15703_ timer\[12\] _02514_ _02475_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__a21oi_1
X_12915_ _06942_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__buf_6
XANTENNA_output211_A net211 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_915 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16683_ _06949_ cpuregs.regs\[19\]\[3\] _03076_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__mux2_1
X_13895_ _03322_ _07678_ _07682_ net158 VGND VGND VPWR VPWR _07694_ sky130_fd_sc_hd__a22o_1
XANTENNA__11932__S _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13713__A net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15634_ _07778_ _03237_ _02461_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__and3_1
X_18422_ clknet_leaf_188_clk _01487_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09910__B _04631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12846_ _06922_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08807__A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14528__B _07942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13976__B1 _07681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18353_ clknet_leaf_50_clk _01421_ VGND VGND VPWR VPWR reg_next_pc\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_173_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15565_ decoded_imm\[27\] _02216_ _02197_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__a21o_1
XANTENNA__13432__B _05259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12777_ _06885_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13440__A2 _05259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17304_ clknet_leaf_170_clk _00478_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14516_ decoded_imm_j\[17\] _07943_ VGND VGND VPWR VPWR _08177_ sky130_fd_sc_hd__nand2_1
X_11728_ _06252_ _03343_ _06253_ _06278_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15717__A1 _07441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18284_ clknet_leaf_8_clk _01352_ VGND VGND VPWR VPWR is_alu_reg_reg sky130_fd_sc_hd__dfxtp_1
X_15496_ _02332_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_155_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17235_ clknet_leaf_109_clk _00409_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14447_ decoded_imm_j\[12\] _07932_ VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12763__S _06869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11659_ _06217_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17166_ clknet_leaf_123_clk _00340_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08604__C1 _03272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14378_ _07995_ VGND VGND VPWR VPWR _08050_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16117_ _03218_ _03199_ _02676_ _02678_ _02775_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__o41a_1
X_13329_ cpuregs.regs\[20\]\[0\] cpuregs.regs\[21\]\[0\] cpuregs.regs\[22\]\[0\] cpuregs.regs\[23\]\[0\]
+ _04207_ _04208_ VGND VGND VPWR VPWR _07196_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_133_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17097_ clknet_leaf_142_clk _00271_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16142__A1 net226 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10962__B1 _05221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16048_ _03402_ decoded_imm_j\[12\] _03403_ _02612_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__a22o_1
XANTENNA__15350__C1 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08870_ _03635_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__buf_4
X_17999_ clknet_leaf_80_clk _01136_ VGND VGND VPWR VPWR irq_mask\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12003__S _06446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10031__B decoded_imm\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09883__A1 _03385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11842__S _06359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13623__A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09422_ _03317_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__buf_4
XANTENNA__11690__A1 alu_out_q\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08717__A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11117__S1 _05277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09353_ cpuregs.regs\[4\]\[1\] cpuregs.regs\[5\]\[1\] cpuregs.regs\[6\]\[1\] cpuregs.regs\[7\]\[1\]
+ _04085_ _04087_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13431__A2 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09284_ instr_maskirq VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_43_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14454__A _03364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08452__A _03196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10402__C1 _03301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16091__D _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16133__A1 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15567__S0 _01979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14144__B1 _07826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15892__B1 _02625_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10921__S _05390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09797__S1 _04277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10705__B1 _05356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08999_ _03759_ _03760_ _03230_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__mux2_1
XANTENNA__13009__S _07021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10961_ _05226_ _05334_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__nand2_2
XANTENNA__11130__A0 _05205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12700_ _06842_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13680_ net81 decoded_imm\[22\] VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__or2_1
XANTENNA__11681__A1 alu_out_q\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15947__A1 _04016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10892_ _05225_ _05569_ _05578_ _05581_ VGND VGND VPWR VPWR alu_out\[14\] sky130_fd_sc_hd__a211o_1
XANTENNA__15947__B2 _02669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12631_ _06805_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12149__A _06077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13422__A2 _04241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15896__C_N _02613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12630__A0 _06216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15350_ _02189_ _02191_ _02194_ _03683_ _02018_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__a221o_1
X_12562_ cpuregs.regs\[2\]\[15\] _06565_ _06763_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14301_ irq_pending\[8\] irq_pending\[9\] irq_pending\[10\] irq_pending\[11\] VGND
+ VGND VPWR VPWR _07978_ sky130_fd_sc_hd__or4_1
XFILLER_0_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11513_ _06078_ cpuregs.regs\[10\]\[0\] _06086_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15281_ cpuregs.regs\[24\]\[11\] cpuregs.regs\[25\]\[11\] cpuregs.regs\[26\]\[11\]
+ cpuregs.regs\[27\]\[11\] _02074_ _02075_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__mux4_1
XANTENNA__12583__S _06774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _06216_ cpuregs.regs\[28\]\[15\] _06726_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17020_ clknet_leaf_3_clk _00194_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14232_ reg_next_pc\[11\] _05834_ _07901_ _07929_ VGND VGND VPWR VPWR _07930_ sky130_fd_sc_hd__o211a_2
X_11444_ _06029_ irq_pending\[11\] _06039_ net3 VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15580__C1 _02027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14163_ _07879_ _07880_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11500__B _06065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15558__S0 _02069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11375_ _05960_ _03878_ _05966_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_78_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14135__B1 _07834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13114_ _07005_ cpuregs.regs\[7\]\[30\] _07045_ VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__mux2_1
X_10326_ _04052_ _05031_ _05035_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__a21oi_1
X_14094_ count_instr\[34\] _07828_ _07790_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15907__B mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output259_A net259 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _07042_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__clkbuf_1
X_17922_ clknet_leaf_26_clk _08391_ VGND VGND VPWR VPWR reg_out\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _04967_ _04968_ _04222_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__mux2_1
X_10188_ _04320_ _04901_ _04068_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__o21a_1
X_17853_ clknet_leaf_104_clk _01022_ VGND VGND VPWR VPWR reg_next_pc\[30\] sky130_fd_sc_hd__dfxtp_1
X_16804_ _03144_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10132__A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17784_ clknet_leaf_85_clk _00953_ VGND VGND VPWR VPWR count_instr\[55\] sky130_fd_sc_hd__dfxtp_1
X_14996_ _03303_ _04022_ _04447_ _01878_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__a31o_1
XANTENNA__09921__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13947_ _07730_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__clkbuf_1
X_16735_ _07001_ cpuregs.regs\[19\]\[28\] _03098_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__mux2_1
XANTENNA__13443__A _07211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11672__A1 alu_out_q\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15399__C1 _01968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16666_ _03070_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__clkbuf_1
X_13878_ _07681_ VGND VGND VPWR VPWR _07682_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_157_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18405_ clknet_leaf_138_clk _01470_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_15617_ cpuregs.regs\[4\]\[31\] cpuregs.regs\[5\]\[31\] cpuregs.regs\[6\]\[31\] cpuregs.regs\[7\]\[31\]
+ _02046_ _02047_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__mux4_1
X_12829_ _06913_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16597_ _06999_ cpuregs.regs\[18\]\[27\] _03026_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11424__A1 _06026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15548_ _01959_ _02373_ _02381_ _01933_ decoded_imm\[26\] VGND VGND VPWR VPWR _02382_
+ sky130_fd_sc_hd__a32o_2
X_18336_ clknet_leaf_37_clk _01404_ VGND VGND VPWR VPWR mem_16bit_buffer\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09712__S1 _04219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08971__S _03730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18267_ clknet_leaf_26_clk _01338_ VGND VGND VPWR VPWR decoded_imm\[25\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_112_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_150_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_150_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__12493__S _06726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15479_ _03709_ _02315_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17218_ clknet_leaf_185_clk _00392_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18198_ clknet_leaf_43_clk _01269_ VGND VGND VPWR VPWR instr_slti sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17149_ clknet_leaf_2_clk _00323_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10307__A reg_pc\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09971_ cpuregs.regs\[16\]\[16\] cpuregs.regs\[17\]\[16\] cpuregs.regs\[18\]\[16\]
+ cpuregs.regs\[19\]\[16\] _04477_ _04478_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15309__S _01984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08922_ cpuregs.regs\[12\]\[3\] cpuregs.regs\[13\]\[3\] cpuregs.regs\[14\]\[3\] cpuregs.regs\[15\]\[3\]
+ _03641_ _03684_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__mux4_1
X_08853_ _03617_ _03618_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08784_ net129 VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09305__A0 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12668__S _06825_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11112__B1 _05517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09400__S0 _04123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10466__A2 _05170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11663__A1 alu_out_q\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10010__S1 _04478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12860__A0 _06266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09405_ cpuregs.regs\[8\]\[2\] cpuregs.regs\[9\]\[2\] cpuregs.regs\[10\]\[2\] cpuregs.regs\[11\]\[2\]
+ _04123_ _04058_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09336_ _00069_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11415__A1 _03892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09267_ _03737_ _03996_ _04004_ _03853_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_141_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_141_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11601__A _06165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09198_ _03730_ _03867_ _03848_ _03829_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10077__S1 _04284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16603__S _03003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08595__A1 _03309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11160_ net127 net113 _04668_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08910__A _03674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10111_ cpuregs.regs\[8\]\[20\] cpuregs.regs\[9\]\[20\] cpuregs.regs\[10\]\[20\]
+ cpuregs.regs\[11\]\[20\] _04275_ _04278_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__mux4_1
X_11091_ _03442_ _05220_ _05251_ _05765_ _05766_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__a221o_1
XANTENNA__10651__S _05287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09725__B decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ cpuregs.regs\[16\]\[18\] cpuregs.regs\[17\]\[18\] cpuregs.regs\[18\]\[18\]
+ cpuregs.regs\[19\]\[18\] _04758_ _04759_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_73_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13340__A1 _04215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10154__A1 _04483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12151__B cpuregs.waddr\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15743__A _07778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14850_ _01786_ _01787_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13801_ _05143_ _07236_ _07593_ _07238_ VGND VGND VPWR VPWR _07638_ sky130_fd_sc_hd__o211a_1
X_14781_ _01739_ _01740_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__nor2_1
XANTENNA__11103__B1 _05213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09847__A1 _04391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11993_ _06274_ cpuregs.regs\[21\]\[22\] _06446_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__mux2_1
XANTENNA__14359__A _03378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16520_ _02993_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13732_ _04959_ _07236_ _07530_ _07238_ VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__o211a_1
XANTENNA__09460__B decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10944_ _05627_ _05629_ _05390_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__mux2_1
XANTENNA__11654__A1 alu_out_q\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16451_ _06989_ cpuregs.regs\[29\]\[22\] _02954_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13663_ _07507_ _07509_ _07225_ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__a21bo_1
X_10875_ _05478_ _05554_ _05556_ _05565_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15402_ _02242_ _02243_ _03719_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__mux2_1
XANTENNA__10209__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12614_ _06796_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12603__A0 _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16382_ _02920_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__clkbuf_1
X_13594_ net74 decoded_imm\[16\] VGND VGND VPWR VPWR _07445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18121_ clknet_leaf_55_clk _01225_ VGND VGND VPWR VPWR latched_branch sky130_fd_sc_hd__dfxtp_4
XFILLER_0_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15333_ _02177_ _02178_ _02002_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12545_ cpuregs.regs\[2\]\[7\] _06548_ _06752_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_132_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_132_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13202__S _07118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18052_ clknet_leaf_52_clk _01157_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_108_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15264_ cpuregs.regs\[20\]\[10\] cpuregs.regs\[21\]\[10\] cpuregs.regs\[22\]\[10\]
+ cpuregs.regs\[23\]\[10\] _02022_ _02023_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__mux4_1
XFILLER_0_123_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12476_ _06150_ cpuregs.regs\[28\]\[7\] _06715_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17003_ clknet_leaf_154_clk _00177_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11230__B _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14215_ _05856_ _06134_ VGND VGND VPWR VPWR _07918_ sky130_fd_sc_hd__or2_1
XANTENNA__15918__A mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_5 _01992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11427_ irq_mask\[3\] _06030_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__or2_1
X_15195_ cpuregs.regs\[8\]\[7\] cpuregs.regs\[9\]\[7\] cpuregs.regs\[10\]\[7\] cpuregs.regs\[11\]\[7\]
+ _02046_ _02047_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__mux4_1
XANTENNA__10917__B1 _05334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08586__A1 _03298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output86_A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14146_ count_instr\[50\] count_instr\[49\] VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__and2_1
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11358_ cpuregs.raddr2\[0\] _03636_ _05968_ _05972_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10309_ _04984_ _04987_ _04985_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10561__S _05264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15320__A2 _02009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14077_ count_instr\[29\] _07818_ _07775_ VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__a21oi_1
X_11289_ _03575_ _05829_ _05914_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__o21ai_4
XFILLER_0_67_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17905_ clknet_leaf_88_clk _01074_ VGND VGND VPWR VPWR count_cycle\[50\] sky130_fd_sc_hd__dfxtp_1
X_13028_ cpuregs.regs\[3\]\[21\] _06578_ _07032_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__mux2_1
XANTENNA__15653__A _02476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17836_ clknet_leaf_59_clk _01005_ VGND VGND VPWR VPWR reg_next_pc\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17767_ clknet_leaf_94_clk _00936_ VGND VGND VPWR VPWR count_instr\[38\] sky130_fd_sc_hd__dfxtp_1
X_14979_ irq_mask\[2\] _01864_ _01868_ _08335_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11645__A1 alu_out_q\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16718_ _03075_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__buf_6
XANTENNA__09933__S1 _04469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17698_ clknet_leaf_75_clk _00867_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16649_ _03061_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_106_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09121_ _03783_ _03213_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__nor2_2
XFILLER_0_123_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18319_ clknet_leaf_37_clk _01387_ VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_123_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_123_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08714__B net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13112__S _07068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11421__A _03305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09052_ mem_16bit_buffer\[2\] _03813_ _03728_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16423__S _02932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09774__B1 _04468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11008__S0 _05264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09954_ _03638_ _04642_ _04664_ _03302_ _04674_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_55_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08905_ _03669_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__buf_6
XANTENNA__10136__A1 _03303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09885_ reg_pc\[14\] decoded_imm\[14\] VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__xnor2_1
X_08836_ instr_bge VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16272__A0 _06947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15075__B2 _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09561__A _04276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08767_ net121 net89 VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__nand2_1
XANTENNA__15170__S1 _02023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10500__A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08698_ net111 net79 VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10660_ _05225_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08905__A _03669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09319_ _04053_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10646__S _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10591_ _03524_ net95 _03518_ _03510_ _05264_ _05235_ VGND VGND VPWR VPWR _05294_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_134_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_114_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_114_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_90_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12330_ cpuregs.regs\[26\]\[3\] _06540_ _06641_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__mux2_1
XANTENNA__14338__B1 _07905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12261_ cpuregs.regs\[25\]\[3\] _06540_ _06604_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14642__A _07966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14000_ count_instr\[5\] count_instr\[4\] count_instr\[3\] _07761_ VGND VGND VPWR
+ VPWR _07767_ sky130_fd_sc_hd__and4_1
XFILLER_0_160_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13561__A1 _03275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11212_ reg_next_pc\[8\] reg_out\[8\] _05834_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09765__B1 _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12192_ _06200_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__buf_2
XANTENNA__09860__S0 _04487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11143_ _03407_ _05414_ net101 _04422_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__a22o_2
Xoutput75 net75 VGND VGND VPWR VPWR cpi_rs1[17] sky130_fd_sc_hd__clkbuf_1
Xoutput86 net86 VGND VGND VPWR VPWR cpi_rs1[27] sky130_fd_sc_hd__buf_1
Xoutput97 net97 VGND VGND VPWR VPWR cpi_rs1[8] sky130_fd_sc_hd__buf_1
X_11074_ _05600_ _05645_ _05745_ _05748_ _05750_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__a2111o_1
X_15951_ instr_fence _02617_ _02636_ _02672_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__a22o_1
XANTENNA__10127__B2 _04024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10025_ net75 VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__clkbuf_4
X_14902_ _01825_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10222__S1 _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15882_ _02634_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__buf_4
XANTENNA__16263__B1 _03292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13077__A0 _06968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17621_ clknet_leaf_100_clk _00790_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14833_ count_cycle\[46\] _01774_ _01717_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__a21oi_1
XANTENNA_output124_A net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15161__S1 _02014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14764_ count_cycle\[22\] count_cycle\[23\] count_cycle\[24\] _01722_ VGND VGND VPWR
+ VPWR _01729_ sky130_fd_sc_hd__and4_2
XANTENNA__12101__S _06496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17552_ clknet_leaf_130_clk _00721_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _06208_ cpuregs.regs\[21\]\[14\] _06435_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13715_ _07554_ _07557_ VGND VGND VPWR VPWR _07558_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_123_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _02984_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__clkbuf_1
X_10927_ _03484_ _05613_ _05517_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17483_ clknet_leaf_126_clk _00652_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14695_ _08337_ _07815_ _08338_ VGND VGND VPWR VPWR _08339_ sky130_fd_sc_hd__and3b_1
XANTENNA__16508__S _02979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13646_ _04810_ _07271_ _07487_ _07493_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__o22a_1
X_16434_ _06972_ cpuregs.regs\[29\]\[14\] _02943_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10858_ _03499_ _03556_ _03557_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10850__A2 _05357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15774__C1 _02476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09679__S0 _04085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16365_ _02911_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__clkbuf_1
X_13577_ _07422_ _07423_ _07427_ _07429_ VGND VGND VPWR VPWR _07430_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_105_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_105_clk sky130_fd_sc_hd__clkbuf_2
X_10789_ _05483_ _05416_ _05295_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18104_ clknet_leaf_90_clk _01208_ VGND VGND VPWR VPWR timer\[19\] sky130_fd_sc_hd__dfxtp_1
X_15316_ cpuregs.regs\[0\]\[13\] cpuregs.regs\[1\]\[13\] cpuregs.regs\[2\]\[13\] cpuregs.regs\[3\]\[13\]
+ _01985_ _01986_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__mux4_1
XFILLER_0_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12528_ cpuregs.waddr\[2\] cpuregs.waddr\[4\] cpuregs.waddr\[3\] _06083_ VGND VGND
+ VPWR VPWR _06750_ sky130_fd_sc_hd__or4b_4
XFILLER_0_125_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16296_ _02874_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18035_ clknet_leaf_66_clk _00011_ VGND VGND VPWR VPWR irq_pending\[19\] sky130_fd_sc_hd__dfxtp_1
X_15247_ _02020_ _02089_ _02097_ _01960_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__o211a_4
XTAP_TAPCELL_ROW_10_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12459_ _06081_ _06082_ _06384_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__and3_4
XFILLER_0_169_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15870__A_N _02612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09756__B1 _04082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15178_ cpuregs.regs\[0\]\[6\] cpuregs.regs\[1\]\[6\] cpuregs.regs\[2\]\[6\] cpuregs.regs\[3\]\[6\]
+ _02030_ _02031_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__mux4_1
XANTENNA__09851__S0 _04512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15829__B1 _03910_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14129_ _07856_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_165_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09508__B1 _04227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10669__A2 _04602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09670_ cpuregs.regs\[4\]\[8\] cpuregs.regs\[5\]\[8\] cpuregs.regs\[6\]\[8\] cpuregs.regs\[7\]\[8\]
+ _04072_ _04074_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15057__A1 _03657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08621_ is_slli_srli_srai _03387_ is_jalr_addi_slti_sltiu_xori_ori_andi VGND VGND
+ VPWR VPWR _03396_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_143_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17819_ clknet_leaf_66_clk _00988_ VGND VGND VPWR VPWR reg_pc\[27\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_143_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08552_ irq_mask\[31\] irq_pending\[31\] VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10826__C1 _05390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08483_ instr_srli instr_lhu instr_sb instr_lw VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08725__A net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15780__A2 _03298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12247__A _06342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09104_ _03814_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09035_ _03795_ _03796_ _03231_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09556__A _04065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10452__S1 _04087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09937_ _04483_ _04653_ _04657_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_70_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17923__D _08394_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15293__A _01984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09868_ _04133_ _04590_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__nand2_1
XANTENNA__16245__A0 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ net115 net83 VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__and2b_1
X_09799_ _04289_ _04523_ _04225_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__a21o_1
XANTENNA__15143__S1 _01997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08619__B irq_active VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13017__S _07021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11830_ _06184_ cpuregs.regs\[11\]\[11\] _06359_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11761_ _06306_ _06118_ _06307_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_68_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16328__S _02881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13500_ _04602_ _07276_ VGND VGND VPWR VPWR _07358_ sky130_fd_sc_hd__or2_1
XANTENNA__13541__A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10712_ _03526_ _05410_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__or2_1
XANTENNA__10293__B1 _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14480_ _07986_ _08136_ _07994_ VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__a21o_1
X_11692_ _06226_ reg_next_pc\[19\] _06244_ _06246_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__a211o_2
XANTENNA__15220__A1 _02012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13431_ _04251_ _07271_ _07286_ _07293_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_101_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10643_ _05331_ _05344_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16150_ net268 net230 _02786_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__mux2_1
X_13362_ net78 decoded_imm\[1\] VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10574_ _03530_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10596__A1 _05288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11793__A0 _06336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10140__S0 _04282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15101_ _01958_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__buf_4
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12313_ cpuregs.regs\[25\]\[28\] _06592_ _06626_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__mux2_1
XANTENNA__12591__S _06774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15468__A _01984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16081_ decoded_imm\[31\] _02750_ _02745_ mem_rdata_q\[31\] _02748_ VGND VGND VPWR
+ VPWR _01344_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13293_ _06980_ cpuregs.regs\[5\]\[18\] _07165_ VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15032_ _03303_ _04022_ _05009_ _01898_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12244_ _06335_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__buf_2
XFILLER_0_122_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14091__B _07815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09833__S0 _04071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12175_ _06549_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11126_ _05517_ _03436_ _05796_ _05798_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__o31a_1
XANTENNA__13298__A0 _06984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output241_A net241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16983_ clknet_leaf_163_clk _00157_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_11057_ _05600_ _05635_ _05728_ _05732_ _05734_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__a2111o_1
X_15934_ mem_rdata_q\[2\] mem_rdata_q\[18\] mem_rdata_q\[3\] mem_rdata_q\[19\] VGND
+ VGND VPWR VPWR _02660_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_108_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10008_ _04725_ _04726_ _04078_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13435__B decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ _02612_ _02613_ _03940_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__nor3b_2
XTAP_TAPCELL_ROW_88_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17604_ clknet_leaf_7_clk _00773_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14816_ count_cycle\[40\] _01762_ _01764_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18584_ clknet_leaf_189_clk _01649_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15796_ instr_lh _03291_ _02582_ latched_is_lh VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17535_ clknet_leaf_163_clk _00704_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14747_ _03239_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__clkbuf_4
X_11959_ _06141_ cpuregs.regs\[21\]\[6\] _06424_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14547__A _07943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17466_ clknet_leaf_112_clk _00635_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_14678_ _08319_ _08320_ _08325_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08545__A _03320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13629_ _04611_ _04913_ _05258_ VGND VGND VPWR VPWR _07478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16417_ _06955_ cpuregs.regs\[29\]\[6\] _02932_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17397_ clknet_leaf_101_clk _00566_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16348_ _02902_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10587__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11784__A0 _06328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15378__A _03658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16279_ _02865_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15514__A2 _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15809__C _03864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13525__A1 _04466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09376__A _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18018_ clknet_leaf_64_clk _00023_ VGND VGND VPWR VPWR irq_pending\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15097__B _01955_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08952__A1 _03657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09722_ irq_mask\[9\] _04448_ timer\[9\] _04024_ _04027_ VGND VGND VPWR VPWR _04449_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__15317__S _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12530__A _06751_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16227__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09653_ _04100_ _04372_ _04381_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__or3_4
X_08604_ irq_mask\[1\] irq_active _03269_ _03272_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__o211a_1
XANTENNA__08977__B_N _03206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09584_ cpuregs.regs\[16\]\[6\] cpuregs.regs\[17\]\[6\] cpuregs.regs\[18\]\[6\] cpuregs.regs\[19\]\[6\]
+ _04217_ _04219_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08535_ _03312_ _03313_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__nand2_1
XANTENNA__12676__S _06825_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13361__A _04040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08466_ _03249_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__inv_2
XANTENNA__08455__A _03196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13213__A0 _06968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09417__C1 _04150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14961__A0 net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11775__A0 _06320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10122__S0 _04282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10673__S1 _05237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14192__A latched_branch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15061__S0 _03670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13300__S _07176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09286__A instr_timer VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09018_ _03728_ _03764_ _03765_ _03766_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_20_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10290_ cpuregs.regs\[4\]\[25\] cpuregs.regs\[5\]\[25\] cpuregs.regs\[6\]\[25\] cpuregs.regs\[7\]\[25\]
+ _04291_ _04292_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09196__B2 _03885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16611__S _03040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15269__A1 decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13980_ _07737_ _07752_ VGND VGND VPWR VPWR _07753_ sky130_fd_sc_hd__and2_1
XANTENNA__10189__S0 _04084_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12931_ _06974_ cpuregs.regs\[31\]\[15\] _06964_ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__mux2_1
XANTENNA__15784__B_N is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10502__A1 _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10502__B2 _05206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15650_ cpu_state\[0\] _02474_ _02472_ mem_do_wdata VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__a2bb2o_1
X_12862_ _06274_ cpuregs.regs\[6\]\[22\] _06928_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _06114_ cpuregs.regs\[11\]\[3\] _06348_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__mux2_1
X_14601_ _08241_ _08243_ _08239_ VGND VGND VPWR VPWR _08255_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_103_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ decoded_imm\[28\] _02216_ _02197_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ cpuregs.regs\[9\]\[22\] _06580_ _06891_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17320_ clknet_leaf_132_clk _00494_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14532_ _07946_ _08185_ VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__nor2_1
X_11744_ _06291_ _06292_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17251_ clknet_leaf_132_clk _00425_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14463_ decoded_imm_j\[13\] _07934_ VGND VGND VPWR VPWR _08128_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11675_ _06231_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__buf_2
XFILLER_0_153_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16582__A _03003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10018__B1 net300 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13414_ _07276_ VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__buf_2
XANTENNA__09959__B1 decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16202_ _03849_ _02821_ _02822_ _01821_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10626_ _05281_ _05285_ _05303_ _05328_ VGND VGND VPWR VPWR alu_out\[1\] sky130_fd_sc_hd__a211o_1
X_17182_ clknet_leaf_167_clk _00356_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14394_ _03368_ _08064_ VGND VGND VPWR VPWR _08065_ sky130_fd_sc_hd__nand2_1
XANTENNA__11766__A0 _06312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16133_ net291 net127 _02771_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13345_ _03387_ _07208_ _07211_ reg_next_pc\[0\] VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_3_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10557_ _05260_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_118_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08812__B net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16064_ _03403_ _02610_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13276_ _07153_ VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__buf_6
X_10488_ cpuregs.regs\[0\]\[31\] cpuregs.regs\[1\]\[31\] cpuregs.regs\[2\]\[31\] cpuregs.regs\[3\]\[31\]
+ _04325_ _04277_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__mux4_1
X_15015_ irq_mask\[17\] _01880_ _01889_ _01876_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12227_ cpuregs.regs\[24\]\[24\] _06584_ _06576_ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__mux2_1
XANTENNA__10416__S1 _04284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16521__S _02990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12158_ _06104_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__buf_2
XANTENNA__15355__S1 _01971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11109_ _03445_ _05770_ _03594_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__a21o_1
XANTENNA__08781__A_N net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16966_ clknet_leaf_138_clk _00140_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_12089_ _06114_ cpuregs.regs\[23\]\[3\] _06496_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15917_ instr_add _02617_ _02614_ _02653_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__a22o_1
XANTENNA__13691__A0 _04913_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16897_ clknet_leaf_30_clk _00042_ VGND VGND VPWR VPWR mem_rdata_q\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15661__A _03301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18636_ clknet_leaf_131_clk _01696_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_15848_ _05969_ _03810_ _03864_ _02608_ _05973_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__a41o_1
XFILLER_0_59_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18567_ clknet_leaf_154_clk _01632_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15779_ _03376_ _07899_ _03363_ _07905_ _06186_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17518_ clknet_leaf_137_clk _00687_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18498_ clknet_leaf_138_clk _01563_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10352__S0 _04207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17449_ clknet_leaf_184_clk _00618_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10009__B1 _04082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15291__S0 _01982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15600__S _01907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14943__A0 net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09414__A2 _04014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13120__S _07082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput210 net210 VGND VGND VPWR VPWR mem_la_addr[26] sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput221 net221 VGND VGND VPWR VPWR mem_la_addr[7] sky130_fd_sc_hd__clkbuf_1
XANTENNA__11509__B1 _03293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput232 net232 VGND VGND VPWR VPWR mem_la_wdata[16] sky130_fd_sc_hd__buf_1
XFILLER_0_64_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput243 net243 VGND VGND VPWR VPWR mem_la_wdata[26] sky130_fd_sc_hd__buf_1
XFILLER_0_101_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput254 net254 VGND VGND VPWR VPWR mem_la_wdata[7] sky130_fd_sc_hd__buf_1
XFILLER_0_11_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput265 net265 VGND VGND VPWR VPWR mem_wdata[11] sky130_fd_sc_hd__buf_1
Xoutput276 net276 VGND VGND VPWR VPWR mem_wdata[21] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput287 net287 VGND VGND VPWR VPWR mem_wdata[31] sky130_fd_sc_hd__clkbuf_1
Xoutput298 net298 VGND VGND VPWR VPWR mem_wstrb[3] sky130_fd_sc_hd__clkbuf_1
XANTENNA__15671__A1 _02484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09705_ _04430_ _04431_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__or2_1
XANTENNA__09045__S _03730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_94_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09636_ cpuregs.regs\[0\]\[7\] cpuregs.regs\[1\]\[7\] cpuregs.regs\[2\]\[7\] cpuregs.regs\[3\]\[7\]
+ _04274_ _04317_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__mux4_1
XFILLER_0_168_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14226__A2 _07906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10591__S0 _05264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09567_ _04272_ _04288_ _04297_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08504__A_N _03196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08518_ _03298_ _03276_ _03289_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_65_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09498_ _04228_ _04229_ _04211_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08449_ mem_state\[0\] mem_state\[1\] VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__or2_1
XANTENNA__15187__B1 _02039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11460__A2 irq_pending\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14934__A0 net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11460_ _06041_ irq_pending\[18\] _06048_ net10 VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10411_ reg_pc\[28\] decoded_imm\[28\] _05115_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__nand3_1
XFILLER_0_116_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11391_ _03977_ _06000_ _03965_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__or3b_1
XFILLER_0_104_721 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13030__S _07032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13130_ _06953_ cpuregs.regs\[4\]\[5\] _07082_ VGND VGND VPWR VPWR _07088_ sky130_fd_sc_hd__mux2_1
X_10342_ _05049_ _05050_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10971__A1 _05255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13061_ _07051_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__clkbuf_1
X_10273_ _04954_ _04957_ _04955_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__o21ai_2
XANTENNA__16341__S _02896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_305 VGND VGND VPWR VPWR alphacore_305/HI cpi_insn[3] sky130_fd_sc_hd__conb_1
Xalphacore_316 VGND VGND VPWR VPWR alphacore_316/HI cpi_insn[14] sky130_fd_sc_hd__conb_1
X_12012_ _06458_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08916__A1 _03677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_327 VGND VGND VPWR VPWR alphacore_327/HI cpi_insn[25] sky130_fd_sc_hd__conb_1
XANTENNA__09744__A _04469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_338 VGND VGND VPWR VPWR alphacore_338/HI mem_la_addr[1] sky130_fd_sc_hd__conb_1
Xalphacore_349 VGND VGND VPWR VPWR alphacore_349/HI trace_data[10] sky130_fd_sc_hd__conb_1
XANTENNA__11920__A0 _06257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16820_ _03153_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12170__A _06140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16751_ _06531_ cpuregs.regs\[13\]\[0\] _03116_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__mux2_1
X_13963_ _07741_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_85_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_2
X_15702_ timer\[11\] timer\[10\] _02508_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_85_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12914_ _06174_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__buf_2
X_13894_ _07693_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__clkbuf_1
X_16682_ _03079_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14217__A2 _07906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_927 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18421_ clknet_leaf_15_clk _01486_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13713__B decoded_imm\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15633_ _02460_ mem_do_prefetch _03380_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__mux2_1
X_12845_ _06208_ cpuregs.regs\[6\]\[14\] _06917_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output204_A net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14097__A _06053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18352_ clknet_leaf_40_clk _01420_ VGND VGND VPWR VPWR mem_la_firstword_reg sky130_fd_sc_hd__dfxtp_1
XANTENNA__13976__B2 net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12776_ cpuregs.regs\[9\]\[14\] _06563_ _06880_ VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15564_ _01969_ _02388_ _02396_ _02027_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__o211a_2
XFILLER_0_83_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17303_ clknet_leaf_162_clk _00477_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_11727_ reg_out\[23\] alu_out_q\[23\] _06068_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__mux2_1
XANTENNA__11233__B _05868_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14515_ _08148_ _08165_ _08173_ _08175_ VGND VGND VPWR VPWR _08176_ sky130_fd_sc_hd__o211a_1
X_15495_ net114 _02331_ _03272_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18283_ clknet_leaf_32_clk _01351_ VGND VGND VPWR VPWR is_alu_reg_imm sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_155_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15273__S0 _01976_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17234_ clknet_leaf_114_clk _00408_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_172_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11658_ _06216_ cpuregs.regs\[10\]\[15\] _06176_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__mux2_1
X_14446_ _07899_ _07930_ _08050_ _08112_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__a31o_1
XFILLER_0_154_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10609_ _05013_ net85 _05263_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10564__S _05264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17165_ clknet_leaf_123_clk _00339_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_14377_ _08048_ VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__inv_2
X_11589_ _06071_ reg_next_pc\[8\] _06154_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08542__B irq_pending\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16116_ _02686_ _02774_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13328_ _04272_ _07194_ VGND VGND VPWR VPWR _07195_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_133_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17096_ clknet_leaf_142_clk _00270_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09028__B_N _03213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15656__A _07208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13259_ _07156_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__clkbuf_1
X_16047_ mem_rdata_q\[31\] _02726_ _02633_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__a21o_2
XANTENNA__14560__A _07998_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08969__S _03730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09654__A _04051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09580__A1 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17998_ clknet_leaf_103_clk _01135_ VGND VGND VPWR VPWR irq_mask\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16850__A0 _06565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16949_ clknet_leaf_53_clk _00077_ VGND VGND VPWR VPWR cpu_state\[3\] sky130_fd_sc_hd__dfxtp_4
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09421_ _04045_ _04154_ _04113_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18619_ clknet_leaf_16_clk _00093_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__dfxtp_4
XANTENNA__13623__B decoded_imm\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08717__B net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09352_ _04086_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__buf_6
XANTENNA__11978__A0 _06216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_150_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11442__A2 irq_pending\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09283_ count_instr\[0\] _04012_ count_cycle\[0\] _04014_ _04019_ VGND VGND VPWR
+ VPWR _04020_ sky130_fd_sc_hd__a221o_1
XFILLER_0_142_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16426__S _02943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13719__A1 _07217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15264__S0 _02022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14454__B _07986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_983 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_165_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15567__S1 _01980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10953__B2 _05281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08998_ mem_rdata_q\[11\] net35 _03208_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11318__B _05929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_67_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_170_Right_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10960_ _05644_ _05589_ _05331_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__mux2_1
XANTENNA__11130__A1 _05174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09619_ _04347_ _04348_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10891_ _05414_ _05579_ _05580_ _05298_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__o211a_1
XANTENNA__15947__A2 _02650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11334__A reg_next_pc\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12630_ _06216_ cpuregs.regs\[30\]\[15\] _06799_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10316__S0 _04123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12561_ _06768_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12864__S _06928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15255__S0 _02022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14300_ _07973_ _07974_ _07975_ _07976_ VGND VGND VPWR VPWR _07977_ sky130_fd_sc_hd__or4_1
XANTENNA__14907__A0 net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11512_ _06085_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__buf_6
XFILLER_0_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15280_ cpuregs.regs\[28\]\[11\] cpuregs.regs\[29\]\[11\] cpuregs.regs\[30\]\[11\]
+ cpuregs.regs\[31\]\[11\] _01999_ _02000_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12492_ _06731_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14231_ _05856_ _06180_ VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__or2_1
X_11443_ irq_mask\[11\] _06030_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10384__S _04369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11197__A1 _05829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14162_ count_instr\[54\] _07876_ _07877_ VGND VGND VPWR VPWR _07880_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_150_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11374_ cpuregs.raddr2\[3\] _05983_ _05984_ _05985_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_78_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15558__S1 _02070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13113_ _07078_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10325_ _04068_ _05034_ _00073_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__a21o_1
X_14093_ count_instr\[34\] count_instr\[33\] count_instr\[32\] _07824_ VGND VGND VPWR
+ VPWR _07831_ sky130_fd_sc_hd__and4_2
XANTENNA__14380__A decoded_imm_j\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15907__C mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17921_ clknet_leaf_54_clk _08380_ VGND VGND VPWR VPWR reg_out\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09474__A _04053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13044_ cpuregs.regs\[3\]\[29\] _06594_ _07032_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10256_ cpuregs.regs\[0\]\[24\] cpuregs.regs\[1\]\[24\] cpuregs.regs\[2\]\[24\] cpuregs.regs\[3\]\[24\]
+ _04290_ _04276_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__mux4_1
XANTENNA__10157__C1 _04027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output154_A net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12104__S _06507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17852_ clknet_leaf_104_clk _01021_ VGND VGND VPWR VPWR reg_next_pc\[29\] sky130_fd_sc_hd__dfxtp_1
X_10187_ cpuregs.regs\[4\]\[22\] cpuregs.regs\[5\]\[22\] cpuregs.regs\[6\]\[22\] cpuregs.regs\[7\]\[22\]
+ _04280_ _04059_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__mux4_1
X_16803_ _06586_ cpuregs.regs\[13\]\[25\] _03138_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__mux2_1
XANTENNA__11228__B _05864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12449__A1 _06590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17783_ clknet_leaf_85_clk _00952_ VGND VGND VPWR VPWR count_instr\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14995_ irq_mask\[9\] _01863_ _01714_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_58_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__09314__A1 _03226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
X_16734_ _03106_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__clkbuf_1
X_13946_ _07714_ _07729_ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__and2_1
XANTENNA__08818__A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_858 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16665_ cpuregs.regs\[1\]\[27\] _06311_ _03062_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__mux2_1
X_13877_ _07676_ _07679_ _07680_ VGND VGND VPWR VPWR _07681_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_157_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18404_ clknet_leaf_143_clk _01469_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15616_ _03719_ _02444_ _00068_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__o21a_1
X_12828_ _06141_ cpuregs.regs\[6\]\[6\] _06906_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__mux2_1
X_16596_ _03033_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18335_ clknet_leaf_35_clk _01403_ VGND VGND VPWR VPWR mem_16bit_buffer\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12774__S _06880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15547_ _03639_ _02376_ _02380_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__a21o_1
X_12759_ cpuregs.regs\[9\]\[6\] _06546_ _06869_ VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10632__B1 _05205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18266_ clknet_leaf_26_clk _01337_ VGND VGND VPWR VPWR decoded_imm\[24\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_115_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15478_ cpuregs.regs\[0\]\[23\] cpuregs.regs\[1\]\[23\] cpuregs.regs\[2\]\[23\] cpuregs.regs\[3\]\[23\]
+ _01995_ _01937_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17217_ clknet_leaf_189_clk _00391_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14374__A1 _07899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14429_ instr_jal _07754_ VGND VGND VPWR VPWR _08097_ sky130_fd_sc_hd__nand2_2
X_18197_ clknet_leaf_41_clk _01268_ VGND VGND VPWR VPWR instr_addi sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17148_ clknet_leaf_12_clk _00322_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10307__B decoded_imm\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09970_ cpuregs.regs\[20\]\[16\] cpuregs.regs\[21\]\[16\] cpuregs.regs\[22\]\[16\]
+ cpuregs.regs\[23\]\[16\] _04477_ _04478_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__mux4_1
X_17079_ clknet_leaf_177_clk _00253_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08921_ cpuregs.regs\[8\]\[3\] cpuregs.regs\[9\]\[3\] cpuregs.regs\[10\]\[3\] cpuregs.regs\[11\]\[3\]
+ _03641_ _03684_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08852_ net105 net73 VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__nand2_1
X_08783_ _03517_ _03518_ _03548_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_93_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09305__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11853__S _06370_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16010__A _02611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08728__A net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09400__S1 _04124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13353__B _03274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15929__A2 _02617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16051__A1 decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09404_ cpuregs.regs\[12\]\[2\] cpuregs.regs\[13\]\[2\] cpuregs.regs\[14\]\[2\] cpuregs.regs\[15\]\[2\]
+ _04123_ _04124_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09608__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09335_ _04069_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__buf_4
XFILLER_0_118_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12684__S _06825_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09559__A _04055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09266_ _03892_ _04002_ _03960_ _04003_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_747 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08463__A mem_do_wdata VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09197_ _03840_ _03941_ _03944_ _03751_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__a22o_1
XFILLER_0_172_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11179__A1 net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15314__B1 _03639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09792__A1 _04272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10110_ cpuregs.regs\[12\]\[20\] cpuregs.regs\[13\]\[20\] cpuregs.regs\[14\]\[20\]
+ cpuregs.regs\[15\]\[20\] _04275_ _04278_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11090_ _03441_ _05398_ _05367_ _03440_ _05646_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_101_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10041_ _04233_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_73_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13628__A0 _04810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13544__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13800_ _03631_ _07635_ _07636_ VGND VGND VPWR VPWR _07637_ sky130_fd_sc_hd__nor3_1
X_14780_ count_cycle\[28\] count_cycle\[29\] _01736_ _03240_ VGND VGND VPWR VPWR _01740_
+ sky130_fd_sc_hd__a31o_1
X_11992_ _06448_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10537__S0 _05230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10943_ _03485_ _03488_ _05608_ _05628_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__a31o_1
X_13731_ _05143_ _07277_ _07532_ _07217_ VGND VGND VPWR VPWR _07573_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11064__A _05225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16042__B2 mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16450_ _02956_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__clkbuf_1
X_13662_ _03276_ _07508_ VGND VGND VPWR VPWR _07509_ sky130_fd_sc_hd__and2_1
X_10874_ _05557_ _05558_ _05560_ _05564_ _05250_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__o32a_1
XFILLER_0_39_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14053__B1 _07790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15401_ cpuregs.regs\[8\]\[18\] cpuregs.regs\[9\]\[18\] cpuregs.regs\[10\]\[18\]
+ cpuregs.regs\[11\]\[18\] _03645_ _01991_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12613_ _06150_ cpuregs.regs\[30\]\[7\] _06788_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13593_ _07444_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__clkbuf_1
X_16381_ _06987_ cpuregs.regs\[16\]\[21\] _02918_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18120_ clknet_leaf_54_clk _01224_ VGND VGND VPWR VPWR latched_stalu sky130_fd_sc_hd__dfxtp_2
XFILLER_0_171_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15332_ cpuregs.regs\[24\]\[14\] cpuregs.regs\[25\]\[14\] cpuregs.regs\[26\]\[14\]
+ cpuregs.regs\[27\]\[14\] _02074_ _02075_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__mux4_1
X_12544_ _06759_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08902__S0 _03658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18051_ clknet_leaf_45_clk _01156_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dfxtp_2
XANTENNA__10090__B2 _04023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12475_ _06722_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__clkbuf_1
X_15263_ _02111_ _02112_ _02017_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17002_ clknet_leaf_139_clk _00176_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_11426_ _03412_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_113_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14214_ reg_pc\[5\] _07906_ _07917_ _07912_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__a22o_1
X_15194_ _03646_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_6 _02000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15918__B mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14145_ count_instr\[49\] _07865_ _07867_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11938__S _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11357_ _05971_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15400__S0 _03649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10308_ _05016_ _05017_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__nand2_1
XANTENNA_output79_A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14076_ _07818_ _07819_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__nor2_1
X_11288_ _03841_ _05912_ _05913_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_167_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17904_ clknet_leaf_87_clk _01073_ VGND VGND VPWR VPWR count_cycle\[49\] sky130_fd_sc_hd__dfxtp_1
X_13027_ _07033_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__clkbuf_1
X_10239_ _04875_ _04950_ _04919_ _04886_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__a211o_1
XANTENNA__15934__A mem_rdata_q\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10143__A _04272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16805__A0 _06588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17835_ clknet_leaf_57_clk _01004_ VGND VGND VPWR VPWR reg_next_pc\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13454__A _05257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17766_ clknet_leaf_94_clk _00935_ VGND VGND VPWR VPWR count_instr\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14978_ _04142_ _01865_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16717_ _03097_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09394__S0 _04071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13929_ _07714_ _07717_ VGND VGND VPWR VPWR _07718_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17697_ clknet_leaf_75_clk _00866_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16033__A1 mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15467__S0 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16648_ cpuregs.regs\[1\]\[19\] _06247_ _03051_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14595__A1 _03379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16579_ _03024_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10605__A0 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15219__S0 _02069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09120_ _03798_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__clkbuf_4
X_18318_ clknet_leaf_38_clk _01386_ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09471__B1 _04008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14347__A1 _07988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09051_ _03811_ _03812_ _03231_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18249_ clknet_leaf_23_clk _01320_ VGND VGND VPWR VPWR decoded_imm\[7\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__14347__B2 _08012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16704__S _03087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10369__C1 _04202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14732__B _08350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09774__A1 _03638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09774__B2 _03226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09953_ _04667_ _04670_ _04673_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_55_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08904_ _00064_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__clkbuf_8
X_09884_ irq_pending\[13\] _04008_ _04596_ _04606_ VGND VGND VPWR VPWR _08373_ sky130_fd_sc_hd__o22a_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09842__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08835_ is_slti_blt_slt _03431_ _03600_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__and3_1
X_08766_ net121 net89 VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__or2_2
XFILLER_0_169_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08458__A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11097__B1 _05517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08697_ _03461_ _03462_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__and2_1
XANTENNA__10439__A3 _05145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16024__B2 mem_rdata_q\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14195__A _03298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09318_ _04052_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_97_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10590_ _04039_ _04198_ _04160_ _04251_ _05239_ _05237_ VGND VGND VPWR VPWR _05293_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09462__B1 _04156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11331__B _05948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09249_ _03902_ _03885_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15535__B1 _00068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14338__B2 reg_next_pc\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10228__A _04940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12260_ _06607_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_999 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09214__B1 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14642__B _07988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11211_ _05850_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_75_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09765__A1 _04053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09736__B decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12191_ _06560_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15299__C1 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11142_ _03407_ _05413_ net100 _04422_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__a22o_2
XANTENNA__09860__S1 _04469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput76 net76 VGND VGND VPWR VPWR cpi_rs1[18] sky130_fd_sc_hd__buf_1
Xoutput87 net87 VGND VGND VPWR VPWR cpi_rs1[28] sky130_fd_sc_hd__clkbuf_1
XANTENNA__15754__A _02476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14510__A1 reg_next_pc\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11073_ _03449_ _05357_ _05749_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__o21ai_1
X_15950_ _03305_ mem_rdata_q\[2\] _02671_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__and3_1
XANTENNA__14510__B2 _07960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput98 net98 VGND VGND VPWR VPWR cpi_rs1[9] sky130_fd_sc_hd__buf_1
XANTENNA__10127__A2 _04448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10024_ count_cycle\[17\] _04014_ _04742_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__a21o_1
X_14901_ net214 net183 _01824_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__mux2_1
XANTENNA__09752__A _04086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12589__S _06774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15881_ _02633_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10898__A _05292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_920 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17620_ clknet_leaf_152_clk _00789_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_14832_ _01774_ _01775_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14274__B1 _07942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11088__A0 _05086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17551_ clknet_leaf_145_clk _00720_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_14763_ _01728_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11975_ _06439_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output117_A net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09898__S _04222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16502_ cpuregs.regs\[17\]\[14\] _06563_ _02979_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__mux2_1
XANTENNA__15449__S0 _02085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13714_ _07555_ _07556_ VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10926_ _03483_ _05608_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_123_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17482_ clknet_leaf_175_clk _00651_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14694_ count_cycle\[0\] count_cycle\[1\] count_cycle\[2\] VGND VGND VPWR VPWR _08338_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10930__S0 _05237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16433_ _02947_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14577__A1 _08232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10857_ _05361_ _05536_ _05537_ _05548_ VGND VGND VPWR VPWR alu_out\[12\] sky130_fd_sc_hd__a31o_2
X_13645_ _03631_ _07492_ _07271_ VGND VGND VPWR VPWR _07493_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13213__S _07129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09679__S1 _04087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16364_ _06970_ cpuregs.regs\[16\]\[13\] _02907_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10788_ net98 _03510_ _03518_ net95 _05236_ _05309_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__mux4_1
X_13576_ reg_pc\[14\] _07211_ _07428_ _07221_ VGND VGND VPWR VPWR _07429_ sky130_fd_sc_hd__a211o_1
XFILLER_0_143_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18103_ clknet_leaf_80_clk _01207_ VGND VGND VPWR VPWR timer\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15315_ cpuregs.regs\[4\]\[13\] cpuregs.regs\[5\]\[13\] cpuregs.regs\[6\]\[13\] cpuregs.regs\[7\]\[13\]
+ _02022_ _02023_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__mux4_1
XFILLER_0_147_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12527_ _06749_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__clkbuf_1
X_16295_ _06970_ cpuregs.regs\[15\]\[13\] _02870_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18034_ clknet_leaf_66_clk _00010_ VGND VGND VPWR VPWR irq_pending\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13537__C1 _07221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15621__S0 _03645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15246_ _02091_ _02093_ _02096_ _02088_ _02018_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_10_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12458_ _06712_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_169_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09756__A1 _04070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13449__A net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11409_ _05969_ _03913_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15177_ _03684_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__buf_6
X_12389_ _06675_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08550__B _03326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15829__A1 decoded_imm_j\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09851__S1 _04513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14128_ _07778_ _07854_ _07855_ VGND VGND VPWR VPWR _07856_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15664__A _02484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14059_ count_instr\[23\] _07805_ _07807_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__o21a_1
XANTENNA__11315__A1 _05044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10749__S0 _05277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12499__S _06726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10669__A3 _04611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08620_ _03304_ _03393_ _03394_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__a21oi_1
X_17818_ clknet_leaf_66_clk _00987_ VGND VGND VPWR VPWR reg_pc\[26\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_118_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08551_ irq_mask\[16\] irq_pending\[16\] VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__and2b_2
X_17749_ clknet_leaf_86_clk _00918_ VGND VGND VPWR VPWR count_instr\[20\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11618__A2 _03335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15603__S _02110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08482_ instr_beq instr_waitirq instr_srai instr_slli VGND VGND VPWR VPWR _03266_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_147_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12528__A cpuregs.waddr\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08725__B net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09103_ _03770_ _03776_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16434__S _02943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12962__S _06985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14743__A _03239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09034_ mem_rdata_q\[6\] net61 _03227_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09936_ _04053_ _04656_ _04095_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_70_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _04584_ _04586_ _04589_ _04053_ _04095_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ net84 VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__inv_2
XANTENNA__12202__S _06555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09798_ _04521_ _04522_ _04321_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__mux2_1
XANTENNA__09358__S0 _04056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08749_ _03513_ _03514_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__nand2b_2
XANTENNA__16609__S _03040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11760_ reg_pc\[26\] reg_pc\[25\] _06283_ reg_pc\[27\] VGND VGND VPWR VPWR _06307_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _03544_ _05409_ _05390_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__mux2_1
XANTENNA__10293__A1 _04430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13541__B decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11691_ _03409_ _03358_ _06066_ _06245_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13767__C1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10642_ _05240_ _05342_ _05343_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__o21ai_1
X_13430_ _03631_ _07290_ _07292_ _07271_ VGND VGND VPWR VPWR _07293_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_101_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10045__A1 _04430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13361_ _04040_ decoded_imm\[1\] VGND VGND VPWR VPWR _07227_ sky130_fd_sc_hd__nand2_1
XANTENNA__15508__B1 _02017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10573_ _05243_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__buf_4
XANTENNA__09986__B2 _04014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12872__S _06928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10140__S1 _04285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15100_ _03396_ _03679_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09747__A _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12312_ _06634_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__clkbuf_1
X_13292_ _07173_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__clkbuf_1
X_16080_ decoded_imm\[30\] _02750_ _02745_ mem_rdata_q\[30\] _02748_ VGND VGND VPWR
+ VPWR _01343_ sky130_fd_sc_hd__a221o_1
XFILLER_0_161_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_125_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15031_ irq_mask\[25\] _01863_ _03240_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12243_ _06595_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10392__S _04222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12173__A _06149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09833__S1 _04073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12174_ cpuregs.regs\[24\]\[7\] _06548_ _06534_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11125_ _05517_ _05797_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__nand2_1
X_16982_ clknet_leaf_116_clk _00156_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09482__A _04068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11056_ _03452_ _05357_ _05733_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__o21ai_1
X_15933_ _02655_ _02658_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__and2_2
XANTENNA_output234_A net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10007_ cpuregs.regs\[24\]\[17\] cpuregs.regs\[25\]\[17\] cpuregs.regs\[26\]\[17\]
+ cpuregs.regs\[27\]\[17\] _04072_ _04074_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ instr_bne _02618_ _02620_ _02622_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_125_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12112__S _06507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10520__A2 _05220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17603_ clknet_leaf_7_clk _00772_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14815_ count_cycle\[40\] _01762_ _01717_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__a21oi_1
X_18583_ clknet_leaf_17_clk _01648_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08779__B_N _03524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15795_ _03292_ _03226_ _03282_ _03305_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__o211a_1
XANTENNA__16519__S _02990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11951__S _06424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17534_ clknet_leaf_125_clk _00703_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_14746_ count_cycle\[18\] _08368_ _01716_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__o21a_1
XFILLER_0_171_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11958_ _06430_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08826__A net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10909_ _05596_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17465_ clknet_leaf_160_clk _00634_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14677_ _08121_ _08323_ _08324_ VGND VGND VPWR VPWR _08325_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_15_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11889_ _06393_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08545__B _03321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16416_ _02938_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13628_ _04810_ _04744_ _07276_ VGND VGND VPWR VPWR _07477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17396_ clknet_leaf_179_clk _00565_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12782__S _06880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16347_ _06953_ cpuregs.regs\[16\]\[5\] _02896_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__mux2_1
X_13559_ _04456_ _05258_ _07412_ _07216_ VGND VGND VPWR VPWR _07413_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10587__A2 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16278_ _06953_ cpuregs.regs\[15\]\[5\] _02859_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__mux2_1
X_18017_ clknet_leaf_64_clk _00012_ VGND VGND VPWR VPWR irq_pending\[1\] sky130_fd_sc_hd__dfxtp_1
X_15229_ net129 _01906_ _02079_ _02080_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__o22a_1
XFILLER_0_140_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09376__B _04038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16475__A1 _06536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09392__A _00071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09721_ _04308_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09588__S0 _04274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09652_ _04206_ _04375_ _04380_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08603_ _03250_ _03380_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__nor2_1
X_09583_ cpuregs.regs\[20\]\[6\] cpuregs.regs\[21\]\[6\] cpuregs.regs\[22\]\[6\] cpuregs.regs\[23\]\[6\]
+ _04217_ _04219_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__mux4_1
XANTENNA__15333__S _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11861__S _06370_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08534_ reg_sh\[4\] reg_sh\[3\] reg_sh\[2\] VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__nor3_2
XFILLER_0_49_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09331__S _04065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11472__B1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15738__B1 _02488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13361__B decoded_imm\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08465_ _03246_ _03248_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__or2_2
XFILLER_0_159_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10027__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14961__A1 net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14473__A _06863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10122__S1 _04285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08640__A1 _03407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09017_ _03743_ _03748_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__nand2_2
XFILLER_0_103_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15061__S1 _03671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12724__A0 _06312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15269__A2 _02009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09919_ reg_pc\[14\] decoded_imm\[14\] _04608_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__a21o_1
XANTENNA__10189__S1 _04086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13028__S _07032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12930_ _06215_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10502__A2 _05205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12861_ _06930_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16339__S _02896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11771__S _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13552__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14600_ _08212_ _07959_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_103_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _06351_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15580_ _02020_ _02403_ _02411_ _02027_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__o211a_2
XANTENNA__09656__B1 instr_rdinstr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08646__A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12792_ _06893_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_120_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10266__A1 _04328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14531_ _08177_ _08180_ _08189_ VGND VGND VPWR VPWR _08191_ sky130_fd_sc_hd__nand3_1
X_11743_ reg_pc\[25\] _06283_ _06101_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_83_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17250_ clknet_leaf_183_clk _00424_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09408__B1 _04133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14462_ _08084_ _08086_ _08094_ _08124_ VGND VGND VPWR VPWR _08127_ sky130_fd_sc_hd__or4_1
X_11674_ _06226_ reg_next_pc\[17\] _06228_ _06230_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__a211o_4
XFILLER_0_36_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16201_ _02685_ _02821_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13413_ _05209_ VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__buf_2
XANTENNA__09503__S0 _04232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10625_ _05255_ _05261_ _05321_ _05327_ _05225_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__a32o_1
XFILLER_0_154_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17181_ clknet_leaf_2_clk _00355_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15479__A _03709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14393_ _08052_ _08058_ _08057_ _08062_ VGND VGND VPWR VPWR _08064_ sky130_fd_sc_hd__a31o_1
XANTENNA__14383__A _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11800__A _06342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16132_ _02783_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__clkbuf_1
X_13344_ _07210_ VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__clkbuf_4
X_10556_ _05259_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__buf_4
XFILLER_0_134_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output184_A net184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16063_ decoded_imm\[19\] _02611_ _02736_ _02744_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__o22a_1
X_13275_ _07164_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__clkbuf_1
X_10487_ cpuregs.regs\[4\]\[31\] cpuregs.regs\[5\]\[31\] cpuregs.regs\[6\]\[31\] cpuregs.regs\[7\]\[31\]
+ _04325_ _04277_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__mux4_1
X_15014_ _04737_ _01885_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12226_ _06288_ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__buf_2
XFILLER_0_121_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12157_ _06537_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14322__S _07998_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14468__B1 _08012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11108_ _05219_ _05774_ _05782_ VGND VGND VPWR VPWR alu_out\[29\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16965_ clknet_leaf_149_clk _00139_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_12088_ _06499_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_142_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16209__A1 _06081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11039_ _03455_ _05367_ _05222_ _03454_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__a2bb2o_1
X_15916_ _02652_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__buf_2
X_16896_ clknet_leaf_30_clk _00041_ VGND VGND VPWR VPWR mem_rdata_q\[15\] sky130_fd_sc_hd__dfxtp_1
X_18635_ clknet_leaf_129_clk _01695_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15661__B _04024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15847_ _03798_ _02607_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18566_ clknet_leaf_146_clk _01631_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_15778_ _05201_ _02486_ _02570_ _02545_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13982__A_N instr_waitirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17517_ clknet_leaf_148_clk _00686_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11454__B1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14729_ count_cycle\[13\] _08359_ _08361_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18497_ clknet_leaf_156_clk _01562_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10352__S1 _04208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17448_ clknet_leaf_175_clk _00617_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16393__A0 _06999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08990__S _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_151_Left_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11206__A0 _04342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10009__A1 _04231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14943__A1 net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15291__S1 _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17379_ clknet_leaf_14_clk _00548_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13401__S _05257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09387__A _04077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12017__S _06460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput200 net200 VGND VGND VPWR VPWR mem_la_addr[16] sky130_fd_sc_hd__buf_1
XANTENNA__11509__A1 latched_branch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16712__S _03087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput211 net211 VGND VGND VPWR VPWR mem_la_addr[27] sky130_fd_sc_hd__buf_1
XFILLER_0_101_917 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput222 net222 VGND VGND VPWR VPWR mem_la_addr[8] sky130_fd_sc_hd__clkbuf_1
Xoutput233 net233 VGND VGND VPWR VPWR mem_la_wdata[17] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput244 net244 VGND VGND VPWR VPWR mem_la_wdata[27] sky130_fd_sc_hd__buf_1
Xoutput255 net255 VGND VGND VPWR VPWR mem_la_wdata[8] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput266 net266 VGND VGND VPWR VPWR mem_wdata[12] sky130_fd_sc_hd__clkbuf_1
Xoutput277 net277 VGND VGND VPWR VPWR mem_wdata[22] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput288 net288 VGND VGND VPWR VPWR mem_wdata[3] sky130_fd_sc_hd__clkbuf_1
Xoutput299 net299 VGND VGND VPWR VPWR trap sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_160_Left_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09704_ cpuregs.regs\[0\]\[9\] cpuregs.regs\[1\]\[9\] cpuregs.regs\[2\]\[9\] cpuregs.regs\[3\]\[9\]
+ _04325_ _04277_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09635_ cpuregs.regs\[4\]\[7\] cpuregs.regs\[5\]\[7\] cpuregs.regs\[6\]\[7\] cpuregs.regs\[7\]\[7\]
+ _04274_ _04317_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__mux4_1
XFILLER_0_168_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10591__S1 _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09566_ _04289_ _04295_ _04296_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10248__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08517_ cpu_state\[1\] VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13985__A2 _07755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09497_ cpuregs.regs\[0\]\[4\] cpuregs.regs\[1\]\[4\] cpuregs.regs\[2\]\[4\] cpuregs.regs\[3\]\[4\]
+ _04207_ _04208_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__mux4_1
XANTENNA__15187__A1 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08448_ _03227_ _03228_ _03231_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10410_ _05084_ _05115_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09297__A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11390_ _03954_ _03987_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10341_ reg_pc\[27\] decoded_imm\[27\] VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14698__B1 _07877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10971__A2 _05394_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13060_ _06951_ cpuregs.regs\[7\]\[4\] _07046_ VGND VGND VPWR VPWR _07051_ sky130_fd_sc_hd__mux2_1
X_10272_ irq_pending\[24\] _04049_ _04958_ _03385_ _04983_ VGND VGND VPWR VPWR _08385_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xalphacore_306 VGND VGND VPWR VPWR alphacore_306/HI cpi_insn[4] sky130_fd_sc_hd__conb_1
X_12011_ _06343_ cpuregs.regs\[21\]\[31\] _06423_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__mux2_1
XANTENNA__11766__S _06258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xalphacore_317 VGND VGND VPWR VPWR alphacore_317/HI cpi_insn[15] sky130_fd_sc_hd__conb_1
XANTENNA__08916__A2 _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_328 VGND VGND VPWR VPWR alphacore_328/HI cpi_insn[26] sky130_fd_sc_hd__conb_1
Xalphacore_339 VGND VGND VPWR VPWR alphacore_339/HI trace_data[0] sky130_fd_sc_hd__conb_1
XFILLER_0_100_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15762__A _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16750_ _03115_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__buf_6
X_13962_ _07737_ _07740_ VGND VGND VPWR VPWR _07741_ sky130_fd_sc_hd__and2_1
X_15701_ _02477_ _02512_ _02513_ _02481_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__o211a_1
X_12913_ _06962_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16681_ _06947_ cpuregs.regs\[19\]\[2\] _03076_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__mux2_1
X_13893_ _07691_ _07692_ VGND VGND VPWR VPWR _07693_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16611__A1 _06095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18420_ clknet_leaf_176_clk _01485_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_15632_ _04271_ instr_jalr VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12844_ _06921_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14622__B1 _07997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11436__B1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18351_ clknet_leaf_36_clk _01419_ VGND VGND VPWR VPWR mem_rdata_q\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13976__A2 _07677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15563_ _02390_ _02392_ _02395_ _02004_ _02088_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__a221o_1
X_12775_ _06884_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17302_ clknet_leaf_128_clk _00476_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_14514_ decoded_imm_j\[16\] _07941_ _08131_ _08174_ VGND VGND VPWR VPWR _08175_ sky130_fd_sc_hd__a22oi_1
X_11726_ reg_pc\[23\] _06268_ _06276_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__o21a_1
X_18282_ clknet_leaf_24_clk _01350_ VGND VGND VPWR VPWR is_beq_bne_blt_bge_bltu_bgeu
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15494_ _01959_ _02322_ _02330_ _01933_ decoded_imm\[23\] VGND VGND VPWR VPWR _02331_
+ sky130_fd_sc_hd__a32o_4
XTAP_TAPCELL_ROW_155_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15273__S1 _01977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17233_ clknet_leaf_160_clk _00407_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14445_ reg_next_pc\[11\] _07947_ _08111_ _08033_ VGND VGND VPWR VPWR _08112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11657_ _06215_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_172_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13221__S _07129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16127__A0 net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10608_ _05306_ _05310_ _05246_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__mux2_1
XANTENNA__08604__A1 irq_mask\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17164_ clknet_leaf_149_clk _00338_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14376_ _07919_ _08036_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11588_ irq_state\[1\] _03359_ _06065_ _06153_ _06074_ VGND VGND VPWR VPWR _06154_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16115_ _02681_ _02682_ _02773_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13327_ _07192_ _07193_ _04287_ VGND VGND VPWR VPWR _07194_ sky130_fd_sc_hd__mux2_1
X_10539_ _05242_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__clkbuf_4
X_17095_ clknet_leaf_147_clk _00269_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10962__A2 _05398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16046_ decoded_imm\[11\] _02720_ _02734_ _02735_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__o22a_1
X_13258_ _06945_ cpuregs.regs\[5\]\[1\] _07154_ VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15656__B _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15350__B2 _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11676__S _06176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15148__S _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13457__A _04262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12209_ _06572_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09654__B _04382_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10175__B1 _04017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13189_ _07119_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__clkbuf_1
X_17997_ clknet_leaf_103_clk _01134_ VGND VGND VPWR VPWR irq_mask\[13\] sky130_fd_sc_hd__dfxtp_1
X_16948_ clknet_leaf_53_clk _00076_ VGND VGND VPWR VPWR cpu_state\[2\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__13664__A1 _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10478__B2 _04165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16879_ _06594_ cpuregs.regs\[14\]\[29\] _03174_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__mux2_1
XANTENNA__08540__B1 instr_waitirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09420_ reg_pc\[1\] decoded_imm\[1\] VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__nor2_1
X_18618_ clknet_leaf_9_clk _00092_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09715__S0 _04072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09351_ _00070_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__buf_6
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18549_ clknet_leaf_14_clk _01614_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09282_ count_instr\[32\] _04016_ _04018_ count_cycle\[32\] VGND VGND VPWR VPWR _04019_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15264__S1 _02023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10755__S _05390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10402__A1 _04009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16669__A1 _06327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16442__S _02943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15892__A2 _02635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10705__A2 _05221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08997_ mem_rdata_q\[27\] net52 _03208_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__mux2_1
XANTENNA__11318__C _05932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10469__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10013__S0 _04280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14198__A _07905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11130__A2 _05143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13306__S _07176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09618_ reg_pc\[6\] decoded_imm\[6\] VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10890_ _05414_ _05436_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09706__S0 _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09549_ _04055_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__buf_6
XANTENNA__09087__A1 _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16617__S _03040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10316__S1 _04124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12560_ cpuregs.regs\[2\]\[14\] _06563_ _06763_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14645__B _07967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15255__S1 _02023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11511_ _06080_ _06084_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__nand2_2
X_12491_ _06208_ cpuregs.regs\[28\]\[14\] _06726_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__mux2_1
XANTENNA__08643__B _03274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ reg_pc\[10\] _07926_ _07928_ _07912_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__a22o_1
X_11442_ _06029_ irq_pending\[10\] _06038_ net2 VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__a31o_1
XANTENNA__15580__A1 _02020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14161_ count_instr\[54\] count_instr\[53\] _07874_ VGND VGND VPWR VPWR _07879_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11373_ _05969_ _03634_ _03889_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_150_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13112_ _07003_ cpuregs.regs\[7\]\[29\] _07068_ VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__mux2_1
X_10324_ _05032_ _05033_ _04063_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__mux2_1
X_14092_ _07830_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11496__S _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15907__D mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17920_ clknet_leaf_64_clk _08369_ VGND VGND VPWR VPWR reg_out\[0\] sky130_fd_sc_hd__dfxtp_1
X_10255_ cpuregs.regs\[4\]\[24\] cpuregs.regs\[5\]\[24\] cpuregs.regs\[6\]\[24\] cpuregs.regs\[7\]\[24\]
+ _04290_ _04276_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__mux4_1
X_13043_ _07041_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10252__S0 _04216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17851_ clknet_leaf_104_clk _01020_ VGND VGND VPWR VPWR reg_next_pc\[28\] sky130_fd_sc_hd__dfxtp_1
X_10186_ _04369_ _04899_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__or2_1
X_16802_ _03143_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__clkbuf_1
X_17782_ clknet_leaf_85_clk _00951_ VGND VGND VPWR VPWR count_instr\[53\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15191__S0 _01936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13646__A1 _04810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14994_ irq_mask\[8\] _01864_ _01877_ _01876_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__a211o_1
XANTENNA__09490__A _04063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09314__A2 _04043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16733_ _06999_ cpuregs.regs\[19\]\[27\] _03098_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__mux2_1
X_13945_ _03332_ _07727_ _07728_ net143 VGND VGND VPWR VPWR _07729_ sky130_fd_sc_hd__a22o_1
XANTENNA__12120__S _06507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16664_ _03069_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__clkbuf_1
X_13876_ _03271_ instr_retirq VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__nor2_1
XANTENNA__15399__B2 _02017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18403_ clknet_leaf_147_clk _01468_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_15615_ cpuregs.regs\[20\]\[31\] cpuregs.regs\[21\]\[31\] cpuregs.regs\[22\]\[31\]
+ cpuregs.regs\[23\]\[31\] _01995_ _01937_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__mux4_1
XANTENNA__16060__A2 decoded_imm_j\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11244__B _05877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12827_ _06912_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__clkbuf_1
X_16595_ _06997_ cpuregs.regs\[18\]\[26\] _03026_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__mux2_1
XANTENNA__16527__S _02990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18334_ clknet_leaf_36_clk _01402_ VGND VGND VPWR VPWR mem_16bit_buffer\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15546_ _03675_ _02379_ _03657_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__a21o_1
X_12758_ _06875_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14555__B _07952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11709_ _06260_ _06118_ _06261_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__and3b_1
XFILLER_0_38_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18265_ clknet_leaf_25_clk _01336_ VGND VGND VPWR VPWR decoded_imm\[23\] sky130_fd_sc_hd__dfxtp_4
X_15477_ net113 _01905_ _02313_ _02314_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_135_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12689_ _06175_ cpuregs.regs\[12\]\[10\] _06836_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__mux2_1
XANTENNA__08553__B irq_pending\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17216_ clknet_leaf_174_clk _00390_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_14428_ _08082_ _08094_ VGND VGND VPWR VPWR _08096_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18196_ clknet_leaf_29_clk _01267_ VGND VGND VPWR VPWR instr_sh sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17147_ clknet_leaf_12_clk _00321_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14359_ _03378_ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10396__B1 _00073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09665__A reg_pc\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10491__S0 _04329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17078_ clknet_leaf_127_clk _00252_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08920_ _03662_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__buf_6
X_16029_ _02712_ _02716_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13885__A1 _03326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11896__A0 _06166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08851_ net105 net73 VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15606__S _02110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08782_ _03517_ _03518_ _03522_ _03546_ _03547_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__a221o_1
XANTENNA__13637__A1 _07274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08728__B net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16036__C1 _02634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13126__S _07082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09403_ _04064_ _04136_ _04068_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12965__S _06985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12073__A0 _06320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09334_ _04068_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__buf_6
XFILLER_0_164_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10485__S _04321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09265_ _03942_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08463__B _03218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09196_ _03853_ _03942_ _03943_ _03869_ _03885_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__a32o_1
XFILLER_0_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11179__A2 _04710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12376__A1 _06586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09241__A1 _03878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15314__A1 _01989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10139__B1 _04014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12205__S _06555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10040_ _04232_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_73_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13628__A1 _04744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08919__A _03654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09927__S0 _04085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13544__B decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11991_ _06266_ cpuregs.regs\[21\]\[21\] _06446_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__mux2_1
XANTENNA__11103__A2 _05215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11345__A _03228_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13036__S _07032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13730_ _03275_ _07570_ _07571_ VGND VGND VPWR VPWR _07572_ sky130_fd_sc_hd__and3_1
XANTENNA__16578__A0 _06980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10942_ net106 net74 _05620_ _03487_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13661_ _07488_ _07502_ _07504_ _07505_ _07501_ VGND VGND VPWR VPWR _07508_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_27_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10873_ _05287_ _05418_ _05563_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__o21a_1
XANTENNA__16347__S _02896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15400_ cpuregs.regs\[12\]\[18\] cpuregs.regs\[13\]\[18\] cpuregs.regs\[14\]\[18\]
+ cpuregs.regs\[15\]\[18\] _03649_ _03643_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__mux4_1
X_12612_ _06795_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16380_ _02919_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__clkbuf_1
X_13592_ _04642_ _07443_ _07374_ VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15331_ cpuregs.regs\[28\]\[14\] cpuregs.regs\[29\]\[14\] cpuregs.regs\[30\]\[14\]
+ cpuregs.regs\[31\]\[14\] _01999_ _02000_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__mux4_1
XANTENNA__11811__A0 _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12543_ cpuregs.regs\[2\]\[6\] _06546_ _06752_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__mux2_1
XANTENNA__08902__S1 _03659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10395__S _04077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12176__A _06156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11080__A _05218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18050_ clknet_leaf_45_clk _01155_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_53_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10090__A2 _04021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15262_ cpuregs.regs\[4\]\[10\] cpuregs.regs\[5\]\[10\] cpuregs.regs\[6\]\[10\] cpuregs.regs\[7\]\[10\]
+ _02013_ _02014_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__mux4_1
X_12474_ _06141_ cpuregs.regs\[28\]\[6\] _06715_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17001_ clknet_leaf_141_clk _00175_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_14213_ reg_next_pc\[5\] _05834_ _07901_ _07916_ VGND VGND VPWR VPWR _07917_ sky130_fd_sc_hd__o211a_2
XFILLER_0_152_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11425_ _03305_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__buf_2
X_15193_ _03669_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__buf_6
XANTENNA__09232__A1 _03895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11410__A1_N _06003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 _02070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09232__B2 _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10917__A2 _05213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14144_ count_instr\[49\] _07865_ _07826_ VGND VGND VPWR VPWR _07867_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09485__A _04216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08586__A3 _03364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11356_ _05969_ _03851_ _05970_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10307_ reg_pc\[26\] decoded_imm\[26\] VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__or2_1
XANTENNA__15400__S1 _03643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14075_ count_instr\[28\] _07814_ _07790_ VGND VGND VPWR VPWR _07819_ sky130_fd_sc_hd__o21ai_1
X_11287_ _05904_ _05906_ _05911_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_167_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17903_ clknet_leaf_87_clk _01072_ VGND VGND VPWR VPWR count_cycle\[48\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11878__A0 _06078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13026_ cpuregs.regs\[3\]\[20\] _06575_ _07032_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__mux2_1
X_10238_ _04821_ _04876_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__or2b_1
XANTENNA__09940__C1 _04188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10169_ irq_pending\[21\] _04008_ _04874_ _04883_ VGND VGND VPWR VPWR _08382_ sky130_fd_sc_hd__o22a_1
X_17834_ clknet_leaf_58_clk _01003_ VGND VGND VPWR VPWR reg_next_pc\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16111__A _02770_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17765_ clknet_leaf_92_clk _00934_ VGND VGND VPWR VPWR count_instr\[36\] sky130_fd_sc_hd__dfxtp_1
X_14977_ irq_mask\[1\] _01864_ _01867_ _08335_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15950__A _03305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13928_ _03356_ _07704_ _07705_ net137 VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16716_ _06982_ cpuregs.regs\[19\]\[19\] _03087_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__mux2_1
X_17696_ clknet_leaf_39_clk _00865_ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dfxtp_2
XANTENNA__09394__S1 _04073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_164_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16033__A2 _02711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16647_ _03060_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15467__S1 _01997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13859_ cpuregs.regs\[0\]\[26\] VGND VGND VPWR VPWR _07669_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16578_ _06980_ cpuregs.regs\[18\]\[18\] _03015_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10605__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15219__S1 _02070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18317_ clknet_leaf_38_clk _01385_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_179_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15529_ _01969_ _02355_ _02363_ _02027_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__o211a_2
XFILLER_0_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09379__B decoded_imm\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09050_ net55 mem_rdata_q\[2\] _03729_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18248_ clknet_leaf_23_clk _01319_ VGND VGND VPWR VPWR decoded_imm\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_154_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16741__A0 _07007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18179_ clknet_leaf_22_clk _01250_ VGND VGND VPWR VPWR decoded_imm_j\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09774__A2 _04466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08982__A0 mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09952_ cpu_state\[6\] _04672_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_38_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12025__S _06460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10334__A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11869__A0 _06336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08903_ _03666_ _03667_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__or2_1
XANTENNA__10216__S0 _04472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09883_ _03385_ _04600_ _04601_ _04605_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__a31o_1
XANTENNA__10136__A3 _04847_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08834_ _03434_ _03599_ _03596_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08739__A net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08765_ _03530_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15860__A _02613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08696_ net112 net80 VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12695__S _06836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14476__A decoded_imm_j\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13380__A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12046__A0 _06216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15783__A1 _03298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14195__B _03196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13794__A0 _05143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10057__C1 _04237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09317_ _00072_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_97_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_934 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15535__A1 _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09248_ mem_rdata_q\[28\] _03987_ _03757_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
X_09179_ _03916_ _03922_ _03925_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11210_ _04360_ _05849_ _05827_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12190_ cpuregs.regs\[24\]\[12\] _06559_ _06555_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__mux2_1
XANTENNA__10455__S0 _04232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11141_ _03407_ _05286_ net130 _04422_ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__a22o_2
XANTENNA__10244__A reg_pc\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15394__S0 _01936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16630__S _03051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput77 net77 VGND VGND VPWR VPWR cpi_rs1[19] sky130_fd_sc_hd__buf_1
X_11072_ _03448_ _05397_ _05221_ _03447_ _05646_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__o221a_1
Xoutput88 net88 VGND VGND VPWR VPWR cpi_rs1[29] sky130_fd_sc_hd__clkbuf_1
XANTENNA__14510__A2 _07948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput99 net99 VGND VGND VPWR VPWR cpi_rs2[0] sky130_fd_sc_hd__clkbuf_1
X_10023_ _04018_ count_cycle\[49\] _04009_ _04741_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__a211o_1
X_14900_ _01823_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__16799__A0 _06582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15146__S0 _01999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15880_ _02632_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__16263__A2 _07944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14831_ count_cycle\[45\] _01771_ _01723_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15770__A _02484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11088__A1 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17550_ clknet_leaf_136_clk _00719_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14762_ _01726_ _08350_ _01727_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__and3b_1
X_11974_ _06201_ cpuregs.regs\[21\]\[13\] _06435_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__mux2_1
X_16501_ _02983_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13713_ net83 decoded_imm\[24\] VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__or2_1
XANTENNA__15449__S1 _02086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10925_ _03485_ _03564_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__or2_1
X_17481_ clknet_leaf_186_clk _00650_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_123_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14693_ count_cycle\[0\] count_cycle\[1\] count_cycle\[2\] VGND VGND VPWR VPWR _08337_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_123_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16432_ _06970_ cpuregs.regs\[29\]\[13\] _02943_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__mux2_1
XANTENNA__11803__A cpuregs.waddr\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13644_ _07490_ _07491_ VGND VGND VPWR VPWR _07492_ sky130_fd_sc_hd__xnor2_1
X_10856_ _05298_ _05538_ _05547_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14577__A2 _07954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16363_ _02910_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__clkbuf_1
X_13575_ _03387_ _04631_ VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__nor2_1
XANTENNA__14982__C1 _08335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10787_ _05225_ _05470_ _05474_ _05482_ VGND VGND VPWR VPWR alu_out\[8\] sky130_fd_sc_hd__a211o_1
XANTENNA__10599__B1 _05220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16805__S _03138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18102_ clknet_leaf_91_clk _01206_ VGND VGND VPWR VPWR timer\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15314_ _01989_ _02160_ _03639_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10063__A2 _04753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12526_ _06343_ cpuregs.regs\[28\]\[31\] _06714_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__mux2_1
XANTENNA__10694__S0 _05277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16294_ _02873_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18033_ clknet_leaf_66_clk _00009_ VGND VGND VPWR VPWR irq_pending\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13537__B1 _07211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11949__S _06424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15245_ _02094_ _02095_ _03687_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15621__S1 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12457_ cpuregs.regs\[27\]\[31\] _06598_ _06677_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09205__B2 _03888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output91_A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11012__A1 _05461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15010__A _04659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12813__A_N _06081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11408_ _05981_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13449__B decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15176_ _03649_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__buf_6
X_12388_ cpuregs.regs\[26\]\[31\] _06598_ _06640_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__mux2_1
XANTENNA__08550__C _03327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08964__B1 _03726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14127_ count_instr\[44\] _07852_ VGND VGND VPWR VPWR _07855_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11339_ _05174_ _05838_ _05955_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__a21bo_1
X_14058_ count_instr\[23\] _07805_ _07775_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10749__S1 _05288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13465__A _03518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13009_ cpuregs.regs\[3\]\[12\] _06559_ _07021_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__mux2_1
X_17817_ clknet_leaf_64_clk _00986_ VGND VGND VPWR VPWR reg_pc\[25\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_143_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15680__A _04335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08550_ _03325_ _03326_ _03327_ _03328_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__or4_1
X_17748_ clknet_leaf_86_clk _00917_ VGND VGND VPWR VPWR count_instr\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08481_ _03261_ _03262_ _03263_ _03264_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__or4_1
XFILLER_0_159_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14296__A irq_pending\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17679_ clknet_leaf_116_clk _00848_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11713__A _06265_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12579__A1 _06582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_28_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09102_ _03782_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16714__A0 _06980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15839__B _03885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11859__S _06370_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09033_ mem_rdata_q\[22\] net47 _03227_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_954 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16016__A is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15855__A _03305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15376__S0 _01908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09935_ _04654_ _04655_ _04320_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15066__S _03664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09866_ _04587_ _04588_ _04064_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__mux2_1
XANTENNA__15128__S0 _01982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08817_ net86 VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ cpuregs.regs\[16\]\[11\] cpuregs.regs\[17\]\[11\] cpuregs.regs\[18\]\[11\]
+ cpuregs.regs\[19\]\[11\] _04325_ _04277_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08748_ net130 net98 VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__nand2_1
XANTENNA__09358__S1 _04091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08679_ _03443_ _03444_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12019__A0 _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13314__S _07176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10710_ _03527_ _05389_ _03528_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11690_ reg_out\[19\] alu_out_q\[19\] _06068_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13767__B1 decoded_imm\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10641_ _04033_ _05237_ _05232_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11342__B _05957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16625__S _03040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13360_ _07226_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15508__A1 _01989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10572_ _05274_ _05275_ _05240_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__mux2_1
XANTENNA__09986__A2 _04016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_165_Right_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12990__A1 _06540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12311_ cpuregs.regs\[25\]\[27\] _06590_ _06626_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16181__A1 net246 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13291_ _06978_ cpuregs.regs\[5\]\[17\] _07165_ VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15030_ _03303_ _04022_ _04979_ _01897_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__a31o_1
X_12242_ cpuregs.regs\[24\]\[29\] _06594_ _06576_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12742__A1 cpuregs.waddr\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12742__B2 _06861_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15367__S0 _02022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16360__S _02907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12173_ _06149_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11124_ _03438_ _05783_ _03595_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__a21o_1
X_16981_ clknet_leaf_119_clk _00155_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__14495__A1 _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11055_ _03451_ _05397_ _05221_ _03450_ _05646_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__o221a_1
X_15932_ mem_rdata_q\[29\] mem_rdata_q\[24\] mem_rdata_q\[31\] mem_rdata_q\[30\] VGND
+ VGND VPWR VPWR _02658_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_155_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09371__B1 _04105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10006_ cpuregs.regs\[28\]\[17\] cpuregs.regs\[29\]\[17\] cpuregs.regs\[30\]\[17\]
+ cpuregs.regs\[31\]\[17\] _04072_ _04074_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__mux4_1
X_15863_ _02621_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__clkbuf_2
X_18651_ clknet_leaf_167_clk _01711_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11517__B latched_compr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output227_A net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15444__B1 _02197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11009__S _05277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14814_ _01762_ _01763_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__nor2_1
X_17602_ clknet_leaf_188_clk _00771_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_18582_ clknet_leaf_52_clk _01647_ VGND VGND VPWR VPWR reg_sh\[1\] sky130_fd_sc_hd__dfxtp_1
X_15794_ latched_branch _02578_ _02581_ _06026_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__o211a_1
XANTENNA__15995__A1 _03885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15995__B2 _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14828__B _01753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14745_ _01714_ _01715_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__nor2_1
X_17533_ clknet_leaf_114_clk _00702_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11957_ _06132_ cpuregs.regs\[21\]\[5\] _06424_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__mux2_1
XANTENNA__11533__A _06104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14547__C _07950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10908_ _05557_ _05316_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__nand2_1
XANTENNA__15005__A _04592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17464_ clknet_leaf_164_clk _00633_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14676_ _07898_ _07969_ _08050_ _07904_ reg_next_pc\[30\] VGND VGND VPWR VPWR _08324_
+ sky130_fd_sc_hd__a32o_1
X_11888_ _06132_ cpuregs.regs\[20\]\[5\] _06387_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08545__C _03322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16415_ _06953_ cpuregs.regs\[29\]\[5\] _02932_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__mux2_1
X_13627_ _07474_ _07475_ VGND VGND VPWR VPWR _07476_ sky130_fd_sc_hd__xnor2_1
X_10839_ _05219_ _05521_ _05526_ _05531_ VGND VGND VPWR VPWR alu_out\[11\] sky130_fd_sc_hd__o211ai_4
X_17395_ clknet_leaf_153_clk _00564_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16535__S _02967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16346_ _02901_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__clkbuf_1
X_13558_ _03566_ _05258_ VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10587__A3 _04708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12509_ _06740_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__clkbuf_1
X_16277_ _02864_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__clkbuf_1
X_13489_ _07345_ _07346_ _03631_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15228_ decoded_imm\[8\] _02009_ _01963_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__a21o_1
XANTENNA__14183__B1 _07877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18016_ clknet_leaf_104_clk _00001_ VGND VGND VPWR VPWR irq_pending\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10419__S0 _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08937__B1 _03675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15159_ _01936_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__buf_8
XANTENNA__16270__S _02859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09720_ _04133_ _04438_ _04446_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__and3_4
XANTENNA__09588__S1 _04317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12303__S _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09651_ _04214_ _04379_ _04081_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__a21o_1
X_08602_ _03378_ _03379_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__nand2_1
X_09582_ irq_pending\[5\] _04008_ _04312_ VGND VGND VPWR VPWR _08396_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08533_ cpu_state\[4\] VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13461__A2 _07211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13134__S _07082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11472__A1 _06054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08464_ net66 _03247_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__nand2_2
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10059__A _04776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14410__A1 _08071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10027__A2 _04745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08752__A net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16163__A1 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14174__B1 _07877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09016_ _03758_ _03763_ _03770_ _03777_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15910__A1 instr_slli VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10506__B instr_slli VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10735__B1 _05218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15674__B1 _02488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09918_ reg_pc\[15\] decoded_imm\[15\] VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10522__A net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10499__C1 _03302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11337__B _05948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09849_ _04018_ count_cycle\[45\] _04014_ count_cycle\[13\] _04571_ VGND VGND VPWR
+ VPWR _04572_ sky130_fd_sc_hd__a221o_1
XANTENNA__11160__A0 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12860_ _06266_ cpuregs.regs\[6\]\[21\] _06928_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__mux2_1
XANTENNA__15521__S0 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09105__B1 _03864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11811_ _06105_ cpuregs.regs\[11\]\[2\] _06348_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__mux2_1
XANTENNA__13552__B decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12791_ cpuregs.regs\[9\]\[21\] _06578_ _06891_ VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08646__B _03394_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13044__S _07032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14530_ _08177_ _08180_ _08189_ VGND VGND VPWR VPWR _08190_ sky130_fd_sc_hd__a21o_1
XANTENNA__15729__A1 _04777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11742_ reg_pc\[25\] _06283_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_120_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14461_ _08104_ _08114_ _08124_ _08107_ _08125_ VGND VGND VPWR VPWR _08126_ sky130_fd_sc_hd__o221a_1
X_11673_ _03409_ _03348_ _06066_ _06229_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__a22o_1
XANTENNA__16355__S _02896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14664__A _07968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16200_ _03730_ _02678_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__nor2_1
X_13412_ _04037_ _05260_ _07273_ _07274_ VGND VGND VPWR VPWR _07275_ sky130_fd_sc_hd__o211a_1
X_10624_ _05325_ _05326_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10649__S0 _05239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09959__A2 decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17180_ clknet_leaf_12_clk _00354_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09503__S1 _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14392_ _08052_ _08058_ _08057_ _08062_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__and4_1
XFILLER_0_52_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14383__B _03378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16131_ net290 net126 _02771_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13343_ instr_lui _07209_ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__nor2_2
X_10555_ _05258_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__16154__A1 net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10974__A0 _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14165__B1 _07877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16062_ _03402_ decoded_imm_j\[19\] _03403_ mem_rdata_q\[19\] VGND VGND VPWR VPWR
+ _02744_ sky130_fd_sc_hd__a22o_1
X_13274_ _06961_ cpuregs.regs\[5\]\[9\] _07154_ VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10486_ _04206_ _05190_ _04225_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__a21oi_1
X_15013_ irq_mask\[16\] _01880_ _01888_ _01876_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__a211o_1
XANTENNA_output177_A net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12225_ _06583_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09493__A _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12156_ cpuregs.regs\[24\]\[1\] _06536_ _06534_ VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11107_ _05554_ _05700_ _05775_ _05781_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__o211a_1
XANTENNA__13219__S _07129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11528__A _06098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10432__A _05138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16964_ clknet_leaf_115_clk _00138_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12087_ _06105_ cpuregs.regs\[23\]\[2\] _06496_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16209__A2 _06862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11038_ _05477_ _05487_ _05254_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__o21bai_2
X_15915_ _02610_ _02647_ _02651_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__and3_1
X_16895_ clknet_leaf_34_clk _00040_ VGND VGND VPWR VPWR mem_rdata_q\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13663__B1_N _07225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13345__A1_N _03387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18634_ clknet_leaf_146_clk _01694_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15968__A1 net262 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15846_ _03804_ _03794_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13979__B1 _07681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18565_ clknet_leaf_138_clk _01630_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_15777_ _02569_ _02567_ _02486_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12989_ _07013_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17516_ clknet_leaf_162_clk _00685_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_14728_ count_cycle\[13\] _08359_ _07826_ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18496_ clknet_leaf_157_clk _01561_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17447_ clknet_leaf_181_clk _00616_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12793__S _06891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14659_ _08288_ _08306_ _08307_ VGND VGND VPWR VPWR _08308_ sky130_fd_sc_hd__and3_1
XFILLER_0_172_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_180_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_180_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_171_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17378_ clknet_leaf_189_clk _00547_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16329_ _02891_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_870 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput201 net201 VGND VGND VPWR VPWR mem_la_addr[17] sky130_fd_sc_hd__buf_1
XFILLER_0_3_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput212 net212 VGND VGND VPWR VPWR mem_la_addr[28] sky130_fd_sc_hd__buf_1
XFILLER_0_140_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11509__A2 latched_store VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15609__S _02110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput223 net223 VGND VGND VPWR VPWR mem_la_addr[9] sky130_fd_sc_hd__buf_1
XFILLER_0_113_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput234 net234 VGND VGND VPWR VPWR mem_la_wdata[18] sky130_fd_sc_hd__buf_1
XANTENNA__10717__A0 _03524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput245 net245 VGND VGND VPWR VPWR mem_la_wdata[28] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput256 net256 VGND VGND VPWR VPWR mem_la_wdata[9] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput267 net267 VGND VGND VPWR VPWR mem_wdata[13] sky130_fd_sc_hd__clkbuf_1
Xoutput278 net278 VGND VGND VPWR VPWR mem_wdata[23] sky130_fd_sc_hd__clkbuf_1
Xoutput289 net289 VGND VGND VPWR VPWR mem_wdata[4] sky130_fd_sc_hd__buf_1
XFILLER_0_10_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12033__S _06460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09703_ _04369_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11142__B1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12968__S _06985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15408__B1 _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13653__A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09634_ net62 net258 _04035_ net48 _04362_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__a221o_2
XANTENNA__15959__A1 _03757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08747__A net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09565_ _04237_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__buf_6
XFILLER_0_167_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08516_ mem_wordsize\[2\] VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_65_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09496_ cpuregs.regs\[4\]\[4\] cpuregs.regs\[5\]\[4\] cpuregs.regs\[6\]\[4\] cpuregs.regs\[7\]\[4\]
+ _04207_ _04208_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08447_ _03230_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_171_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_171_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__15187__A2 _01906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08482__A instr_beq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09497__S0 _04207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12208__S _06555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09810__A1 _04391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10340_ reg_pc\[27\] decoded_imm\[27\] VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10271_ _03638_ _04959_ _04752_ _04960_ _04982_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12010_ _06457_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09574__B1 _04225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_307 VGND VGND VPWR VPWR alphacore_307/HI cpi_insn[5] sky130_fd_sc_hd__conb_1
Xalphacore_318 VGND VGND VPWR VPWR alphacore_318/HI cpi_insn[16] sky130_fd_sc_hd__conb_1
Xalphacore_329 VGND VGND VPWR VPWR alphacore_329/HI cpi_insn[27] sky130_fd_sc_hd__conb_1
XFILLER_0_100_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15111__A2 _03726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13961_ _03347_ _07727_ _07728_ net148 VGND VGND VPWR VPWR _07740_ sky130_fd_sc_hd__a22o_1
XANTENNA__15762__B _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15700_ _01881_ _02479_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__nand2_1
X_12912_ _06961_ cpuregs.regs\[31\]\[9\] _06943_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__mux2_1
X_16680_ _03078_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__clkbuf_1
X_13892_ _03327_ _07678_ _07682_ net157 VGND VGND VPWR VPWR _07692_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_85_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ _02459_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__clkbuf_1
X_12843_ _06201_ cpuregs.regs\[6\]\[13\] _06917_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12179__A _06165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14622__A1 _07998_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15562_ _02393_ _02394_ _01907_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__mux2_1
X_18350_ clknet_leaf_35_clk _01418_ VGND VGND VPWR VPWR mem_rdata_q\[5\] sky130_fd_sc_hd__dfxtp_1
X_12774_ cpuregs.regs\[9\]\[13\] _06561_ _06880_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17301_ clknet_leaf_113_clk _00475_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_14513_ _08141_ _08172_ VGND VGND VPWR VPWR _08174_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11725_ reg_pc\[23\] _06268_ _06093_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18281_ clknet_leaf_43_clk _00035_ VGND VGND VPWR VPWR is_sltiu_bltu_sltu sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15493_ _03639_ _02325_ _02329_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16085__S _03635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_162_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_162_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14394__A _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17232_ clknet_leaf_110_clk _00406_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_14444_ _08102_ _08103_ _08109_ _08110_ VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_154_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11656_ _06186_ reg_next_pc\[15\] _06212_ _06214_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__a211o_2
XFILLER_0_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09488__S0 _04217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10607_ _05307_ _05308_ _05309_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17163_ clknet_leaf_150_clk _00337_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16127__A1 _05414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14375_ _06863_ _08036_ _07919_ VGND VGND VPWR VPWR _08047_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10947__A0 _04754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08604__A2 irq_active VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11587_ reg_out\[8\] alu_out_q\[8\] _06067_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__mux2_1
XANTENNA__12118__S _06507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11022__S _05230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14138__B1 _07834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16114_ _03199_ _02674_ _02676_ _02673_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__o31a_1
X_13326_ cpuregs.regs\[24\]\[0\] cpuregs.regs\[25\]\[0\] cpuregs.regs\[26\]\[0\] cpuregs.regs\[27\]\[0\]
+ _04758_ _04759_ VGND VGND VPWR VPWR _07193_ sky130_fd_sc_hd__mux4_1
X_10538_ net121 VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15335__C1 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17094_ clknet_leaf_139_clk _00268_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11957__S _06424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10972__A1_N _05220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16045_ _02715_ decoded_imm_j\[11\] mem_rdata_q\[7\] _03309_ _02633_ VGND VGND VPWR
+ VPWR _02735_ sky130_fd_sc_hd__a221o_1
XANTENNA__10861__S _05363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13738__A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13257_ _07155_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__clkbuf_1
X_10469_ net56 _04745_ _04666_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09427__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12208_ cpuregs.regs\[24\]\[18\] _06571_ _06555_ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__mux2_1
XANTENNA__13457__B _05257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13188_ _06941_ cpuregs.regs\[8\]\[0\] _07118_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__mux2_1
X_12139_ _06312_ cpuregs.regs\[23\]\[27\] _06518_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__mux2_1
XANTENNA__13649__C1 _07274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17996_ clknet_leaf_65_clk _01133_ VGND VGND VPWR VPWR irq_mask\[12\] sky130_fd_sc_hd__dfxtp_1
X_16947_ clknet_leaf_61_clk _00075_ VGND VGND VPWR VPWR cpu_state\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13664__A2 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10478__A2 _04012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12872__A0 _06312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16878_ _03183_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08540__A1 decoder_trigger VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18617_ clknet_leaf_16_clk _00091_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__dfxtp_4
X_15829_ decoded_imm_j\[16\] _05987_ _03910_ _02587_ _02596_ VGND VGND VPWR VPWR _01246_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14613__A1 _07958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15810__B1 _03954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12624__A0 _06193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09350_ _04084_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__buf_8
XANTENNA__09715__S1 _04074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18548_ clknet_leaf_170_clk _01613_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09281_ _04017_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__buf_4
XFILLER_0_145_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_153_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_153_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18479_ clknet_leaf_20_clk _01544_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16723__S _03098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15877__A0 instr_jalr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11867__S _06370_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13648__A _04959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10166__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15629__B1 _01932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08996_ mem_rdata_q\[31\] _03756_ _03757_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09861__A _04369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11318__D _05937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10469__A2 _04745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10013__S1 _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11130__A3 _05086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09617_ reg_pc\[6\] decoded_imm\[6\] VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09548_ cpuregs.regs\[12\]\[5\] cpuregs.regs\[13\]\[5\] cpuregs.regs\[14\]\[5\] cpuregs.regs\[15\]\[5\]
+ _04275_ _04278_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__mux4_1
XANTENNA__09706__S1 _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_144_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_144_clk sky130_fd_sc_hd__clkbuf_2
X_09479_ _04078_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__buf_8
XANTENNA__08834__A2 _03599_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11631__A _06192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11510_ cpuregs.waddr\[2\] _06081_ _06082_ _06083_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_108_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10641__A2 _05237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12490_ _06730_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11441_ irq_mask\[10\] _06030_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_22_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11350__B _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10247__A net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14942__A _01823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14160_ _07876_ _07878_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11372_ _03895_ _05962_ _05967_ _05981_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_150_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14661__B _07968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13111_ _07077_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10323_ cpuregs.regs\[0\]\[26\] cpuregs.regs\[1\]\[26\] cpuregs.regs\[2\]\[26\] cpuregs.regs\[3\]\[26\]
+ _04055_ _04058_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_78_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10681__S _05239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14091_ _07828_ _07815_ _07829_ VGND VGND VPWR VPWR _07830_ sky130_fd_sc_hd__and3b_1
XFILLER_0_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13042_ cpuregs.regs\[3\]\[28\] _06592_ _07032_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__mux2_1
X_10254_ _04211_ _04963_ _04965_ _04328_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__o211a_1
XANTENNA__10157__B2 _04024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17850_ clknet_leaf_107_clk _01019_ VGND VGND VPWR VPWR reg_next_pc\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10252__S1 _04376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10185_ cpuregs.regs\[0\]\[22\] cpuregs.regs\[1\]\[22\] cpuregs.regs\[2\]\[22\] cpuregs.regs\[3\]\[22\]
+ _04056_ _04091_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__mux4_1
XANTENNA__16293__A0 _06968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16801_ _06584_ cpuregs.regs\[13\]\[24\] _03138_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__mux2_1
X_17781_ clknet_leaf_86_clk _00950_ VGND VGND VPWR VPWR count_instr\[52\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13646__A2 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15191__S1 _03647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14389__A decoded_imm_j\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14993_ _04414_ _01869_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__nor2_1
X_16732_ _03105_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__clkbuf_1
X_13944_ _07681_ VGND VGND VPWR VPWR _07728_ sky130_fd_sc_hd__buf_2
XANTENNA__12401__S _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16045__B1 mem_rdata_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13875_ _03292_ cpu_state\[2\] VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__nand2_2
X_16663_ cpuregs.regs\[1\]\[26\] _06303_ _03062_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__mux2_1
X_18402_ clknet_leaf_137_clk _01467_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_157_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15614_ _03709_ _02442_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__or2_1
X_12826_ _06132_ cpuregs.regs\[6\]\[5\] _06906_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__mux2_1
XANTENNA__13803__C1 _07221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16594_ _03032_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09710__S _04321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18333_ clknet_leaf_35_clk _01401_ VGND VGND VPWR VPWR mem_16bit_buffer\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15545_ _02377_ _02378_ _03713_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__mux2_1
X_12757_ cpuregs.regs\[9\]\[5\] _06544_ _06869_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_135_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_135_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16109__A mem_do_wdata VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13232__S _07140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11708_ reg_pc\[20\] reg_pc\[19\] _06234_ reg_pc\[21\] VGND VGND VPWR VPWR _06261_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15476_ decoded_imm\[22\] _02216_ _02197_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18264_ clknet_leaf_26_clk _01335_ VGND VGND VPWR VPWR decoded_imm\[22\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_155_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12688_ _06824_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__buf_6
XFILLER_0_86_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11260__B _05881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17215_ clknet_leaf_179_clk _00389_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_14427_ _08087_ _08094_ VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11639_ _06186_ reg_next_pc\[13\] _06197_ _06199_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__a211o_4
XFILLER_0_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18195_ clknet_leaf_41_clk _01266_ VGND VGND VPWR VPWR instr_sb sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16543__S _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14374__A3 _07992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17146_ clknet_leaf_187_clk _00320_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14358_ _03368_ _08027_ _08028_ _08031_ VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__a31o_1
XFILLER_0_170_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10396__A1 _04052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13309_ _07182_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17077_ clknet_leaf_116_clk _00251_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14289_ reg_pc\[29\] _07953_ _07968_ _07960_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__a22o_1
XANTENNA__09665__B decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10491__S1 _04218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09538__B1 _04017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16028_ decoded_imm\[4\] _02720_ _02723_ _02724_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08850_ _03608_ _03521_ _03612_ _03615_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__or4_1
XFILLER_0_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08996__S _03757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08781_ net127 net95 VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__and2b_1
X_17979_ clknet_leaf_43_clk _01116_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13604__A2_N _04702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10620__A _05322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12311__S _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09402_ cpuregs.regs\[4\]\[2\] cpuregs.regs\[5\]\[2\] cpuregs.regs\[6\]\[2\] cpuregs.regs\[7\]\[2\]
+ _04071_ _04073_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15795__C1 _03305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09333_ _00072_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__inv_6
XFILLER_0_158_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1004 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_126_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_126_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__16019__A mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09264_ _03737_ _04001_ _03763_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_146_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16453__S _02954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09195_ _03916_ _03925_ _03941_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13573__A1 _04466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_985 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09856__A _04487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11584__A0 _06150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13378__A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10139__A1 _04018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11336__B1 _05952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13089__A0 _06980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09591__A _04320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08979_ mem_rdata_q\[30\] net56 _03208_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__mux2_1
XANTENNA__11639__A1 _06186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12221__S _06576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09927__S1 _04087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11990_ _06447_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09701__B1 _04018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10941_ _03488_ _05612_ _03568_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13660_ _07501_ _07506_ VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__nand2_1
XANTENNA__14589__B1 _08071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10872_ _05287_ _05562_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_27_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12611_ _06141_ cpuregs.regs\[30\]\[6\] _06788_ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13591_ _07437_ _07440_ _07442_ _07284_ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_117_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_117_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_155_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13052__S _07046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15330_ _02012_ _02175_ _02017_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12542_ _06758_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_152_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15261_ _02110_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12891__S _06943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12473_ _06721_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14212_ _05856_ _06128_ VGND VGND VPWR VPWR _07916_ sky130_fd_sc_hd__or2_1
X_17000_ clknet_leaf_142_clk _00174_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11424_ _06026_ _06027_ _06028_ net12 VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__a31o_1
X_15192_ _03719_ _02044_ _00067_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__o21a_1
XANTENNA__08670__A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_8 _02166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14143_ _07865_ _07866_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_130_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11355_ _03199_ _03310_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__nand2_4
XANTENNA__12192__A _06200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10306_ reg_pc\[26\] decoded_imm\[26\] VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_394 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14074_ count_instr\[28\] count_instr\[27\] count_instr\[26\] _07811_ VGND VGND VPWR
+ VPWR _07818_ sky130_fd_sc_hd__and4_2
X_11286_ _05904_ _05906_ _05911_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output257_A net257 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17902_ clknet_leaf_87_clk _01071_ VGND VGND VPWR VPWR count_cycle\[47\] sky130_fd_sc_hd__dfxtp_1
X_13025_ _07009_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__buf_6
X_10237_ _04877_ _04886_ _04919_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_167_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17833_ clknet_leaf_57_clk _01002_ VGND VGND VPWR VPWR reg_next_pc\[10\] sky130_fd_sc_hd__dfxtp_1
X_10168_ _03384_ _04878_ _04879_ _04882_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__a31o_1
XANTENNA__08829__B net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13227__S _07129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15008__A _04631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17764_ clknet_leaf_92_clk _00933_ VGND VGND VPWR VPWR count_instr\[35\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12131__S _06518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10099_ _04749_ _04784_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_128_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14976_ _04101_ _01865_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_145_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16715_ _03096_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09006__A _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13927_ _07716_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15950__B mem_rdata_q\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17695_ clknet_leaf_169_clk _00864_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11970__S _06435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16646_ cpuregs.regs\[1\]\[18\] _06239_ _03051_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__mux2_1
X_13858_ _07668_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08845__A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13252__A0 _07007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12809_ cpuregs.regs\[9\]\[30\] _06596_ _06868_ VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09456__C1 _04188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16577_ _03023_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_108_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_108_clk sky130_fd_sc_hd__clkbuf_2
X_13789_ _05174_ _05086_ _05227_ VGND VGND VPWR VPWR _07627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18316_ clknet_leaf_36_clk _01384_ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dfxtp_1
X_15528_ _02357_ _02359_ _02362_ _02037_ _02006_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__a221o_1
XANTENNA__15529__C1 _02027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09471__A2 _04197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18247_ clknet_leaf_23_clk _01318_ VGND VGND VPWR VPWR decoded_imm\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_142_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15459_ _02020_ _02289_ _02297_ _01960_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__o211a_2
XFILLER_0_5_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10369__A1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18178_ clknet_leaf_31_clk _01249_ VGND VGND VPWR VPWR decoded_imm_j\[19\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_40_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10369__B2 _05077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17129_ clknet_leaf_134_clk _00303_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08982__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09951_ latched_is_lh _04670_ _04671_ _04420_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_38_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08902_ cpuregs.regs\[24\]\[2\] cpuregs.regs\[25\]\[2\] cpuregs.regs\[26\]\[2\] cpuregs.regs\[27\]\[2\]
+ _03658_ _03659_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _03637_ _04602_ _04604_ _03225_ _04266_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__a221o_1
XANTENNA__10216__S1 _04473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _03446_ _03591_ _03598_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08739__B net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08764_ net124 VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08695_ net112 net80 VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__or2_1
XFILLER_0_170_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11880__S _06387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13380__B decoded_imm\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15783__A2 _04006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09316_ instr_retirq VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10152__S0 _04579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09247_ _03754_ _03733_ _03731_ _03753_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__a22o_2
XFILLER_0_106_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16183__S _02770_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15091__S0 _03669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09586__A _04215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09178_ _03798_ _03853_ _03927_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15100__B _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10455__S1 _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15299__B2 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11140_ _03407_ _05324_ net129 _04422_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__a22o_2
XFILLER_0_101_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11309__A0 _05013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10244__B decoded_imm\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15394__S1 _01937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput67 net67 VGND VGND VPWR VPWR cpi_rs1[0] sky130_fd_sc_hd__buf_1
XANTENNA__15527__S _01907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput78 net78 VGND VGND VPWR VPWR cpi_rs1[1] sky130_fd_sc_hd__buf_1
X_11071_ _05277_ _05746_ _05747_ _05251_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__o211a_1
Xoutput89 net89 VGND VGND VPWR VPWR cpi_rs1[2] sky130_fd_sc_hd__clkbuf_1
X_10022_ count_instr\[49\] _04104_ _04011_ count_instr\[17\] VGND VGND VPWR VPWR _04741_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15146__S1 _02000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14830_ count_cycle\[43\] count_cycle\[44\] count_cycle\[45\] _01768_ VGND VGND VPWR
+ VPWR _01774_ sky130_fd_sc_hd__and4_2
XFILLER_0_98_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14761_ count_cycle\[22\] _01722_ count_cycle\[23\] VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__a21o_1
X_11973_ _06438_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16358__S _02907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16500_ cpuregs.regs\[17\]\[13\] _06561_ _02979_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__mux2_1
X_13712_ net83 decoded_imm\[24\] VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__nand2_1
X_10924_ _05279_ _05597_ _05607_ _05611_ VGND VGND VPWR VPWR alu_out\[16\] sky130_fd_sc_hd__a211o_1
XANTENNA__09150__B2 _03888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14692_ count_cycle\[0\] count_cycle\[1\] _08336_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__a21oi_1
X_17480_ clknet_leaf_13_clk _00649_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08665__A instr_beq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10391__S0 _04273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16431_ _02946_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__clkbuf_1
X_13643_ _07473_ _07475_ _07472_ VGND VGND VPWR VPWR _07491_ sky130_fd_sc_hd__a21boi_1
X_10855_ _05542_ _05546_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__nand2_1
XANTENNA__11803__B cpuregs.waddr\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13574_ _07190_ _07424_ _07426_ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__or3_1
X_16362_ _06968_ cpuregs.regs\[16\]\[12\] _02907_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10786_ _05476_ _05478_ _05399_ _05481_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_137_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18101_ clknet_leaf_90_clk _01205_ VGND VGND VPWR VPWR timer\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15313_ cpuregs.regs\[16\]\[13\] cpuregs.regs\[17\]\[13\] cpuregs.regs\[18\]\[13\]
+ cpuregs.regs\[19\]\[13\] _02013_ _02014_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__mux4_1
X_12525_ _06748_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16293_ _06968_ cpuregs.regs\[15\]\[12\] _02870_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13537__A1 _07209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18032_ clknet_leaf_80_clk _00008_ VGND VGND VPWR VPWR irq_pending\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15244_ cpuregs.regs\[20\]\[9\] cpuregs.regs\[21\]\[9\] cpuregs.regs\[22\]\[9\] cpuregs.regs\[23\]\[9\]
+ _02074_ _02075_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__mux4_1
X_12456_ _06711_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11407_ cpuregs.raddr1\[1\] _06006_ _06014_ _06015_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_169_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15010__B _01885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15175_ _02012_ _02028_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16821__S _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12387_ _06674_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11030__S _05390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output84_A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14126_ count_instr\[44\] _07852_ VGND VGND VPWR VPWR _07854_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11338_ _03229_ _05953_ _05954_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__or3_1
XANTENNA__08964__B2 _03638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11965__S _06424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15437__S _01907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14057_ _07805_ _07806_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__nor2_1
XANTENNA__13746__A _05037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11269_ _05876_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__buf_2
XANTENNA__16239__A0 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13008_ _07023_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09913__B1 _03252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13465__B decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17816_ clknet_leaf_68_clk _00985_ VGND VGND VPWR VPWR reg_pc\[24\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_50_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17747_ clknet_leaf_86_clk _00916_ VGND VGND VPWR VPWR count_instr\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12276__A1 _06554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15680__B _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14959_ net215 net184 _01846_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__mux2_1
XANTENNA__16268__S _02859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09141__A1 _03895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08480_ instr_ori instr_xori instr_addi instr_bgeu VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17678_ clknet_leaf_144_clk _00847_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16411__A0 _06949_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10382__S0 _04216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13225__A0 _06980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16629_ _03039_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13776__A1 _04959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11787__B1 _06101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09101_ _03853_ _03776_ _03855_ _03860_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15839__C _03895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09032_ mem_16bit_buffer\[5\] _03793_ _03727_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16016__B is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12036__S _06471_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16731__S _03098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15376__S1 _01909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09934_ cpuregs.regs\[8\]\[15\] cpuregs.regs\[9\]\[15\] cpuregs.regs\[10\]\[15\]
+ cpuregs.regs\[11\]\[15\] _04487_ _04469_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09865_ cpuregs.regs\[8\]\[13\] cpuregs.regs\[9\]\[13\] cpuregs.regs\[10\]\[13\]
+ cpuregs.regs\[11\]\[13\] _04280_ _04091_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__mux4_1
XANTENNA__15128__S1 _03639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08469__B instr_rdinstr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08816_ _03459_ _03581_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__or2_1
X_09796_ cpuregs.regs\[20\]\[11\] cpuregs.regs\[21\]\[11\] cpuregs.regs\[22\]\[11\]
+ cpuregs.regs\[23\]\[11\] _04325_ _04277_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__mux4_1
X_08747_ net130 net98 VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08678_ net120 net88 VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__nand2_2
XANTENNA__08485__A _03254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15205__A1 _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13767__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10640_ net89 _03242_ _03609_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11778__B1 _06101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10571_ net90 _05205_ _05229_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__mux2_1
XANTENNA__16207__A _04156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15064__S0 _03670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12310_ _06633_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13290_ _07172_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12241_ _06327_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__buf_2
XFILLER_0_106_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16469__A0 _07007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_163_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12742__A2 _06862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12172_ _06547_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15765__B _03425_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15367__S1 _02023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11123_ _03444_ _05785_ _03435_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13566__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16980_ clknet_leaf_105_clk _00154_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_164_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11054_ _05277_ _05730_ _05731_ _05251_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__o211a_1
X_15931_ instr_srai _02650_ _02657_ mem_rdata_q\[30\] VGND VGND VPWR VPWR _01287_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_178_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15781__A _07778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10005_ _04483_ _04723_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__nand2_1
X_18650_ clknet_leaf_163_clk _01710_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_15862_ _03309_ _03304_ _02610_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15444__A1 decoded_imm\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17601_ clknet_leaf_16_clk _00770_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14813_ count_cycle\[39\] _01759_ _01723_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__o21ai_1
X_18581_ clknet_leaf_52_clk _01646_ VGND VGND VPWR VPWR reg_sh\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_output122_A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09659__C1 _03301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15793_ _03302_ _02579_ _02580_ _02578_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__or4b_1
XFILLER_0_99_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15995__A2 _03880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17532_ clknet_leaf_107_clk _00701_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_14744_ count_cycle\[16\] count_cycle\[17\] count_cycle\[18\] _08365_ VGND VGND VPWR
+ VPWR _01715_ sky130_fd_sc_hd__and4_2
X_11956_ _06429_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10907_ _05361_ _05584_ _05585_ _05595_ VGND VGND VPWR VPWR alu_out\[15\] sky130_fd_sc_hd__a31o_1
XFILLER_0_129_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17463_ clknet_leaf_122_clk _00632_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_11887_ _06392_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14675_ _08321_ _08322_ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14955__A0 net212 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16414_ _02937_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13626_ _07459_ _07463_ VGND VGND VPWR VPWR _07475_ sky130_fd_sc_hd__nand2_1
X_10838_ _05399_ _05529_ _05530_ _05478_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08545__D _03323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17394_ clknet_leaf_140_clk _00563_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11769__B1 _06101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12430__A1 _06571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16345_ _06951_ cpuregs.regs\[16\]\[4\] _02896_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10769_ _05361_ _05453_ _05454_ _05465_ VGND VGND VPWR VPWR alu_out\[7\] sky130_fd_sc_hd__a31o_1
X_13557_ _04611_ _04566_ _05227_ VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15055__S0 _03658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13240__S _07140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14707__B1 _07877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12508_ _06274_ cpuregs.regs\[28\]\[22\] _06737_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13488_ _07345_ _07346_ VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__nor2_1
X_16276_ _06951_ cpuregs.regs\[15\]\[4\] _02859_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18015_ clknet_leaf_76_clk _01152_ VGND VGND VPWR VPWR irq_mask\[31\] sky130_fd_sc_hd__dfxtp_1
X_15227_ _01969_ _02065_ _02078_ _01960_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__o211a_4
X_12439_ cpuregs.regs\[27\]\[22\] _06580_ _06700_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__mux2_1
XANTENNA__10419__S1 _04478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16551__S _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08937__A1 _03657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15158_ _03653_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__buf_6
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14109_ _07842_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15089_ _03666_ _01947_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13694__A0 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09362__A1 _04070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15691__A _02486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09650_ _04377_ _04378_ _04222_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08601_ instr_jal _03367_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__nor2_2
XANTENNA__13446__A0 _04262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09581_ _03385_ _04261_ _04267_ _04311_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__a211o_1
X_08532_ _03238_ _03311_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10355__S0 _04057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08463_ mem_do_wdata _03218_ _03241_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15630__S _03272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13749__A1 _03276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15294__S0 _02069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09015_ _03776_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15371__B1 _02027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15910__A2 _02635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10075__A _04289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16461__S _02954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13921__A1 _03352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09050__A0 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10196__C1 _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16871__A0 _06586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09917_ irq_pending\[14\] _04049_ _04610_ _04638_ VGND VGND VPWR VPWR _08374_ sky130_fd_sc_hd__a211o_1
XANTENNA__16697__A _03075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_97_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__11337__C _05952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09848_ count_instr\[45\] _04016_ _04012_ count_instr\[13\] VGND VGND VPWR VPWR _04571_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11160__A1 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15426__A1 _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09779_ _04501_ _04502_ _04503_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__or3_1
XANTENNA__15521__S1 _01997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11810_ _06350_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15106__A _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12790_ _06892_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_103_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _06290_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11353__B _03864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16636__S _03051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11672_ reg_out\[17\] alu_out_q\[17\] _06068_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__mux2_1
X_14460_ decoded_imm_j\[12\] _07932_ VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10623_ _03535_ _03536_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__xnor2_1
X_13411_ _07216_ VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14391_ _08060_ _08061_ VGND VGND VPWR VPWR _08062_ sky130_fd_sc_hd__nand2_1
XANTENNA__10649__S1 _05237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13060__S _07046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_106_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16130_ _02782_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__clkbuf_1
X_13342_ is_lui_auipc_jal VGND VGND VPWR VPWR _07209_ sky130_fd_sc_hd__clkinv_4
X_10554_ _05257_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__buf_2
XFILLER_0_63_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10974__A1 _04810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15362__B1 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13273_ _07163_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__clkbuf_1
X_16061_ decoded_imm\[18\] _02720_ _02736_ _02743_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__o22a_1
X_10485_ _05188_ _05189_ _04321_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__mux2_1
XANTENNA__14680__A _07971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13912__A1 _03333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15012_ _04702_ _01885_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12224_ cpuregs.regs\[24\]\[23\] _06582_ _06576_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__mux2_1
X_12155_ _06095_ VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__buf_2
X_11106_ _05281_ _05777_ _05780_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__a21oi_1
X_12086_ _06498_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__clkbuf_1
X_16963_ clknet_leaf_130_clk _00137_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_88_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_2
X_11037_ _03456_ _05220_ _05600_ _05618_ _05715_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__a221o_1
X_15914_ _03277_ is_alu_reg_reg VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__and2_1
XANTENNA__15942__C mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16894_ clknet_leaf_35_clk _00039_ VGND VGND VPWR VPWR mem_rdata_q\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08822__A_N net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18633_ clknet_leaf_138_clk _01693_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_15845_ _02606_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08837__B _03600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15016__A _04776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13979__B2 net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18564_ clknet_leaf_143_clk _01629_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15776_ timer\[31\] VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12988_ cpuregs.regs\[3\]\[2\] _06538_ _07010_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17515_ clknet_leaf_127_clk _00684_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09014__A _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14727_ _08359_ _08360_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11454__A2 irq_pending\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18495_ clknet_leaf_131_clk _01560_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11939_ _06419_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15276__S0 _01985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14928__A0 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_276 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17446_ clknet_leaf_167_clk _00615_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14658_ _07966_ _07967_ _08232_ VGND VGND VPWR VPWR _08307_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13609_ net75 decoded_imm\[17\] VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17377_ clknet_leaf_17_clk _00546_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14589_ _08241_ _08243_ _08071_ VGND VGND VPWR VPWR _08244_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_172_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__10414__B1 _04014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16328_ _07003_ cpuregs.regs\[15\]\[29\] _02881_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_922 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15353__B1 _02197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16259_ mem_rdata_q\[6\] _03878_ _03914_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput202 net202 VGND VGND VPWR VPWR mem_la_addr[18] sky130_fd_sc_hd__buf_1
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput213 net213 VGND VGND VPWR VPWR mem_la_addr[29] sky130_fd_sc_hd__buf_1
XFILLER_0_113_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11509__A3 _03195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput224 net224 VGND VGND VPWR VPWR mem_la_read sky130_fd_sc_hd__clkbuf_1
Xoutput235 net235 VGND VGND VPWR VPWR mem_la_wdata[19] sky130_fd_sc_hd__buf_1
XANTENNA__10717__A1 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput246 net246 VGND VGND VPWR VPWR mem_la_wdata[29] sky130_fd_sc_hd__buf_1
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput257 net257 VGND VGND VPWR VPWR mem_la_write sky130_fd_sc_hd__clkbuf_1
XANTENNA__15105__B1 _01962_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput268 net268 VGND VGND VPWR VPWR mem_wdata[14] sky130_fd_sc_hd__clkbuf_1
Xoutput279 net279 VGND VGND VPWR VPWR mem_wdata[24] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_79_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_156_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09702_ count_instr\[41\] _04016_ count_cycle\[9\] _04014_ _04428_ VGND VGND VPWR
+ VPWR _04429_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11142__A1 _03407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16605__A0 _07007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15408__A1 _01959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11142__B2 _04422_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15408__B2 decoded_imm\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13653__B decoded_imm\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09633_ _03242_ net39 _04361_ net67 mem_wordsize\[1\] VGND VGND VPWR VPWR _04362_
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__08747__B net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13145__S _07093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16081__A1 decoded_imm\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16081__B2 mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09564_ _04293_ _04294_ _04223_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08515_ _03296_ VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__buf_2
XFILLER_0_33_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09495_ net301 VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__buf_8
XANTENNA__12984__S _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14919__A0 net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08446_ mem_la_secondword _03229_ _03191_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__or3_2
XANTENNA__09859__A _04206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08482__B instr_waitirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09497__S1 _04208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15895__A1 is_alu_reg_imm VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10270_ _04268_ _04962_ _04981_ _04149_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__o211a_1
XANTENNA__10708__A1 _05255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09574__A1 _04289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xalphacore_308 VGND VGND VPWR VPWR alphacore_308/HI cpi_insn[6] sky130_fd_sc_hd__conb_1
XANTENNA__12224__S _06576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_319 VGND VGND VPWR VPWR alphacore_319/HI cpi_insn[17] sky130_fd_sc_hd__conb_1
XANTENNA__15647__A1 _03309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13960_ _07739_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12911_ _06165_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__buf_2
XANTENNA__10679__S _05239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13891_ _06053_ VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__16072__A1 decoded_imm\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14607__C1 _07898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15630_ net123 _02458_ _03272_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__mux2_1
XANTENNA__16072__B2 mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12842_ _06920_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10319__S0 _04071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15561_ cpuregs.regs\[8\]\[27\] cpuregs.regs\[9\]\[27\] cpuregs.regs\[10\]\[27\]
+ cpuregs.regs\[11\]\[27\] _02074_ _02075_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__mux4_1
X_12773_ _06883_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16366__S _02907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12894__S _06943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10644__A0 _04466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15258__S0 _01990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17300_ clknet_leaf_105_clk _00474_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08932__S0 _03641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14512_ _08140_ _08151_ _08172_ VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__or3_1
X_18280_ clknet_leaf_43_clk _00034_ VGND VGND VPWR VPWR is_slti_blt_slt sky130_fd_sc_hd__dfxtp_1
X_11724_ _06275_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__clkbuf_1
X_15492_ _03675_ _02328_ _03657_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17231_ clknet_leaf_124_clk _00405_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _03409_ _03356_ _06066_ _06213_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14443_ _08106_ _08108_ VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__nand2_1
XANTENNA__12195__A _06207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09488__S1 _04219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10606_ _05231_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__clkbuf_4
X_17162_ clknet_leaf_147_clk _00336_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14374_ _07899_ _07917_ _07992_ _08046_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__a31o_1
X_11586_ reg_pc\[8\] _06146_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10947__A1 _04744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16113_ _05829_ _02768_ _02772_ net193 VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__a22o_1
X_10537_ _04251_ _04262_ _04342_ _04360_ _05230_ _05240_ VGND VGND VPWR VPWR _05241_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_134_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13325_ cpuregs.regs\[28\]\[0\] cpuregs.regs\[29\]\[0\] cpuregs.regs\[30\]\[0\] cpuregs.regs\[31\]\[0\]
+ _04282_ _04285_ VGND VGND VPWR VPWR _07192_ sky130_fd_sc_hd__mux4_1
X_17093_ clknet_leaf_156_clk _00267_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15430__S0 _01979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15886__B2 is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16044_ is_sb_sh_sw _02712_ mem_rdata_q\[31\] VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__o21a_1
XANTENNA__13738__B decoded_imm\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10468_ net90 VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__clkbuf_4
X_13256_ _06941_ cpuregs.regs\[5\]\[0\] _07154_ VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12207_ _06239_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13187_ _07117_ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__buf_6
X_10399_ _05106_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__inv_2
XANTENNA__10175__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11372__A1 _03895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12138_ _06525_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__clkbuf_1
X_17995_ clknet_leaf_65_clk _01132_ VGND VGND VPWR VPWR irq_mask\[11\] sky130_fd_sc_hd__dfxtp_1
X_16946_ clknet_leaf_53_clk _00074_ VGND VGND VPWR VPWR cpu_state\[0\] sky130_fd_sc_hd__dfxtp_1
X_12069_ _06304_ cpuregs.regs\[22\]\[26\] _06482_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__08848__A net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16877_ _06592_ cpuregs.regs\[14\]\[28\] _03174_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16063__A1 decoded_imm\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15497__S0 _01970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18616_ clknet_leaf_9_clk _00090_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__dfxtp_1
X_15828_ decoded_imm_j\[15\] _05987_ _03781_ _02587_ _02596_ VGND VGND VPWR VPWR _01245_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__14613__A2 _07959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18547_ clknet_leaf_162_clk _01612_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_15759_ _02554_ _02555_ _02556_ _02545_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__o211a_1
XANTENNA__16276__S _02859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09280_ instr_rdcycleh VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18478_ clknet_leaf_106_clk _01543_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08583__A irq_active VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17429_ clknet_leaf_106_clk _00598_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12309__S _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12044__S _06471_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10166__A2 _04745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15629__A1 _01959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15629__B2 decoded_imm\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08995_ _03227_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_167_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08758__A net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08477__B instr_sub VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09616_ _04046_ _04342_ _04345_ _03225_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__a22o_1
XANTENNA__14065__B1 _07790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09547_ _04277_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__buf_4
XFILLER_0_167_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08493__A _03275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09478_ cpuregs.regs\[24\]\[4\] cpuregs.regs\[25\]\[4\] cpuregs.regs\[26\]\[4\] cpuregs.regs\[27\]\[4\]
+ _04207_ _04208_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__mux4_1
XFILLER_0_109_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15565__B1 _02197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08429_ _03214_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13576__C1 _07221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11440_ _06029_ irq_pending\[9\] _06037_ net32 VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_22_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13040__A1 _06590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11051__A0 _05044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11371_ _05970_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_150_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15412__S0 _03670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13110_ _07001_ cpuregs.regs\[7\]\[28\] _07068_ VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__mux2_1
X_10322_ cpuregs.regs\[4\]\[26\] cpuregs.regs\[5\]\[26\] cpuregs.regs\[6\]\[26\] cpuregs.regs\[7\]\[26\]
+ _04055_ _04058_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__mux4_1
X_14090_ count_instr\[32\] _07824_ count_instr\[33\] VGND VGND VPWR VPWR _07829_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13041_ _07040_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10253_ _04369_ _04964_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__or2_1
XANTENNA__10157__A2 _04448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15773__B _02560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10184_ _04054_ _04897_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__nand2_1
X_16800_ _03142_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__clkbuf_1
X_17780_ clknet_leaf_86_clk _00949_ VGND VGND VPWR VPWR count_instr\[51\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11106__A1 _05281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14992_ irq_mask\[7\] _01864_ _01875_ _01876_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__a211o_1
XANTENNA__09263__S _03757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16731_ _06997_ cpuregs.regs\[19\]\[26\] _03098_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__mux2_1
X_13943_ _07677_ VGND VGND VPWR VPWR _07727_ sky130_fd_sc_hd__buf_2
XFILLER_0_72_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16045__B2 _03309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10865__B1 _05357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16662_ _03068_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__clkbuf_1
X_13874_ _07677_ VGND VGND VPWR VPWR _07678_ sky130_fd_sc_hd__buf_2
XANTENNA__14056__B1 _07790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15253__C1 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18401_ clknet_leaf_157_clk _01466_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15613_ cpuregs.regs\[16\]\[31\] cpuregs.regs\[17\]\[31\] cpuregs.regs\[18\]\[31\]
+ cpuregs.regs\[19\]\[31\] _01995_ _01937_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__mux4_1
X_12825_ _06911_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output202_A net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16593_ _06995_ cpuregs.regs\[18\]\[25\] _03026_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__mux2_1
XANTENNA__13803__B1 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12918__A _06183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18332_ clknet_leaf_36_clk _01400_ VGND VGND VPWR VPWR mem_16bit_buffer\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15544_ cpuregs.regs\[8\]\[26\] cpuregs.regs\[9\]\[26\] cpuregs.regs\[10\]\[26\]
+ cpuregs.regs\[11\]\[26\] _03640_ _03642_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__mux4_1
XANTENNA__09499__A _04052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12756_ _06874_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11290__A0 reg_next_pc\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11707_ reg_pc\[21\] reg_pc\[20\] _06242_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__and3_1
X_18263_ clknet_leaf_26_clk _01334_ VGND VGND VPWR VPWR decoded_imm\[21\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_127_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12129__S _06518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15475_ _01969_ _02304_ _02312_ _02027_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__o211a_4
XFILLER_0_25_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12687_ _06835_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17214_ clknet_leaf_167_clk _00388_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14426_ decoded_imm_j\[10\] _07928_ VGND VGND VPWR VPWR _08094_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_170_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11260__C _05885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11638_ _03409_ _03352_ _06066_ _06198_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__a22o_1
X_18194_ clknet_leaf_28_clk _01265_ VGND VGND VPWR VPWR instr_lhu sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11968__S _06435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17145_ clknet_leaf_15_clk _00319_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_986 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14357_ _07986_ _08029_ _08030_ _07994_ _07915_ VGND VGND VPWR VPWR _08031_ sky130_fd_sc_hd__a32o_1
XFILLER_0_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11569_ reg_pc\[6\] reg_pc\[5\] _06121_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__and3_1
XANTENNA__15403__S0 _03661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09438__S _04064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13308_ _06995_ cpuregs.regs\[5\]\[25\] _07176_ VGND VGND VPWR VPWR _07182_ sky130_fd_sc_hd__mux2_1
X_17076_ clknet_leaf_112_clk _00250_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_14288_ _05941_ _06325_ _07944_ _05947_ VGND VGND VPWR VPWR _07968_ sky130_fd_sc_hd__o211a_2
XPHY_EDGE_ROW_139_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15964__A net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16027_ _02715_ decoded_imm_j\[4\] _02716_ mem_rdata_q\[11\] _02633_ VGND VGND VPWR
+ VPWR _02724_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13239_ _07145_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12799__S _06891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08780_ _03526_ _03544_ _03545_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__o21ai_2
X_17978_ clknet_leaf_44_clk _01115_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16929_ clknet_leaf_130_clk _00110_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16036__B2 mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10112__S _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14047__B1 _07790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_148_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09401_ _00071_ _04134_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09332_ _04054_ _04066_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11281__A0 _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09202__A _03767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09263_ mem_rdata_q\[30\] _04000_ _03757_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09194_ _03799_ _03926_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14762__B _08350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11878__S _06387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_157_Left_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13378__B decoded_imm\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15085__S _03713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14286__B1 _07944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08488__A _03239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08978_ mem_rdata_q\[14\] net38 _03208_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__mux2_1
XANTENNA__09388__S0 _04072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_166_Left_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16027__B2 mem_rdata_q\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10940_ _05361_ _05616_ _05626_ VGND VGND VPWR VPWR alu_out\[17\] sky130_fd_sc_hd__a21o_1
XFILLER_0_168_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10957__S _05517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10871_ _05561_ _05483_ _05295_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12738__A _06186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12610_ _06794_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15114__A _01968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13590_ _07281_ _07441_ _07305_ reg_pc\[15\] VGND VGND VPWR VPWR _07442_ sky130_fd_sc_hd__a22o_1
XANTENNA__11272__A0 _04754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12541_ cpuregs.regs\[2\]\[5\] _06544_ _06752_ VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__mux2_1
XANTENNA__16644__S _03051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15260_ _03664_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_152_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12472_ _06132_ cpuregs.regs\[28\]\[5\] _06715_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14211_ reg_pc\[4\] _07906_ _07915_ _07912_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11423_ _03412_ irq_mask\[1\] irq_pending\[1\] VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__or3b_1
XFILLER_0_34_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15191_ cpuregs.regs\[12\]\[7\] cpuregs.regs\[13\]\[7\] cpuregs.regs\[14\]\[7\] cpuregs.regs\[15\]\[7\]
+ _01936_ _03647_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08670__B net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 _02166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14142_ count_instr\[48\] _07862_ _07834_ VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11354_ _03215_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_130_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10305_ _04990_ _05012_ _05015_ _04007_ irq_pending\[25\] VGND VGND VPWR VPWR _08386_
+ sky130_fd_sc_hd__o32a_1
XANTENNA__15784__A _03630_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14073_ _07817_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__clkbuf_1
X_11285_ reg_out\[21\] _05909_ _05910_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12524__A0 _06336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10236_ _04391_ _04920_ _04921_ _04948_ VGND VGND VPWR VPWR _08384_ sky130_fd_sc_hd__a31o_1
X_17901_ clknet_leaf_94_clk _01070_ VGND VGND VPWR VPWR count_cycle\[46\] sky130_fd_sc_hd__dfxtp_1
X_13024_ _07031_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_167_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17832_ clknet_leaf_57_clk _01001_ VGND VGND VPWR VPWR reg_next_pc\[9\] sky130_fd_sc_hd__dfxtp_1
X_10167_ _03637_ _04880_ _04673_ _04881_ _04048_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__a221o_1
XANTENNA__09940__B2 _04023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15474__C1 _02006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17763_ clknet_leaf_90_clk _00932_ VGND VGND VPWR VPWR count_instr\[34\] sky130_fd_sc_hd__dfxtp_1
X_10098_ _04391_ _04786_ _04814_ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__a21o_1
XANTENNA__15008__B _01885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14975_ irq_mask\[0\] _01864_ _01866_ _08335_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__a211o_1
XANTENNA__10440__B decoded_imm\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16819__S _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16018__A1 decoded_imm\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_145_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16714_ _06980_ cpuregs.regs\[19\]\[18\] _03087_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13926_ _07714_ _07715_ VGND VGND VPWR VPWR _07716_ sky130_fd_sc_hd__and2_1
XANTENNA__09006__B _03747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17694_ clknet_leaf_162_clk _00863_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15226__C1 _02006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16645_ _03059_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15777__B1 _02486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13857_ cpuregs.regs\[0\]\[25\] VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11552__A reg_pc\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13788__C1 _03275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12808_ _06901_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__clkbuf_1
X_16576_ _06978_ cpuregs.regs\[18\]\[17\] _03015_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13788_ _07609_ _07623_ _07625_ _03275_ VGND VGND VPWR VPWR _07626_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09022__A _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18315_ clknet_leaf_36_clk _01383_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dfxtp_1
XANTENNA__11271__B _05899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15527_ _02360_ _02361_ _01907_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12739_ decoded_rd\[0\] _06863_ _06864_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09471__A3 _04203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15624__S0 _03640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18246_ clknet_leaf_25_clk _01317_ VGND VGND VPWR VPWR decoded_imm\[4\] sky130_fd_sc_hd__dfxtp_2
X_15458_ _02291_ _02293_ _02296_ _03683_ _02004_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14409_ reg_next_pc\[8\] _07947_ _08077_ _08078_ VGND VGND VPWR VPWR _08079_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18177_ clknet_leaf_31_clk _01248_ VGND VGND VPWR VPWR decoded_imm_j\[18\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15389_ _02220_ _02225_ _02228_ _02231_ _01968_ _02037_ VGND VGND VPWR VPWR _02232_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__10369__A2 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17128_ clknet_leaf_134_clk _00302_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09950_ _04666_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__inv_2
X_17059_ clknet_leaf_142_clk _00233_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08901_ _00066_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_4_9_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09881_ _04420_ _04603_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_55_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16257__A1 _03895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08832_ _03434_ _03438_ _03594_ _03597_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__a31o_1
X_08763_ _03527_ _03528_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__nand2b_2
XANTENNA__16729__S _03098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10829__B1 _05301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08694_ net82 VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__inv_2
XANTENNA__13491__A1 _04419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09695__B1 _04422_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13153__S _07093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09315_ irq_pending\[0\] _04008_ _04029_ _04050_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__o22a_1
XANTENNA__10057__B2 _04231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12992__S _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15615__S0 _01995_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10152__S1 _04284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09246_ _03976_ _03978_ _03986_ _03888_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08771__A net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15091__S1 _03646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09177_ _03770_ _03926_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__nor2_2
XANTENNA__15940__B1 _02659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11101__S0 _05324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12506__A0 _06266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11070_ _05689_ _05243_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__or2b_1
Xoutput68 net68 VGND VGND VPWR VPWR cpi_rs1[10] sky130_fd_sc_hd__clkbuf_1
Xoutput79 net79 VGND VGND VPWR VPWR cpi_rs1[20] sky130_fd_sc_hd__buf_1
X_10021_ _04168_ _04738_ _04739_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__a21o_1
XANTENNA__18130__D alu_out\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ count_cycle\[22\] count_cycle\[23\] _01722_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__and3_1
XANTENNA__13482__A1 _07274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11972_ _06193_ cpuregs.regs\[21\]\[12\] _06435_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__mux2_1
XANTENNA__08946__A _03666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13711_ _07508_ _07548_ _07553_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10923_ _03485_ _05609_ _05610_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14691_ count_cycle\[0\] count_cycle\[1\] _07675_ VGND VGND VPWR VPWR _08336_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16430_ _06968_ cpuregs.regs\[29\]\[12\] _02943_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__mux2_1
XANTENNA__10391__S1 _04283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13642_ _07488_ _07489_ VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_123_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10854_ _05414_ _05404_ _05545_ _05250_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16361_ _02909_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__clkbuf_1
X_13573_ _04466_ _07315_ _07425_ _07216_ VGND VGND VPWR VPWR _07426_ sky130_fd_sc_hd__o211a_1
XANTENNA__16374__S _02907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10785_ _05249_ _05480_ _05288_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10599__A2 _05301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18100_ clknet_leaf_90_clk _01204_ VGND VGND VPWR VPWR timer\[15\] sky130_fd_sc_hd__dfxtp_1
X_15312_ _02012_ _02158_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__or2_1
X_12524_ _06336_ cpuregs.regs\[28\]\[30\] _06714_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ _02872_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08681__A net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18031_ clknet_leaf_66_clk _00007_ VGND VGND VPWR VPWR irq_pending\[15\] sky130_fd_sc_hd__dfxtp_1
X_15243_ cpuregs.regs\[16\]\[9\] cpuregs.regs\[17\]\[9\] cpuregs.regs\[18\]\[9\] cpuregs.regs\[19\]\[9\]
+ _01999_ _02000_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12455_ cpuregs.regs\[27\]\[30\] _06596_ _06677_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12407__S _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11406_ _05960_ _03910_ _06003_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_169_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15174_ cpuregs.regs\[4\]\[6\] cpuregs.regs\[5\]\[6\] cpuregs.regs\[6\]\[6\] cpuregs.regs\[7\]\[6\]
+ _02013_ _02014_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12386_ cpuregs.regs\[26\]\[30\] _06596_ _06640_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14125_ _07852_ _07853_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__nor2_1
X_11337_ _05946_ _05948_ _05952_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output77_A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14056_ count_instr\[22\] _07803_ _07790_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__o21ai_1
X_11268_ _05838_ _05895_ _05896_ _05897_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__o31ai_4
XFILLER_0_120_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09913__A1 _04017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09374__C1 _03303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13007_ cpuregs.regs\[3\]\[11\] _06557_ _07021_ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__mux2_1
XANTENNA__13238__S _07140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15019__A _04805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10219_ cpuregs.regs\[24\]\[23\] cpuregs.regs\[25\]\[23\] cpuregs.regs\[26\]\[23\]
+ cpuregs.regs\[27\]\[23\] _04281_ _04470_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__mux4_1
X_11199_ _05836_ _05840_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11720__A1 _06252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09017__A _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11266__B _05894_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17815_ clknet_leaf_63_clk _00984_ VGND VGND VPWR VPWR reg_pc\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15998__B1 _03892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10170__B decoded_imm\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16549__S _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17746_ clknet_leaf_86_clk _00915_ VGND VGND VPWR VPWR count_instr\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14958_ _01854_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13473__A1 _07217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13909_ _07703_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11484__B1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17677_ clknet_leaf_136_clk _00846_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14889_ _07633_ _07636_ _01813_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__nor3_1
XFILLER_0_89_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10382__S1 _04376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16628_ _03050_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10039__B2 _04165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16559_ _06961_ cpuregs.regs\[18\]\[9\] _03004_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__mux2_1
XANTENNA__16284__S _02859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09100_ _03785_ _03788_ _03845_ _03859_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__or4_1
XANTENNA__09687__A _04414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09031_ _03791_ _03792_ _03231_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__mux2_1
X_18229_ clknet_leaf_23_clk _01300_ VGND VGND VPWR VPWR decoded_rd\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15922__B1 _02620_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12317__S _06603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12736__B1 _06861_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15686__C1 _06026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09933_ cpuregs.regs\[12\]\[15\] cpuregs.regs\[13\]\[15\] cpuregs.regs\[14\]\[15\]
+ cpuregs.regs\[15\]\[15\] _04487_ _04469_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10361__A _04051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12052__S _06471_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09864_ cpuregs.regs\[12\]\[13\] cpuregs.regs\[13\]\[13\] cpuregs.regs\[14\]\[13\]
+ cpuregs.regs\[15\]\[13\] _04280_ _04059_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__mux4_1
XANTENNA__11711__A1 _06252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08815_ net114 _03460_ _03474_ _03572_ _03580_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__o221a_1
XANTENNA__08469__C instr_rdcycleh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15989__B1 _06016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09795_ _04518_ _04519_ _04287_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__mux2_1
XANTENNA__16459__S _02954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08746_ _03509_ _03511_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__nand2_2
XANTENNA__09668__B1 _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08766__A net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09763__S0 _04487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08677_ net120 net88 VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13767__A2 decoded_imm\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11778__A1 reg_pc\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10570_ net87 net88 _05263_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12735__B _06860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15064__S1 _03671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16207__B _07898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09229_ _03779_ _03784_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__nor2_1
XANTENNA__15913__B1 _02650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12227__S _06576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10536__A _05239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12240_ _06593_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09199__A2 _03810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10202__B2 _04915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12171_ cpuregs.regs\[24\]\[6\] _06546_ _06534_ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__mux2_1
XANTENNA__15538__S _03653_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15765__C _02560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11122_ _05361_ _05788_ _05795_ VGND VGND VPWR VPWR alu_out\[30\] sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_147_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13566__B decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13058__S _07046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11053_ _05683_ _05243_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__or2b_1
X_15930_ is_alu_reg_imm _02625_ _02654_ _02655_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__and4_1
X_10004_ _04721_ _04722_ _04065_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09371__A2 _04104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15861_ _03940_ _02619_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__nor2_2
XANTENNA__12897__S _06943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ clknet_leaf_169_clk _00769_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15444__A2 _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14812_ count_cycle\[37\] count_cycle\[38\] count_cycle\[39\] _01756_ VGND VGND VPWR
+ VPWR _01762_ sky130_fd_sc_hd__and4_2
X_18580_ clknet_leaf_174_clk _01645_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15792_ _04156_ _06863_ _03368_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__and3_1
XANTENNA__10269__A1 instr_retirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17531_ clknet_leaf_166_clk _00700_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11466__B1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14743_ _03239_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__buf_4
XANTENNA__09754__S0 _04085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11955_ _06125_ cpuregs.regs\[21\]\[4\] _06424_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__mux2_1
XANTENNA_output115_A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12198__A _06215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10906_ _05588_ _05592_ _05594_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__or3b_1
X_17462_ clknet_leaf_97_clk _00631_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14674_ _07968_ _07969_ _08301_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__and3_1
X_11886_ _06125_ cpuregs.regs\[20\]\[4\] _06387_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_103_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16413_ _06951_ cpuregs.regs\[29\]\[4\] _02932_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__mux2_1
X_13625_ _07472_ _07473_ VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__nand2_1
XANTENNA__14955__A1 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10837_ _03530_ _05384_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__nor2_1
X_17393_ clknet_leaf_141_clk _00562_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11769__A1 reg_pc\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16344_ _02900_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__clkbuf_1
X_13556_ _07408_ _07409_ VGND VGND VPWR VPWR _07410_ sky130_fd_sc_hd__xnor2_1
X_10768_ _05255_ _05261_ _05458_ _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__a31o_1
XANTENNA__09300__A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15055__S1 _03659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12507_ _06739_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16275_ _02863_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12137__S _06518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13487_ _03510_ decoded_imm\[8\] VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10699_ _05226_ _05210_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__nor2_2
XFILLER_0_54_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18014_ clknet_leaf_77_clk _01151_ VGND VGND VPWR VPWR irq_mask\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15226_ _02068_ _02072_ _02077_ _02037_ _02006_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__a221o_1
X_12438_ _06702_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11976__S _06435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15157_ cpuregs.regs\[8\]\[6\] cpuregs.regs\[9\]\[6\] cpuregs.regs\[10\]\[6\] cpuregs.regs\[11\]\[6\]
+ _01970_ _01971_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12369_ _06665_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_112_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15668__C1 _06026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14108_ _07840_ _07815_ _07841_ VGND VGND VPWR VPWR _07842_ sky130_fd_sc_hd__and3b_1
XFILLER_0_121_983 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09446__S _04077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15088_ cpuregs.regs\[24\]\[1\] cpuregs.regs\[25\]\[1\] cpuregs.regs\[26\]\[1\] cpuregs.regs\[27\]\[1\]
+ _03669_ _03646_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__mux4_1
XFILLER_0_129_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11277__A _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15972__A mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14039_ count_instr\[17\] _07792_ _07675_ VGND VGND VPWR VPWR _07794_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13694__A1 _04810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10052__S0 _04472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13492__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08600_ _03377_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__buf_2
XANTENNA__16632__A1 _06183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09580_ _04268_ _04270_ _04310_ _03302_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08531_ cpu_state\[6\] cpu_state\[5\] VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__nor2_4
XANTENNA__09745__S0 _04281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17729_ clknet_leaf_101_clk _00898_ VGND VGND VPWR VPWR count_instr\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_121_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10355__S1 _04060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10120__S _04430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08462_ irq_mask\[2\] irq_active _03245_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15294__S1 _02070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1004 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09014_ _03762_ _03775_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__nand2_2
XANTENNA__11886__S _06387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10790__S _05244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09050__A1 mem_rdata_q\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09916_ _03638_ _04611_ _04613_ _03226_ _04637_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__a221o_1
XANTENNA__15882__A _02634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10499__A1 _04010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10043__S0 _04057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09847_ _04391_ _04539_ _04542_ _04570_ VGND VGND VPWR VPWR _08372_ sky130_fd_sc_hd__a31o_1
XANTENNA__11696__B1 _06093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15093__S _03713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16623__A1 _06149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12510__S _06737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09778_ _04462_ _04464_ _04461_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_87_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ net103 net71 VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__C1 _04188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _06289_ cpuregs.regs\[10\]\[24\] _06258_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11671_ reg_pc\[17\] _06218_ _06227_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13410_ _07272_ _07236_ VGND VGND VPWR VPWR _07273_ sky130_fd_sc_hd__nand2_1
XANTENNA__15122__A _01919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10622_ _05323_ _05324_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14390_ decoded_imm_j\[7\] _07921_ VGND VGND VPWR VPWR _08061_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13341_ _07195_ _07199_ _04227_ _07207_ VGND VGND VPWR VPWR _07208_ sky130_fd_sc_hd__a211o_4
X_10553_ _05256_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__buf_2
XFILLER_0_51_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16060_ _03402_ decoded_imm_j\[18\] _03403_ mem_rdata_q\[18\] VGND VGND VPWR VPWR
+ _02743_ sky130_fd_sc_hd__a22o_1
X_13272_ _06959_ cpuregs.regs\[5\]\[8\] _07154_ VGND VGND VPWR VPWR _07163_ sky130_fd_sc_hd__mux2_1
XANTENNA__15362__A1 _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10484_ cpuregs.regs\[24\]\[31\] cpuregs.regs\[25\]\[31\] cpuregs.regs\[26\]\[31\]
+ cpuregs.regs\[27\]\[31\] _04274_ _04317_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__mux4_1
X_15011_ irq_mask\[15\] _01880_ _01887_ _01876_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12223_ _06280_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__buf_2
XFILLER_0_122_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12154_ _06535_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10282__S0 _04275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11105_ _05600_ _05668_ _05778_ _03443_ _05779_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__a221o_1
XANTENNA__15792__A _04156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12085_ _06096_ cpuregs.regs\[23\]\[1\] _06496_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__mux2_1
X_16962_ clknet_leaf_182_clk _00136_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_11036_ _05287_ _05399_ _05714_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__and3_1
X_15913_ is_alu_reg_imm _02625_ _02649_ _02650_ instr_srli VGND VGND VPWR VPWR _01276_
+ sky130_fd_sc_hd__a32o_1
XANTENNA__09975__S0 _04232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output232_A net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16893_ clknet_leaf_35_clk _00038_ VGND VGND VPWR VPWR mem_rdata_q\[12\] sky130_fd_sc_hd__dfxtp_1
X_18632_ clknet_leaf_149_clk _01692_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_15844_ instr_auipc _02605_ _03635_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__mux2_1
XANTENNA__12420__S _06689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14201__A _07901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13979__A2 _07677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15775_ _05170_ _02486_ _02568_ _02545_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__o211a_1
XANTENNA__15016__B _01885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18563_ clknet_leaf_145_clk _01628_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12987_ _07012_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16827__S _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14726_ count_cycle\[12\] _08356_ _07877_ VGND VGND VPWR VPWR _08360_ sky130_fd_sc_hd__o21ai_1
X_17514_ clknet_leaf_175_clk _00683_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18494_ clknet_leaf_182_clk _01559_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_11938_ _06328_ cpuregs.regs\[20\]\[29\] _06409_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14855__B _01753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15276__S1 _01986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17445_ clknet_leaf_2_clk _00614_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14657_ _08272_ _08280_ _08287_ _08295_ VGND VGND VPWR VPWR _08306_ sky130_fd_sc_hd__or4_1
X_11869_ _06336_ cpuregs.regs\[11\]\[30\] _06347_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__mux2_1
X_13608_ _07458_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17376_ clknet_leaf_21_clk _00545_ VGND VGND VPWR VPWR cpuregs.waddr\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_172_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09804__B1 instr_rdcycleh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14588_ _08226_ _08231_ _08242_ VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_45_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_984 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10414__A1 _04018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16327_ _02890_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13539_ _07345_ _07346_ _07352_ _07393_ VGND VGND VPWR VPWR _07394_ sky130_fd_sc_hd__or4bb_1
XANTENNA__16562__S _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15353__A1 decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16258_ _02853_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_934 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput203 net203 VGND VGND VPWR VPWR mem_la_addr[19] sky130_fd_sc_hd__clkbuf_1
XANTENNA__13487__A _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15209_ cpuregs.regs\[20\]\[8\] cpuregs.regs\[21\]\[8\] cpuregs.regs\[22\]\[8\] cpuregs.regs\[23\]\[8\]
+ _01970_ _01971_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__mux4_1
Xoutput214 net214 VGND VGND VPWR VPWR mem_la_addr[2] sky130_fd_sc_hd__buf_1
X_16189_ _03221_ _01821_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput225 net225 VGND VGND VPWR VPWR mem_la_wdata[0] sky130_fd_sc_hd__buf_1
XFILLER_0_3_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput236 net236 VGND VGND VPWR VPWR mem_la_wdata[1] sky130_fd_sc_hd__buf_1
XANTENNA__10717__A2 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput247 net247 VGND VGND VPWR VPWR mem_la_wdata[2] sky130_fd_sc_hd__clkbuf_1
XANTENNA__15105__A1 _05413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput258 net258 VGND VGND VPWR VPWR mem_la_wstrb[0] sky130_fd_sc_hd__buf_1
XANTENNA__13116__A0 _07007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput269 net269 VGND VGND VPWR VPWR mem_wdata[15] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14313__C1 _06860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09701_ count_instr\[9\] _04145_ _04018_ count_cycle\[41\] VGND VGND VPWR VPWR _04428_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09966__S0 _04579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11142__A2 _05413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15408__A2 _02241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09632_ net57 _03242_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__or2b_1
XANTENNA__12330__S _06641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09563_ cpuregs.regs\[0\]\[5\] cpuregs.regs\[1\]\[5\] cpuregs.regs\[2\]\[5\] cpuregs.regs\[3\]\[5\]
+ _04291_ _04292_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__mux4_1
XANTENNA__08797__A_N net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16737__S _03098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08514_ mem_do_wdata net66 _03220_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__and3_1
XFILLER_0_172_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_162_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09494_ _04215_ _04224_ _04225_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08445_ _03199_ mem_do_prefetch VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__nor2_2
XFILLER_0_59_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10785__S _05288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09859__B _04581_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11470__A _06053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_984 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11602__A0 _06166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_177_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16541__A0 _06941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13355__B1 _05211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15895__A2 _02611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10708__A2 _05261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xalphacore_309 VGND VGND VPWR VPWR alphacore_309/HI cpi_insn[7] sky130_fd_sc_hd__conb_1
XFILLER_0_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12330__A1 _06540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12910_ _06960_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__clkbuf_1
X_13890_ _07690_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14607__B1 _07959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10892__A1 _05225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12841_ _06193_ cpuregs.regs\[6\]\[12\] _06917_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__mux2_1
XANTENNA__09709__S0 _04274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15942__B_N mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10319__S1 _04073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ cpuregs.regs\[12\]\[27\] cpuregs.regs\[13\]\[27\] cpuregs.regs\[14\]\[27\]
+ cpuregs.regs\[15\]\[27\] _01999_ _02000_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__mux4_1
XFILLER_0_150_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12772_ cpuregs.regs\[9\]\[12\] _06559_ _06880_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14511_ _08150_ _08166_ VGND VGND VPWR VPWR _08172_ sky130_fd_sc_hd__or2_1
XANTENNA__10644__A1 _04532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15258__S1 _01992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11723_ _06274_ cpuregs.regs\[10\]\[22\] _06258_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08932__S1 _03684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15491_ _02326_ _02327_ _03713_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17230_ clknet_leaf_123_clk _00404_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14442_ _08106_ _08108_ _03368_ VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11654_ reg_out\[15\] alu_out_q\[15\] _06067_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_973 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10605_ net82 net83 _05263_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17161_ clknet_leaf_134_clk _00335_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14373_ reg_next_pc\[5\] _07947_ _08045_ _08033_ VGND VGND VPWR VPWR _08046_ sky130_fd_sc_hd__a22o_1
X_11585_ _06151_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16112_ _03221_ _02676_ _02771_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_24_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13324_ _07190_ VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10536_ _05239_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15335__A1 _01969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17092_ clknet_leaf_157_clk _00266_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output182_A net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13346__B1 _03311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15886__A2 _02635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15430__S1 _01980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16043_ decoded_imm\[10\] _02711_ _02733_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__o21a_1
X_13255_ _07153_ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10467_ _04268_ _05152_ _05172_ _03302_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12206_ _06570_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10255__S0 _04290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13186_ _06383_ _06084_ VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__nand2_2
XFILLER_0_20_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10398_ _05093_ _05097_ net301 _05105_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__a211o_2
XFILLER_0_103_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12137_ _06304_ cpuregs.regs\[23\]\[26\] _06518_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__mux2_1
XANTENNA__13649__A1 _04708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17994_ clknet_leaf_103_clk _01131_ VGND VGND VPWR VPWR irq_mask\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10007__S0 _04072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16945_ clknet_leaf_169_clk _00126_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_12068_ _06488_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08848__B _03518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09722__C1 _04027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11555__A _06124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13246__S _07140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11019_ _05458_ _05597_ _05694_ _05699_ VGND VGND VPWR VPWR alu_out\[23\] sky130_fd_sc_hd__a211o_1
XANTENNA__15027__A _04940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16876_ _03182_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16063__A2 _02611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15497__S1 _01971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09025__A _03213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18615_ clknet_leaf_9_clk _00089_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__dfxtp_2
X_15827_ decoded_imm_j\[14\] _05987_ _03891_ _02587_ _02596_ VGND VGND VPWR VPWR _01244_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16557__S _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13770__A net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15758_ _05037_ _02479_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18546_ clknet_leaf_117_clk _01611_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14585__B _07958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10096__C1 _04202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11832__A0 _06193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14709_ count_cycle\[7\] _08346_ _07826_ VGND VGND VPWR VPWR _08348_ sky130_fd_sc_hd__a21oi_1
X_15689_ timer\[8\] _02500_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__nor2_1
X_18477_ clknet_leaf_161_clk _01542_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15023__B1 _01714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17428_ clknet_leaf_179_clk _00597_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12388__A1 _06598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17359_ clknet_leaf_139_clk _00528_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09253__A1 _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10938__A2 _05301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13888__A1 _03344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10020__C1 _04027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15629__A2 _02449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10571__A0 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08994_ _03752_ _03754_ _03755_ _03753_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09615_ net61 net258 _04035_ net47 _04344_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__a221o_2
XANTENNA__16054__A2 decoded_imm_j\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16467__S _02931_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13680__A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09546_ _04276_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10626__A1 _05281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09477_ cpuregs.regs\[28\]\[4\] cpuregs.regs\[29\]\[4\] cpuregs.regs\[30\]\[4\] cpuregs.regs\[31\]\[4\]
+ _04207_ _04208_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_80_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12296__A _06603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08428_ _03206_ _03213_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__and2_1
XANTENNA__15565__A1 decoded_imm\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11350__D _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11051__A1 _05013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11370_ cpuregs.raddr2\[2\] _05974_ _05980_ _05982_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__a22o_1
XANTENNA__08812__A_N net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15412__S1 _03671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10321_ _05029_ _05030_ _00071_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__mux2_1
XANTENNA__18133__D alu_out\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13879__A1 _03338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10544__A _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14016__A _03304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13040_ cpuregs.regs\[3\]\[27\] _06590_ _07032_ VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__mux2_1
X_10252_ cpuregs.regs\[8\]\[24\] cpuregs.regs\[9\]\[24\] cpuregs.regs\[10\]\[24\]
+ cpuregs.regs\[11\]\[24\] _04216_ _04376_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__mux4_1
X_10183_ _04895_ _04896_ _04065_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__mux2_1
X_14991_ _03240_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13066__S _07046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12303__A1 _06582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13942_ _07726_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16730_ _03104_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16045__A2 decoded_imm_j\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16661_ cpuregs.regs\[1\]\[25\] _06296_ _03062_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__mux2_1
X_13873_ _03301_ _07676_ VGND VGND VPWR VPWR _07677_ sky130_fd_sc_hd__nor2_2
X_15612_ net122 _01906_ _02441_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__o21a_1
X_18400_ clknet_leaf_159_clk _01465_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12824_ _06125_ cpuregs.regs\[6\]\[4\] _06906_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__mux2_1
X_16592_ _03031_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08684__A net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13803__A1 _07304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15543_ cpuregs.regs\[12\]\[26\] cpuregs.regs\[13\]\[26\] cpuregs.regs\[14\]\[26\]
+ cpuregs.regs\[15\]\[26\] _03661_ _03642_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__mux4_1
X_18331_ clknet_leaf_36_clk _01399_ VGND VGND VPWR VPWR mem_16bit_buffer\[2\] sky130_fd_sc_hd__dfxtp_1
X_12755_ cpuregs.regs\[9\]\[4\] _06542_ _06869_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11706_ _06259_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__clkbuf_1
X_18262_ clknet_leaf_26_clk _01333_ VGND VGND VPWR VPWR decoded_imm\[20\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_166_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16753__A0 _06536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15474_ _02306_ _02308_ _02311_ _02004_ _02006_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__a221o_1
X_12686_ _06166_ cpuregs.regs\[12\]\[9\] _06825_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17213_ clknet_leaf_2_clk _00387_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_14425_ _07925_ _08076_ _07928_ VGND VGND VPWR VPWR _08093_ sky130_fd_sc_hd__a21oi_1
X_11637_ reg_out\[13\] alu_out_q\[13\] _06068_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18193_ clknet_leaf_40_clk _01264_ VGND VGND VPWR VPWR instr_lbu sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11260__D _05889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17144_ clknet_leaf_176_clk _00318_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14356_ _07915_ _08016_ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__or2_1
X_11568_ _06116_ reg_next_pc\[6\] _06135_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15403__S1 _03662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13307_ _07181_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__clkbuf_1
X_10519_ _03610_ _05221_ _05222_ _03611_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_122_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17075_ clknet_leaf_19_clk _00249_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_14287_ reg_pc\[28\] _07953_ _07967_ _07960_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__a22o_1
XANTENNA__16840__S _03163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11499_ _06071_ latched_compr _03338_ _06072_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16026_ mem_rdata_q\[24\] _02712_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__and2_1
XANTENNA__09538__A2 _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13238_ _06993_ cpuregs.regs\[8\]\[24\] _07140_ VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__mux2_1
XANTENNA__11984__S _06435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09962__B decoded_imm\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15167__S0 _01990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13169_ _07108_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17977_ clknet_leaf_44_clk _01114_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_137_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15492__B1 _03657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16928_ clknet_leaf_145_clk _00109_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16036__A2 decoded_imm_j\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16859_ _03173_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14596__A _03293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09400_ cpuregs.regs\[0\]\[2\] cpuregs.regs\[1\]\[2\] cpuregs.regs\[2\]\[2\] cpuregs.regs\[3\]\[2\]
+ _04123_ _04124_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15795__A1 _03292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08594__A _03196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09331_ _04061_ _04062_ _04065_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__mux2_1
X_18529_ clknet_leaf_157_clk _01594_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_5_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15547__A1 _03639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09262_ _03753_ _03740_ _03741_ _03850_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__a22o_2
XFILLER_0_146_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09193_ _03940_ _03891_ _03757_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10219__S0 _04281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11336__A2 _05948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12533__A1 _06536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11894__S _06387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08769__A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08977_ _03213_ _03206_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__nor2b_4
XTAP_TAPCELL_ROW_90_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11195__A _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15890__A is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09388__S1 _04074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09701__A2 _04145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10870_ net71 net70 net69 net68 _05264_ _05235_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12738__B _06863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09529_ _04258_ _04259_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18128__D alu_out\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12540_ _06757_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13549__A0 _04566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12471_ _06720_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14210_ _07914_ VGND VGND VPWR VPWR _07915_ sky130_fd_sc_hd__buf_2
XFILLER_0_136_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11422_ irq_pending\[1\] _03308_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__or2_1
XANTENNA__15130__A _01936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15190_ _02041_ _02042_ _03664_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__mux2_1
XANTENNA__10458__S0 _04487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_1013 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14141_ _07864_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__clkbuf_2
X_11353_ _05960_ _03864_ _05967_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__and3_1
XANTENNA__10783__A0 _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10274__A reg_pc\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15397__S0 _02046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10304_ _03680_ _05013_ _04752_ _05014_ _04202_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__a221o_1
X_14072_ _07814_ _07815_ _07816_ VGND VGND VPWR VPWR _07817_ sky130_fd_sc_hd__and3b_1
X_11284_ reg_next_pc\[21\] _05898_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17900_ clknet_leaf_94_clk _01069_ VGND VGND VPWR VPWR count_cycle\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13023_ cpuregs.regs\[3\]\[19\] _06573_ _07021_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__mux2_1
X_10235_ irq_pending\[23\] _04006_ _04944_ _04947_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17831_ clknet_leaf_58_clk _01000_ VGND VGND VPWR VPWR reg_next_pc\[8\] sky130_fd_sc_hd__dfxtp_1
X_10166_ net46 _04745_ _04666_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__a21o_1
XANTENNA__09940__A2 _04021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11309__S _03219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17762_ clknet_leaf_90_clk _00931_ VGND VGND VPWR VPWR count_instr\[33\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10213__S _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10097_ irq_pending\[19\] _04007_ _04809_ _04813_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__o22a_1
X_14974_ _07208_ _01865_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_128_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10299__C1 _04188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16018__A2 _02711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16713_ _03095_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__clkbuf_1
X_13925_ _03353_ _07704_ _07705_ net136 VGND VGND VPWR VPWR _07715_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_145_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17693_ clknet_leaf_125_clk _00862_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15305__A _01989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16644_ cpuregs.regs\[1\]\[17\] _06231_ _03051_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__mux2_1
X_13856_ _07667_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12807_ cpuregs.regs\[9\]\[29\] _06594_ _06891_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13787_ _07624_ _07611_ _07622_ VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16575_ _03022_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16835__S _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10999_ _05679_ _05680_ _05218_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09456__B2 _04187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18314_ clknet_leaf_36_clk _01382_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15526_ cpuregs.regs\[24\]\[25\] cpuregs.regs\[25\]\[25\] cpuregs.regs\[26\]\[25\]
+ cpuregs.regs\[27\]\[25\] _02074_ _02075_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__mux4_1
XANTENNA__09022__B _03213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15529__A1 _01969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12738_ _06186_ _06863_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_167_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15624__S1 _03642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15457_ _02294_ _02295_ _01907_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__mux2_1
X_18245_ clknet_leaf_25_clk _01316_ VGND VGND VPWR VPWR decoded_imm\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_170_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12669_ _06826_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11015__A1 _05323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09449__S _04063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14408_ _03378_ _07921_ _08048_ _07924_ _03293_ VGND VGND VPWR VPWR _08078_ sky130_fd_sc_hd__a32o_1
XFILLER_0_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15388_ _02229_ _02230_ _02110_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__mux2_1
X_18176_ clknet_leaf_31_clk _01247_ VGND VGND VPWR VPWR decoded_imm_j\[17\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17127_ clknet_leaf_142_clk _00301_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14339_ _07998_ _08004_ VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__or2_1
XANTENNA__16570__S _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10184__A _04054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17058_ clknet_leaf_183_clk _00232_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15701__A1 _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08900_ _03660_ _03663_ _03664_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__mux2_1
X_16009_ cpuregs.raddr2\[4\] _06006_ _05986_ _05988_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__o22a_1
XANTENNA__09916__C1 _04637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09880_ net54 _04030_ _04034_ net37 _04423_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__o221a_1
XANTENNA__09692__B _04363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12603__S _06788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10912__A _05244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _03434_ _03595_ _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08762_ net125 net93 VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__nand2_1
XANTENNA__10123__S _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13476__C1 _07221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15560__S0 _01999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08693_ _03457_ _03458_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__nor2_1
XANTENNA__13491__A2 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15768__A1 _05107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09213__A _03935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09314_ _03226_ _04043_ _04047_ _04049_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__a211o_2
XFILLER_0_75_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09998__A2 decoded_imm\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15615__S1 _01937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09245_ _03879_ _03867_ _03923_ _03983_ _03985_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__a311o_1
XFILLER_0_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11006__A1 _05281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09359__S _04064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09176_ _03736_ _03925_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__nor2_1
XANTENNA__15940__B2 _02665_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11101__S1 _05286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15885__A _02611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10094__A _04668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10765__B1 _05215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15153__C1 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13703__B1 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput69 net69 VGND VGND VPWR VPWR cpi_rs1[11] sky130_fd_sc_hd__buf_1
XANTENNA__08499__A _03218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10020_ irq_mask\[17\] _04448_ timer\[17\] _04187_ _04027_ VGND VGND VPWR VPWR _04739_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15551__S0 _01979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ _06437_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13710_ _07526_ _07549_ _07551_ _07552_ _07542_ VGND VGND VPWR VPWR _07553_ sky130_fd_sc_hd__o311a_1
X_10922_ _03485_ _05609_ _05218_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15125__A _01919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15303__S0 _01970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14690_ _08335_ count_cycle\[0\] VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13641_ net77 decoded_imm\[19\] VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_123_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10853_ _05292_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_123_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16655__S _03062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14431__A1 _08035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14964__A _07737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16360_ _06966_ cpuregs.regs\[16\]\[11\] _02907_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__mux2_1
XANTENNA__16708__A0 _06974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13572_ _04754_ _07276_ VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__or2_1
X_10784_ _05479_ _05441_ _05401_ _05342_ _05266_ _05395_ VGND VGND VPWR VPWR _05480_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15311_ cpuregs.regs\[20\]\[13\] cpuregs.regs\[21\]\[13\] cpuregs.regs\[22\]\[13\]
+ cpuregs.regs\[23\]\[13\] _01990_ _01992_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12523_ _06747_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16291_ _06966_ cpuregs.regs\[15\]\[11\] _02870_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__mux2_1
XANTENNA__09777__B decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08681__B net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18030_ clknet_leaf_66_clk _00006_ VGND VGND VPWR VPWR irq_pending\[14\] sky130_fd_sc_hd__dfxtp_1
X_15242_ _01989_ _02092_ _03654_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__o21a_1
X_12454_ _06710_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15931__B2 mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11405_ _03867_ _05994_ _06013_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15173_ _01959_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_169_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12385_ _06673_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14124_ count_instr\[43\] _07849_ _07834_ VGND VGND VPWR VPWR _07853_ sky130_fd_sc_hd__o21ai_1
X_11336_ _05946_ _05948_ _05952_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__a21oi_1
XANTENNA_output262_A net262 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14055_ count_instr\[22\] count_instr\[21\] count_instr\[20\] _07799_ VGND VGND VPWR
+ VPWR _07805_ sky130_fd_sc_hd__and4_2
X_11267_ _04744_ _05838_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13006_ _07022_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10218_ _04483_ _04930_ _04296_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15019__B _01885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11198_ reg_next_pc\[5\] reg_out\[5\] _05834_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__mux2_2
XANTENNA__11720__A2 _03320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17814_ clknet_leaf_63_clk _00983_ VGND VGND VPWR VPWR reg_pc\[22\] sky130_fd_sc_hd__dfxtp_2
X_10149_ cpuregs.regs\[24\]\[21\] cpuregs.regs\[25\]\[21\] cpuregs.regs\[26\]\[21\]
+ cpuregs.regs\[27\]\[21\] _04758_ _04759_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__mux4_1
XANTENNA__15961__C _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17745_ clknet_leaf_87_clk _00914_ VGND VGND VPWR VPWR count_instr\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10878__S _05363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14957_ net213 net182 _01846_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__mux2_1
XANTENNA__09677__A1 _04070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11563__A _06131_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15035__A _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13908_ _07691_ _07702_ VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__and2_1
XANTENNA__11484__A1 _06054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17676_ clknet_leaf_150_clk _00845_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_14888_ _05205_ decoded_imm\[31\] VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__xor2_1
XFILLER_0_159_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16627_ cpuregs.regs\[1\]\[9\] _06165_ _03040_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__mux2_1
XANTENNA__09429__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13839_ cpuregs.regs\[0\]\[16\] VGND VGND VPWR VPWR _07659_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09429__B2 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14422__A1 _08012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10039__A2 _04012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16558_ _03013_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15509_ cpuregs.regs\[20\]\[24\] cpuregs.regs\[21\]\[24\] cpuregs.regs\[22\]\[24\]
+ cpuregs.regs\[23\]\[24\] _02022_ _02023_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16175__A1 net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16489_ cpuregs.regs\[17\]\[8\] _06550_ _02968_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09030_ net60 mem_rdata_q\[5\] _03729_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18228_ clknet_leaf_32_clk _01299_ VGND VGND VPWR VPWR decoded_rd\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12736__A1 _03309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18159_ clknet_leaf_21_clk _01230_ VGND VGND VPWR VPWR do_waitirq sky130_fd_sc_hd__dfxtp_1
XANTENNA__10747__B1 _05356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09932_ _04651_ _04652_ _04121_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _04320_ _04585_ _04068_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_70_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11172__B1 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10361__B _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08814_ _03469_ _03579_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__or2_1
XANTENNA__11711__A2 _03346_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09794_ cpuregs.regs\[24\]\[11\] cpuregs.regs\[25\]\[11\] cpuregs.regs\[26\]\[11\]
+ cpuregs.regs\[27\]\[11\] _04282_ _04285_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08745_ net129 _03510_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08766__B net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13164__S _07104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12672__A0 _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08676_ _03440_ _03441_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__and2b_1
XANTENNA__09763__S1 _04469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10089__A _04805_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16475__S _02968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10435__C1 _04150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09840__A1 _04271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12508__S _06737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09228_ _03749_ _03966_ _03969_ _03739_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__o211a_1
XANTENNA__16207__C _06863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15913__A1 is_alu_reg_imm VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09159_ _03912_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10202__A2 _04006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12170_ _06140_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__buf_2
XFILLER_0_101_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15677__B1 _02488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11121_ _05574_ _05621_ _05789_ _05794_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__a211o_1
XANTENNA__11648__A _06207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18141__D alu_out\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ _05729_ _05702_ _05266_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__mux2_1
XANTENNA__11702__A2 reg_next_pc\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10003_ cpuregs.regs\[16\]\[17\] cpuregs.regs\[17\]\[17\] cpuregs.regs\[18\]\[17\]
+ cpuregs.regs\[19\]\[17\] _04057_ _04060_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__mux4_1
XANTENNA__10910__A0 _04708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15860_ _02613_ _02612_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__or2b_1
XANTENNA__14101__B1 _07834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14811_ _01761_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__clkbuf_1
X_15791_ is_beq_bne_blt_bge_bltu_bgeu instr_jalr _02574_ cpu_state\[3\] VGND VGND
+ VPWR VPWR _02579_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_4_13_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11383__A _03781_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10269__A2 _04979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17530_ clknet_leaf_106_clk _00699_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_14742_ _01713_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__clkbuf_1
X_11954_ _06428_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09754__S1 _04087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10905_ _03618_ _05440_ _05456_ _05478_ _05593_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__o221a_1
X_17461_ clknet_leaf_98_clk _00630_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14673_ _07968_ _08301_ _07969_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__a21oi_1
X_11885_ _06391_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16385__S _02918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output108_A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13624_ net76 decoded_imm\[18\] VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16412_ _02936_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__clkbuf_1
X_10836_ _05377_ _05528_ _05287_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__mux2_1
XANTENNA__09788__A _04283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08692__A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17392_ clknet_leaf_130_clk _00561_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13555_ _07398_ _07401_ VGND VGND VPWR VPWR _07409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16343_ _06949_ cpuregs.regs\[16\]\[3\] _02896_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__mux2_1
X_10767_ _05298_ _05459_ _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__a21o_1
XANTENNA__09292__C1 _03303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12418__S _06689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10727__A _05254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12506_ _06266_ cpuregs.regs\[28\]\[21\] _06737_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16274_ _06949_ cpuregs.regs\[15\]\[3\] _02859_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13486_ _07344_ _07328_ _07325_ VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__a21oi_2
X_10698_ _05397_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__clkbuf_4
X_18013_ clknet_leaf_76_clk _01150_ VGND VGND VPWR VPWR irq_mask\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15225_ _02073_ _02076_ _03687_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12437_ cpuregs.regs\[27\]\[21\] _06578_ _06700_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__mux2_1
XANTENNA__12942__A _06247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13391__A1 _07232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15156_ net126 _01906_ _02008_ _02010_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__o22a_1
X_12368_ cpuregs.regs\[26\]\[21\] _06578_ _06663_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14107_ count_instr\[37\] _07836_ count_instr\[38\] VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__a21o_1
X_11319_ _05934_ _05937_ _05938_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15087_ cpuregs.regs\[28\]\[1\] cpuregs.regs\[29\]\[1\] cpuregs.regs\[30\]\[1\] cpuregs.regs\[31\]\[1\]
+ _01936_ _03647_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_35_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12153__S _06534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12299_ cpuregs.regs\[25\]\[21\] _06578_ _06626_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__mux2_1
X_14038_ _07792_ _07793_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_52_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09028__A _03206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14340__B1 _07997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11154__A0 _05292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10052__S1 _04473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08867__A _03199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13492__B decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15989_ decoded_rd\[0\] _05973_ _06016_ _02704_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__a22o_1
XANTENNA__14643__A1 _08012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08530_ _03237_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17728_ clknet_leaf_74_clk _00897_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09745__S1 _04470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08461_ _03241_ _03244_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17659_ clknet_leaf_72_clk _00828_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_159_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16295__S _02870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_183_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_183_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_147_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16148__A1 net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12328__S _06641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14159__B1 _07877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09013_ _03774_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09637__S _04321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10196__B2 instr_timer VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09681__S0 _04056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13159__S _07093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12063__S _06482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10372__A reg_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09915_ _04632_ _04633_ _04636_ _04149_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__o211a_1
XANTENNA__12998__S _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11145__B1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09846_ irq_pending\[12\] _04007_ _04565_ _04569_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__o22a_1
XANTENNA__10043__S1 _04060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ reg_pc\[11\] decoded_imm\[11\] VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08728_ net103 net71 VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_87_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _03416_ _03423_ _03425_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_1_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_174_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_174_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_139_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11670_ reg_pc\[17\] _06218_ _06093_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10621_ _05230_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09401__A _00071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18136__D alu_out\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10959__A0 _04810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13340_ _04215_ _07202_ _07206_ VGND VGND VPWR VPWR _07207_ sky130_fd_sc_hd__a21oi_1
X_10552_ instr_sra instr_srl instr_srai instr_srli VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15549__S _03272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13271_ _07162_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10483_ cpuregs.regs\[28\]\[31\] cpuregs.regs\[29\]\[31\] cpuregs.regs\[30\]\[31\]
+ cpuregs.regs\[31\]\[31\] _04274_ _04317_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_118_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15010_ _04659_ _01885_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__nor2_1
X_12222_ _06581_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12153_ cpuregs.regs\[24\]\[0\] _06531_ _06534_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__mux2_1
XANTENNA__10282__S1 _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11104_ _03444_ _05398_ _05646_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__o21ai_1
X_16961_ clknet_leaf_183_clk _00135_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12084_ _06497_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15792__B _06863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14689__A _03240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11035_ _05713_ _05667_ _05246_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__mux2_1
X_15912_ _02633_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__buf_4
XANTENNA__12701__S _06836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09975__S1 _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16892_ clknet_leaf_31_clk _00037_ VGND VGND VPWR VPWR mem_rdata_q\[11\] sky130_fd_sc_hd__dfxtp_1
X_18631_ clknet_leaf_160_clk _01691_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_15843_ _03799_ _03885_ _02603_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__and3_1
XANTENNA__15822__B1 decoded_imm_j\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12636__A0 _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18562_ clknet_leaf_138_clk _01627_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10221__S _04430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15774_ timer\[31\] _02567_ _02564_ timer\[30\] _02476_ VGND VGND VPWR VPWR _02568_
+ sky130_fd_sc_hd__a221o_1
X_12986_ cpuregs.regs\[3\]\[1\] _06536_ _07010_ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17513_ clknet_leaf_186_clk _00682_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_14725_ count_cycle\[10\] count_cycle\[11\] count_cycle\[12\] _08353_ VGND VGND VPWR
+ VPWR _08359_ sky130_fd_sc_hd__and4_2
X_18493_ clknet_leaf_184_clk _01558_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11937_ _06418_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_165_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_165_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17444_ clknet_leaf_12_clk _00613_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11868_ _06380_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__clkbuf_1
X_14656_ _03294_ _07968_ _07997_ _08304_ VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13607_ _04708_ _07457_ _07374_ VGND VGND VPWR VPWR _07458_ sky130_fd_sc_hd__mux2_1
X_10819_ _05345_ _05512_ _05287_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17375_ clknet_leaf_21_clk _00544_ VGND VGND VPWR VPWR cpuregs.waddr\[1\] sky130_fd_sc_hd__dfxtp_4
X_11799_ _06116_ reg_next_pc\[31\] _06339_ _06341_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_31_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14587_ _07954_ _07956_ _08221_ VGND VGND VPWR VPWR _08242_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16326_ _07001_ cpuregs.regs\[15\]\[28\] _02881_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__mux2_1
X_13538_ _07364_ _07378_ VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13469_ _07325_ _07326_ _07328_ VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__or3b_1
X_16257_ mem_rdata_q\[5\] _03895_ _03914_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__mux2_1
XANTENNA__15353__A2 _02009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15208_ _02060_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14561__B1 _07997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput204 net204 VGND VGND VPWR VPWR mem_la_addr[20] sky130_fd_sc_hd__buf_1
XANTENNA__13487__B decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput215 net215 VGND VGND VPWR VPWR mem_la_addr[30] sky130_fd_sc_hd__clkbuf_1
X_16188_ net257 net258 _01822_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__a21bo_1
Xoutput226 net226 VGND VGND VPWR VPWR mem_la_wdata[10] sky130_fd_sc_hd__clkbuf_1
XANTENNA__10717__A3 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput237 net237 VGND VGND VPWR VPWR mem_la_wdata[20] sky130_fd_sc_hd__buf_1
XANTENNA__11288__A _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput248 net248 VGND VGND VPWR VPWR mem_la_wdata[30] sky130_fd_sc_hd__buf_1
XANTENNA__15105__A2 _01906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15139_ _01989_ _01993_ _03692_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__o21a_1
Xoutput259 net259 VGND VGND VPWR VPWR mem_la_wstrb[1] sky130_fd_sc_hd__buf_1
X_09700_ _04391_ _04394_ _04395_ _04427_ VGND VGND VPWR VPWR _08399_ sky130_fd_sc_hd__a31o_1
XANTENNA__09966__S1 _04470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12611__S _06788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09631_ _03518_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15408__A3 _02249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11735__B _06118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09562_ cpuregs.regs\[4\]\[5\] cpuregs.regs\[5\]\[5\] cpuregs.regs\[6\]\[5\] cpuregs.regs\[7\]\[5\]
+ _04291_ _04292_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__mux4_1
XFILLER_0_172_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08513_ mem_wordsize\[0\] _03290_ _03295_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__a21o_1
X_09493_ _04081_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_156_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_156_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_65_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15223__A _01937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08444_ _03206_ _03212_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__nand2_2
XFILLER_0_172_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13052__A0 _06941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10367__A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16753__S _03116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08482__D instr_slli VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15369__S _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09875__B decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10814__B _05220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10708__A3 _05394_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15647__A3 _03630_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11118__B1 _05356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12252__A_N cpuregs.waddr\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09829_ cpuregs.regs\[24\]\[12\] cpuregs.regs\[25\]\[12\] cpuregs.regs\[26\]\[12\]
+ cpuregs.regs\[27\]\[12\] _04329_ _04218_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__mux4_1
XANTENNA__14607__A1 _03195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15804__B1 _03895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12840_ _06919_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09709__S1 _04317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12771_ _06882_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_147_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_147_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_68_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15133__A _01984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11722_ _06273_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__buf_2
X_14510_ reg_next_pc\[16\] _07948_ _08171_ _07960_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__a22o_1
XANTENNA__10644__A2 _04566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15490_ cpuregs.regs\[8\]\[23\] cpuregs.regs\[9\]\[23\] cpuregs.regs\[10\]\[23\]
+ cpuregs.regs\[11\]\[23\] _03640_ _03642_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__mux4_1
XFILLER_0_167_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15032__A1 _03303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11653_ _06210_ _06118_ _06211_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__and3b_1
XFILLER_0_83_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14441_ _08087_ _08094_ _08107_ VGND VGND VPWR VPWR _08108_ sky130_fd_sc_hd__o21a_1
XANTENNA__16663__S _03062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14972__A _01863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10604_ _04880_ net81 _05263_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__mux2_1
XANTENNA__11054__C1 _05251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_985 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17160_ clknet_leaf_133_clk _00334_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_14372_ _07917_ _07994_ _08044_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11584_ _06150_ cpuregs.regs\[10\]\[7\] _06086_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09893__S0 _04290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13323_ _07189_ VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__buf_2
X_16111_ _02770_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__buf_4
XFILLER_0_91_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10535_ _05231_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__buf_4
XFILLER_0_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17091_ clknet_leaf_143_clk _00265_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13346__A1 _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13254_ _06422_ _06904_ VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__nand2_4
X_16042_ _02715_ decoded_imm_j\[10\] _02726_ mem_rdata_q\[30\] _02634_ VGND VGND VPWR
+ VPWR _02733_ sky130_fd_sc_hd__a221o_1
X_10466_ _04271_ _05170_ _05171_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_133_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09645__S0 _04325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output175_A net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12205_ cpuregs.regs\[24\]\[17\] _06569_ _06555_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13185_ _07116_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10255__S1 _04276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10397_ _04214_ _05100_ _05104_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15099__A1 _05286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12136_ _06524_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__clkbuf_1
X_17993_ clknet_leaf_103_clk _01130_ VGND VGND VPWR VPWR irq_mask\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13649__A2 _05261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10007__S1 _04074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16944_ clknet_leaf_163_clk _00125_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_12067_ _06297_ cpuregs.regs\[22\]\[25\] _06482_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_8_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11018_ _05219_ _05698_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__nor2_1
XANTENNA__09306__A _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15027__B _01885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12745__A_N cpuregs.waddr\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16875_ _06590_ cpuregs.regs\[14\]\[27\] _03174_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__mux2_1
X_18614_ clknet_leaf_167_clk _01679_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12609__A0 _06132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15826_ decoded_imm_j\[13\] _05983_ _03747_ _02587_ _02596_ VGND VGND VPWR VPWR _01243_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13770__B decoded_imm\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18545_ clknet_leaf_113_clk _01610_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_15757_ timer\[26\] _02552_ _02479_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_138_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_138_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08828__A2 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _07000_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13262__S _07154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15043__A _05200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14708_ _08346_ _08347_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18476_ clknet_leaf_109_clk _01541_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_15688_ timer\[8\] _02503_ _02476_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17427_ clknet_leaf_178_clk _00596_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14639_ _08287_ _08289_ VGND VGND VPWR VPWR _08290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_173_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17358_ clknet_leaf_132_clk _00527_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08880__A _03640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13498__A _03275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16309_ _02858_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16523__A1 _06584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10915__A _05292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17289_ clknet_leaf_135_clk _00463_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09636__S0 _04274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09410__C1 _04027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_1_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15629__A3 _02457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08993_ net39 mem_rdata_q\[15\] _03729_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__mux2_1
XANTENNA__10571__A1 _05205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15218__A _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09216__A _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09614_ _04036_ mem_wordsize\[1\] _04343_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__and3_1
XANTENNA__09650__S _04222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13680__B decoded_imm\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09545_ _04058_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_129_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_129_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13172__S _07104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09476_ _04074_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_80_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10182__S0 _04281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08427_ _03212_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_163_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15888__A _02634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15565__A2 _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16483__S _02968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12516__S _06737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10320_ cpuregs.regs\[12\]\[26\] cpuregs.regs\[13\]\[26\] cpuregs.regs\[14\]\[26\]
+ cpuregs.regs\[15\]\[26\] _04123_ _04124_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10251_ cpuregs.regs\[12\]\[24\] cpuregs.regs\[13\]\[24\] cpuregs.regs\[14\]\[24\]
+ cpuregs.regs\[15\]\[24\] _04217_ _04219_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__mux4_1
XFILLER_0_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10182_ cpuregs.regs\[24\]\[22\] cpuregs.regs\[25\]\[22\] cpuregs.regs\[26\]\[22\]
+ cpuregs.regs\[27\]\[22\] _04281_ _04470_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__mux4_1
XANTENNA__12839__A0 _06184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14990_ _04382_ _01869_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__nor2_1
XANTENNA__11375__B _03878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13941_ _07714_ _07725_ VGND VGND VPWR VPWR _07726_ sky130_fd_sc_hd__and2_1
XANTENNA__15562__S _01907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09180__A1 _03895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13871__A _06053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16660_ _03067_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10865__A2 _05440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15789__C1 _06026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13872_ _06072_ _03298_ VGND VGND VPWR VPWR _07676_ sky130_fd_sc_hd__nand2_1
XANTENNA__15253__A1 _01982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15611_ decoded_imm\[30\] _01933_ _01959_ _02440_ _01934_ VGND VGND VPWR VPWR _02441_
+ sky130_fd_sc_hd__a221o_4
X_12823_ _06910_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__clkbuf_1
X_16591_ _06993_ cpuregs.regs\[18\]\[24\] _03026_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08684__B net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13803__A2 _05170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11391__A _03977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18330_ clknet_leaf_38_clk _01398_ VGND VGND VPWR VPWR mem_16bit_buffer\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15542_ _02374_ _02375_ _03709_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__mux2_1
X_12754_ _06873_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11705_ _06257_ cpuregs.regs\[10\]\[20\] _06258_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__mux2_1
X_18261_ clknet_leaf_29_clk _01332_ VGND VGND VPWR VPWR decoded_imm\[19\] sky130_fd_sc_hd__dfxtp_4
X_12685_ _06834_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__clkbuf_1
X_15473_ _02309_ _02310_ _03687_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__mux2_1
XANTENNA__16393__S _02918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ clknet_leaf_12_clk _00386_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11636_ _06195_ _06196_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__nor2_1
X_14424_ _07925_ _07928_ _08076_ VGND VGND VPWR VPWR _08092_ sky130_fd_sc_hd__and3_1
XFILLER_0_170_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18192_ clknet_leaf_29_clk _01263_ VGND VGND VPWR VPWR instr_lw sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17143_ clknet_leaf_156_clk _00317_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11567_ _06072_ _03321_ _06098_ _06134_ _06118_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__a221o_1
XANTENNA__12426__S _06689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14355_ _07915_ _08016_ VGND VGND VPWR VPWR _08029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11510__B_N _06081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10518_ _05212_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__clkbuf_4
X_13306_ _06993_ cpuregs.regs\[5\]\[24\] _07176_ VGND VGND VPWR VPWR _07181_ sky130_fd_sc_hd__mux2_1
X_14286_ _05941_ _06317_ _07944_ _05942_ VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__o211a_2
XANTENNA__15713__C1 _07775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17074_ clknet_leaf_110_clk _00248_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_11498_ irq_state\[1\] VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08787__A_N net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13237_ _07144_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__clkbuf_1
X_16025_ decoded_imm\[3\] _02720_ _02721_ _02722_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__o22a_1
X_10449_ _05153_ _05154_ _04065_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_161_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13168_ _06991_ cpuregs.regs\[4\]\[23\] _07104_ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__mux2_1
XANTENNA__15167__S1 _01992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12119_ _06515_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__clkbuf_1
X_17976_ clknet_leaf_44_clk _01113_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dfxtp_2
X_13099_ _07071_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15492__A1 _03675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16927_ clknet_leaf_138_clk _00108_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11502__B1 reg_next_pc\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16568__S _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_176_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16858_ _06573_ cpuregs.regs\[14\]\[19\] _03163_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__mux2_1
XANTENNA__08875__A _00064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14596__B _07958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15809_ _05960_ _03634_ _03864_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__and3_1
XANTENNA__15795__A2 _03226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16789_ _03136_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09330_ _04064_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__buf_8
X_18528_ clknet_leaf_160_clk _01593_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09261_ _03840_ _03995_ _03999_ _03888_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_173_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18459_ clknet_leaf_181_clk _01524_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09192_ mem_rdata_q\[14\] VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_99_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09857__S0 _04579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12230__A1 _06586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12336__S _06641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15932__B_N mem_rdata_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10219__S1 _04470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_129_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08769__B net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12071__S _06482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08976_ _03229_ _03237_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_90_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15890__B _02611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12297__A1 _06575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15382__S _02110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09528_ reg_pc\[5\] decoded_imm\[5\] VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_27_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09459_ reg_pc\[3\] decoded_imm\[3\] VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_899 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12470_ _06125_ cpuregs.regs\[28\]\[4\] _06715_ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11421_ _03305_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12221__A1 _06580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10458__S1 _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11150__S _04745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14140_ count_instr\[48\] count_instr\[47\] count_instr\[46\] _07859_ VGND VGND VPWR
+ VPWR _07864_ sky130_fd_sc_hd__and4_1
XFILLER_0_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11352_ _05962_ _05966_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10274__B decoded_imm\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10783__A1 _03518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15397__S1 _02047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10303_ net50 _04811_ _04667_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__a21o_2
XFILLER_0_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14071_ count_instr\[26\] _07811_ count_instr\[27\] VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11283_ _05857_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__buf_2
X_13022_ _07030_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13721__A1 _07232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10234_ _03637_ _04945_ _04673_ _04946_ _04266_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_167_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13077__S _07057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17830_ clknet_leaf_57_clk _00999_ VGND VGND VPWR VPWR reg_next_pc\[7\] sky130_fd_sc_hd__dfxtp_1
X_10165_ net80 VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__buf_4
XFILLER_0_100_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15474__B2 _02004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17761_ clknet_leaf_90_clk _00930_ VGND VGND VPWR VPWR count_instr\[32\] sky130_fd_sc_hd__dfxtp_1
X_10096_ _04046_ _04810_ _04752_ _04812_ _04202_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__a221o_1
X_14973_ _01862_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13805__S _07224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16712_ _06978_ cpuregs.regs\[19\]\[17\] _03087_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__mux2_1
X_13924_ _06053_ VGND VGND VPWR VPWR _07714_ sky130_fd_sc_hd__clkbuf_2
X_17692_ clknet_leaf_119_clk _00861_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08695__A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15226__B2 _02037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10394__S0 _04123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11401__C_N _03867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16643_ _03058_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__clkbuf_1
X_13855_ cpuregs.regs\[0\]\[24\] VGND VGND VPWR VPWR _07667_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12806_ _06900_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__clkbuf_1
X_16574_ _06976_ cpuregs.regs\[18\]\[16\] _03015_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__mux2_1
X_10998_ _03472_ _05678_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__or2_1
X_13786_ _05086_ decoded_imm\[28\] VGND VGND VPWR VPWR _07624_ sky130_fd_sc_hd__nand2_1
XANTENNA__09456__A2 _04021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18313_ clknet_leaf_35_clk _01381_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dfxtp_1
X_15525_ cpuregs.regs\[28\]\[25\] cpuregs.regs\[29\]\[25\] cpuregs.regs\[30\]\[25\]
+ cpuregs.regs\[31\]\[25\] _01999_ _02000_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12737_ _03364_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12945__A _06256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14737__B1 _07826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18244_ clknet_leaf_25_clk _01315_ VGND VGND VPWR VPWR decoded_imm\[2\] sky130_fd_sc_hd__dfxtp_2
X_15456_ cpuregs.regs\[24\]\[21\] cpuregs.regs\[25\]\[21\] cpuregs.regs\[26\]\[21\]
+ cpuregs.regs\[27\]\[21\] _02074_ _02075_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12668_ _06078_ cpuregs.regs\[12\]\[0\] _06825_ VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14407_ _08035_ _08076_ _07995_ _07924_ VGND VGND VPWR VPWR _08077_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08416__A0 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11619_ _06071_ reg_next_pc\[11\] _06181_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12156__S _06534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18175_ clknet_leaf_24_clk _01246_ VGND VGND VPWR VPWR decoded_imm_j\[16\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15387_ cpuregs.regs\[24\]\[17\] cpuregs.regs\[25\]\[17\] cpuregs.regs\[26\]\[17\]
+ cpuregs.regs\[27\]\[17\] _02221_ _02222_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12599_ _06078_ cpuregs.regs\[30\]\[0\] _06788_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17126_ clknet_leaf_137_clk _00300_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14338_ _08002_ _08006_ _08013_ _07905_ reg_next_pc\[2\] VGND VGND VPWR VPWR _00994_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11995__S _06446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17057_ clknet_leaf_183_clk _00231_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_14269_ reg_next_pc\[22\] _05898_ _07942_ _07955_ VGND VGND VPWR VPWR _07956_ sky130_fd_sc_hd__o211a_2
XANTENNA__09916__B1 _04613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16008_ cpuregs.raddr2\[3\] _05983_ _05984_ _05985_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_55_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ net123 net91 VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__and2b_1
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08761_ net125 net93 VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__nor2_1
X_17959_ clknet_leaf_191_clk _01096_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dfxtp_1
XANTENNA__15560__S1 _02000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10829__A2 _05220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08692_ net115 net83 VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14400__A _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15768__A2 _02486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13779__A1 _03275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09213__B _03880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09313_ _04048_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_145_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09244_ _03748_ _03790_ _03984_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__and3_1
XANTENNA__14728__B1 _07826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09175_ _03762_ _03892_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10375__A reg_pc\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16761__S _03116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13400__B1 _07210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15940__A2 _02650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13951__A1 _03320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15885__B _02620_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15377__S _01907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13703__A1 _03631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09375__S _04040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09907__B1 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11714__A0 _06266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11190__A1 _04198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08959_ cpuregs.regs\[16\]\[4\] cpuregs.regs\[17\]\[4\] cpuregs.regs\[18\]\[4\] cpuregs.regs\[19\]\[4\]
+ _03661_ _03662_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__mux4_1
XANTENNA__15551__S1 _01980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_162_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _06184_ cpuregs.regs\[21\]\[11\] _06435_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__mux2_1
XANTENNA__14310__A _03364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16405__A0 _06941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13219__A0 _06974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10921_ _03564_ _05608_ _05390_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__mux2_1
XANTENNA__11653__B _06118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18139__D alu_out\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15303__S1 _01971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13640_ net77 decoded_imm\[19\] VGND VGND VPWR VPWR _07488_ sky130_fd_sc_hd__nand2_1
X_10852_ _05543_ _05510_ _05479_ _05441_ _05266_ _05243_ VGND VGND VPWR VPWR _05544_
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_123_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15978__B_N mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _04602_ _07315_ _07382_ _07254_ VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__o211a_1
X_10783_ _03510_ _03518_ _05229_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_51_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_137_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15310_ _02037_ _02156_ _02006_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__a21o_1
XANTENNA__15141__A _01995_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14719__B1 _07826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12522_ _06328_ cpuregs.regs\[28\]\[29\] _06737_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__mux2_1
X_16290_ _02871_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15241_ cpuregs.regs\[24\]\[9\] cpuregs.regs\[25\]\[9\] cpuregs.regs\[26\]\[9\] cpuregs.regs\[27\]\[9\]
+ _02069_ _02070_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__mux4_1
XANTENNA__16671__S _03039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12453_ cpuregs.regs\[27\]\[29\] _06594_ _06700_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15931__A2 _02650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11404_ _05976_ _06007_ _06008_ _06012_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__or4b_1
XFILLER_0_151_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15172_ _02020_ _02025_ _02006_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_10_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12384_ cpuregs.regs\[26\]\[29\] _06594_ _06663_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09610__A2 _04165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11953__A0 _06114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11335_ reg_out\[30\] _05941_ _05951_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__o21a_1
X_14123_ count_instr\[43\] _07843_ _07848_ VGND VGND VPWR VPWR _07852_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15695__A1 _04447_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14054_ _07803_ _07804_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__nor2_1
X_11266_ _05891_ _05894_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__and2_2
XANTENNA__11705__A0 _06257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output255_A net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13005_ cpuregs.regs\[3\]\[10\] _06554_ _07021_ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__mux2_1
X_10217_ _04928_ _04929_ _04065_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10224__S _04064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11197_ _05829_ _05836_ _05837_ _05839_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__a31o_4
XFILLER_0_20_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17813_ clknet_leaf_63_clk _00982_ VGND VGND VPWR VPWR reg_pc\[21\] sky130_fd_sc_hd__dfxtp_1
X_10148_ cpuregs.regs\[28\]\[21\] cpuregs.regs\[29\]\[21\] cpuregs.regs\[30\]\[21\]
+ cpuregs.regs\[31\]\[21\] _04758_ _04759_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17744_ clknet_leaf_87_clk _00913_ VGND VGND VPWR VPWR count_instr\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_max_cap301_A _04099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14956_ _01853_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__clkbuf_1
X_10079_ _04054_ _04795_ _04225_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_50_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13907_ _03323_ _07678_ _07682_ net162 VGND VGND VPWR VPWR _07702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15035__B _01885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18049__D _01154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17675_ clknet_leaf_160_clk _00844_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_14887_ _03400_ _01811_ _07224_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__o21a_1
XANTENNA__16846__S _03163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16626_ _03049_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13838_ _07658_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09429__A2 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10119__S0 _04275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10894__S _05390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16557_ _06959_ cpuregs.regs\[18\]\[8\] _03004_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__mux2_1
X_13769_ _07558_ _07569_ _07603_ _07605_ _07607_ VGND VGND VPWR VPWR _07608_ sky130_fd_sc_hd__o311a_1
Xclkbuf_leaf_42_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__13270__S _07154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15508_ _01989_ _02343_ _02017_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16488_ _02976_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18227_ clknet_leaf_32_clk _01298_ VGND VGND VPWR VPWR decoded_rd\[0\] sky130_fd_sc_hd__dfxtp_1
X_15439_ _02111_ _02278_ _01968_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__o21a_1
XANTENNA__10195__A _04908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15922__A2 _02617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12736__A2 _03384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09062__A0 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18158_ clknet_leaf_40_clk clear_prefetched_high_word VGND VGND VPWR VPWR clear_prefetched_high_word_q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17109_ clknet_leaf_116_clk _00283_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18089_ clknet_leaf_101_clk _01193_ VGND VGND VPWR VPWR timer\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16883__A0 _06598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15686__A1 _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09931_ cpuregs.regs\[0\]\[15\] cpuregs.regs\[1\]\[15\] cpuregs.regs\[2\]\[15\] cpuregs.regs\[3\]\[15\]
+ _04232_ _04233_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09862_ cpuregs.regs\[4\]\[13\] cpuregs.regs\[5\]\[13\] cpuregs.regs\[6\]\[13\] cpuregs.regs\[7\]\[13\]
+ _04273_ _04283_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_70_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11172__A1 _04038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11172__B2 _03297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08813_ _03472_ _03577_ _03578_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__a21oi_1
X_09793_ cpuregs.regs\[28\]\[11\] cpuregs.regs\[29\]\[11\] cpuregs.regs\[30\]\[11\]
+ cpuregs.regs\[31\]\[11\] _04282_ _04285_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__mux4_1
X_08744_ net97 VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_169_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09668__A2 _04104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11473__B _03428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08675_ net119 net87 VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__nand2_1
XANTENNA__15297__S0 _02074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14949__A0 net209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14784__B _08350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12424__A1 _06565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13180__S _07104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_146_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10530__S0 _05230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15374__B1 _02215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15896__A _02612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09227_ _03895_ _03958_ _03967_ _03927_ _03968_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16491__S _02968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15913__A2 _02625_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09158_ _03911_ _03878_ _03908_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10738__A1 _05277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09089_ _03753_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11120_ _05601_ _05684_ _05791_ _05281_ _05793_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__a221o_1
XANTENNA__15221__S0 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11051_ _05044_ _05013_ _05230_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_164_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10002_ cpuregs.regs\[20\]\[17\] cpuregs.regs\[21\]\[17\] cpuregs.regs\[22\]\[17\]
+ cpuregs.regs\[23\]\[17\] _04472_ _04473_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__mux4_1
XANTENNA__10910__A1 _04642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _01759_ _01753_ _01760_ VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__and3b_1
XANTENNA__15136__A _03642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _04156_ _03292_ _03271_ _07680_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__a31oi_1
XANTENNA__10349__S0 _04207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09134__A _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14741_ _08368_ _08350_ _01712_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__and3b_1
XFILLER_0_87_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11953_ _06114_ cpuregs.regs\[21\]\[3\] _06424_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__mux2_1
XANTENNA__15288__S0 _01973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10904_ _03617_ _05301_ _05356_ _03619_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__o2bb2a_1
X_17460_ clknet_leaf_151_clk _00629_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_805 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14672_ _08309_ _08315_ _08318_ _08055_ VGND VGND VPWR VPWR _08320_ sky130_fd_sc_hd__a31o_1
X_11884_ _06114_ cpuregs.regs\[20\]\[3\] _06387_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16411_ _06949_ cpuregs.regs\[29\]\[3\] _02932_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13623_ net76 decoded_imm\[18\] VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10835_ _05527_ _05460_ _05246_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__mux2_1
X_17391_ clknet_leaf_146_clk _00560_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13612__B1 _03311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08692__B net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16342_ _02899_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__clkbuf_1
X_13554_ _07406_ _07407_ VGND VGND VPWR VPWR _07408_ sky130_fd_sc_hd__nand2_1
X_10766_ _03614_ _05222_ _05251_ _05461_ _05462_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10977__A1 _05544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10727__B _05261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12505_ _06738_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16273_ _02862_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__clkbuf_1
X_13485_ net96 decoded_imm\[7\] VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__or2_1
X_10697_ instr_and instr_andi VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__nor2_2
XANTENNA__15904__A2 _02617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18012_ clknet_leaf_76_clk _01149_ VGND VGND VPWR VPWR irq_mask\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13915__A1 _03335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15224_ cpuregs.regs\[28\]\[8\] cpuregs.regs\[29\]\[8\] cpuregs.regs\[30\]\[8\] cpuregs.regs\[31\]\[8\]
+ _02074_ _02075_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__mux4_1
X_12436_ _06701_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10729__A1 _05361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15155_ decoded_imm\[5\] _02009_ _01963_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__a21o_1
X_12367_ _06664_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15212__S0 _01979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16865__A0 _06580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15668__A1 _07250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output82_A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14106_ count_instr\[35\] _07831_ _07839_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__and3_1
X_11318_ _05925_ _05929_ _05932_ _05937_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__and4_1
XANTENNA__09309__A reg_next_pc\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15086_ _03656_ _01944_ _00068_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__a21o_1
X_12298_ _06627_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14340__A1 _03294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14037_ count_instr\[16\] _07789_ _07790_ VGND VGND VPWR VPWR _07793_ sky130_fd_sc_hd__o21ai_1
X_11249_ _05878_ _05881_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_52_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11154__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10889__S _05413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10362__C1 _04188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16093__A1 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15046__A _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15988_ _03816_ _03737_ _02628_ _02699_ _02703_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__a41o_1
XFILLER_0_89_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17727_ clknet_leaf_74_clk _00896_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dfxtp_1
X_14939_ _01844_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16576__S _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08460_ net67 mem_wordsize\[2\] _03243_ mem_wordsize\[0\] VGND VGND VPWR VPWR _03244_
+ sky130_fd_sc_hd__a22o_1
X_17658_ clknet_leaf_71_clk _00827_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dfxtp_2
XANTENNA__15053__C1 _03654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16609_ cpuregs.regs\[1\]\[0\] _06077_ _03040_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12609__S _06788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17589_ clknet_leaf_98_clk _00758_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11513__S _06086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11090__B1 _05367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09012_ mem_16bit_buffer\[10\] _03773_ _03727_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15451__S0 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10653__A net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10196__A2 _04308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16856__A0 _06571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09681__S1 _04091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10372__B decoded_imm\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09914_ count_cycle\[14\] _04165_ _04635_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__a21o_1
XANTENNA__11145__A1 _03407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11145__B2 _04422_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09845_ _03637_ _04566_ _04568_ _03225_ _04266_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08777__B net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16084__A1 _03767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16084__B2 _03215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ reg_pc\[11\] decoded_imm\[11\] VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__nor2_1
XANTENNA__15831__A1 decoded_imm_j\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _03491_ _03492_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__or2b_2
XTAP_TAPCELL_ROW_87_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09889__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08944__S0 _03649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09510__B2 _04187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08658_ timer\[31\] _03424_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14398__B2 _08033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08589_ _03366_ _03367_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__nor2_4
XFILLER_0_77_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10620_ _05322_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10959__A1 _04754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ _05254_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13270_ _06957_ cpuregs.regs\[5\]\[7\] _07154_ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__mux2_1
X_10482_ _04289_ _05186_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13373__A2 _04262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12221_ cpuregs.regs\[24\]\[22\] _06580_ _06576_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__mux2_1
XANTENNA__18730__A net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12152_ _06533_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__clkbuf_8
X_11103_ _03444_ _05215_ _05213_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__a21o_1
XANTENNA__13874__A _07677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16960_ clknet_leaf_172_clk _00134_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12083_ _06078_ cpuregs.regs\[23\]\[0\] _06496_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__mux2_1
XANTENNA__15792__C _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11136__B2 _04422_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11034_ _05013_ _04959_ _04945_ net81 _05264_ _05232_ VGND VGND VPWR VPWR _05713_
+ sky130_fd_sc_hd__mux4_1
X_15911_ _02611_ _02647_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__and2_1
X_16891_ clknet_leaf_31_clk _00036_ VGND VGND VPWR VPWR mem_rdata_q\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13085__S _07057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16075__A1 decoded_imm\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18630_ clknet_leaf_129_clk _01690_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11394__A _03781_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16075__B2 mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15842_ instr_lui _05987_ _06016_ _02601_ _02604_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__a221o_1
XANTENNA__15283__C1 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18561_ clknet_leaf_156_clk _01626_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15822__B2 _03636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output120_A net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15773_ _03424_ _02560_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__nor2_1
X_12985_ _07011_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output218_A net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17512_ clknet_leaf_173_clk _00681_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14724_ _08358_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08935__S0 _03658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18492_ clknet_leaf_186_clk _01557_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11936_ _06320_ cpuregs.regs\[20\]\[28\] _06409_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17443_ clknet_leaf_14_clk _00612_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14655_ _07998_ _08301_ VGND VGND VPWR VPWR _08304_ sky130_fd_sc_hd__or2_1
X_11867_ _06328_ cpuregs.regs\[11\]\[29\] _06370_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13606_ _03276_ _07449_ _07450_ _07456_ VGND VGND VPWR VPWR _07457_ sky130_fd_sc_hd__a31o_1
XFILLER_0_157_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10818_ _05511_ _05442_ _05295_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__mux2_1
X_17374_ clknet_leaf_20_clk _00543_ VGND VGND VPWR VPWR cpuregs.waddr\[0\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_172_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14586_ _08239_ _08240_ VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__nand2_1
X_11798_ _06072_ _03331_ _06098_ _06340_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11072__B1 _05221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16325_ _02889_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13537_ _07209_ _04562_ _07211_ reg_pc\[12\] _07221_ VGND VGND VPWR VPWR _07392_
+ sky130_fd_sc_hd__a221o_1
X_10749_ _05348_ _05329_ _05351_ _05346_ _05277_ _05288_ VGND VGND VPWR VPWR _05447_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__16425__A _02931_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15433__S0 _02085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15889__B2 is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16256_ _02852_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__clkbuf_1
X_13468_ _07297_ _07311_ _07309_ _07327_ VGND VGND VPWR VPWR _07328_ sky130_fd_sc_hd__a31o_1
XFILLER_0_113_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14010__B1 _07759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15207_ net128 _02059_ _01905_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12419_ _06692_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14561__A1 _03294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16187_ net295 _01822_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__or2_1
Xoutput205 net205 VGND VGND VPWR VPWR mem_la_addr[21] sky130_fd_sc_hd__buf_1
X_13399_ _07259_ _07260_ _07261_ VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput216 net216 VGND VGND VPWR VPWR mem_la_addr[31] sky130_fd_sc_hd__buf_1
XFILLER_0_112_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput227 net227 VGND VGND VPWR VPWR mem_la_wdata[11] sky130_fd_sc_hd__buf_1
Xoutput238 net238 VGND VGND VPWR VPWR mem_la_wdata[21] sky130_fd_sc_hd__clkbuf_1
X_15138_ cpuregs.regs\[24\]\[5\] cpuregs.regs\[25\]\[5\] cpuregs.regs\[26\]\[5\] cpuregs.regs\[27\]\[5\]
+ _01990_ _01992_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__mux4_1
Xoutput249 net249 VGND VGND VPWR VPWR mem_la_wdata[31] sky130_fd_sc_hd__buf_1
XFILLER_0_121_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_34_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15069_ _03679_ _01928_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_4_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__08878__A _03642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16066__A1 instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16066__B2 mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10886__B1 _05367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09630_ _04347_ _04351_ _04356_ _04357_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14077__B1 _07775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09561_ _04276_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__buf_4
XANTENNA__13723__S _07224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08512_ instr_lw _03291_ _03287_ instr_sw _03294_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__a221o_1
XANTENNA__08926__S0 _03658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09492_ _04220_ _04221_ _04223_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16471__B_N _06082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08443_ _03208_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09256__A0 mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13959__A _07737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14001__B1 _07759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13355__A2 _07221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10169__A2 _04008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15385__S _02110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08782__A2 _03518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15647__A4 _07905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16057__A1 decoded_imm\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09828_ _04214_ _04551_ _04237_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_6_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15804__B2 _06016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09759_ cpuregs.regs\[0\]\[10\] cpuregs.regs\[1\]\[10\] cpuregs.regs\[2\]\[10\] cpuregs.regs\[3\]\[10\]
+ _04232_ _04233_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_61_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13633__S _07374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_1008 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12770_ cpuregs.regs\[9\]\[11\] _06557_ _06880_ VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11721_ _06226_ reg_next_pc\[22\] _06270_ _06272_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__a211o_2
XFILLER_0_166_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10644__A3 _04602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15032__A2 _04022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14440_ decoded_imm_j\[10\] _07928_ _08096_ VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__a21oi_1
X_11652_ reg_pc\[14\] reg_pc\[13\] _06187_ reg_pc\[15\] VGND VGND VPWR VPWR _06211_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14240__B1 _07934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10603_ _05304_ _05305_ _05232_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__mux2_1
X_14371_ _08035_ _08036_ _08037_ _08043_ VGND VGND VPWR VPWR _08044_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_107_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11583_ _06149_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__buf_2
XFILLER_0_65_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_172_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16110_ _02769_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__buf_2
XFILLER_0_107_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13322_ _03312_ _03274_ VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09893__S1 _04276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10534_ _04036_ _04160_ _04039_ _04198_ _05235_ _05237_ VGND VGND VPWR VPWR _05238_
+ sky130_fd_sc_hd__mux4_1
X_17090_ clknet_leaf_181_clk _00264_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_70_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13346__A2 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16041_ decoded_imm\[9\] _02711_ _02732_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__o21a_1
XANTENNA__11389__A _03756_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10465_ irq_mask\[30\] _04308_ timer\[30\] _04023_ _04026_ VGND VGND VPWR VPWR _05171_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13253_ _07152_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09645__S1 _04317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12204_ _06231_ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__buf_2
X_13184_ _07007_ cpuregs.regs\[4\]\[31\] _07081_ VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__mux2_1
X_10396_ _04052_ _05103_ _00073_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__a21o_1
XANTENNA__15099__A2 _01906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12135_ _06297_ cpuregs.regs\[23\]\[25\] _06518_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__mux2_1
XANTENNA__12712__S _06847_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17992_ clknet_leaf_104_clk _01129_ VGND VGND VPWR VPWR irq_mask\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08698__A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16943_ clknet_leaf_117_clk _00124_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_12066_ _06487_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16048__B2 _02612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11017_ _03469_ _05697_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__xor2_1
XANTENNA__09722__B2 _04024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09306__B _04038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16874_ _03181_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10332__A2 _04165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18613_ clknet_leaf_163_clk _01678_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_15825_ _05970_ _02594_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__nor2_2
XFILLER_0_59_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15756_ timer\[26\] _02552_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__nor2_1
X_18544_ clknet_leaf_105_clk _01609_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12968_ _06999_ cpuregs.regs\[31\]\[27\] _06985_ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10096__A1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14707_ count_cycle\[6\] _08343_ _07877_ VGND VGND VPWR VPWR _08347_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09322__A _04056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15043__B _01863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10096__B2 _04812_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11919_ _06386_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__buf_6
XFILLER_0_59_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18475_ clknet_leaf_124_clk _01540_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15559__B1 _03692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10468__A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15687_ timer\[0\] _03416_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__or2_1
XANTENNA__16854__S _03163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12159__S _06534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12899_ _06131_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__buf_2
XANTENNA__15023__A2 _01863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17426_ clknet_leaf_140_clk _00595_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13034__A1 _06584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14638_ _08272_ _08280_ _08288_ VGND VGND VPWR VPWR _08289_ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14882__B _01753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17357_ clknet_leaf_127_clk _00526_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14569_ _08219_ _08225_ VGND VGND VPWR VPWR _08226_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11596__A1 _06116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16308_ _02880_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17288_ clknet_leaf_115_clk _00462_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16239_ net53 mem_16bit_buffer\[12\] _02830_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09636__S1 _04317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10020__B2 _04187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12622__S _06799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14403__A decoded_imm_j\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08992_ _03753_ _03203_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_118_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16039__A1 decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09216__B _03892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10142__S _04430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15247__C1 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09613_ net38 net56 _04039_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__mux2_1
XANTENNA__15798__A0 latched_compr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15234__A _01918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09544_ _04274_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10087__A1 _04483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11481__B _03428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09572__S0 _04217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09475_ _04072_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__buf_6
XANTENNA__12069__S _06482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10378__A net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10182__S1 _04470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08426_ mem_16bit_buffer\[1\] _03211_ _03205_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13576__A2 _07211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11587__A1 alu_out_q\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10317__S _04077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11339__A1 _05174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13733__C1 _07283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10250_ count_instr\[24\] _04145_ count_cycle\[24\] _03253_ _04961_ VGND VGND VPWR
+ VPWR _04962_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10181_ cpuregs.regs\[28\]\[22\] cpuregs.regs\[29\]\[22\] cpuregs.regs\[30\]\[22\]
+ cpuregs.regs\[31\]\[22\] _04281_ _04470_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__mux4_1
XANTENNA__14289__B1 _07968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11148__S _04745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13940_ _03358_ _07704_ _07705_ net141 VGND VGND VPWR VPWR _07725_ sky130_fd_sc_hd__a22o_1
X_13871_ _06053_ VGND VGND VPWR VPWR _07675_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15610_ _02430_ _02433_ _02436_ _02439_ _01968_ _03639_ VGND VGND VPWR VPWR _02440_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__15144__A _01995_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12822_ _06114_ cpuregs.regs\[6\]\[3\] _06906_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__mux2_1
X_16590_ _03030_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11275__B1 _05902_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15541_ cpuregs.regs\[28\]\[26\] cpuregs.regs\[29\]\[26\] cpuregs.regs\[30\]\[26\]
+ cpuregs.regs\[31\]\[26\] _03645_ _03647_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__mux4_1
XANTENNA__09563__S0 _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12753_ cpuregs.regs\[9\]\[3\] _06540_ _06869_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__mux2_1
XANTENNA__14983__A _04240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11704_ _06085_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__clkbuf_8
X_18260_ clknet_leaf_31_clk _01331_ VGND VGND VPWR VPWR decoded_imm\[18\] sky130_fd_sc_hd__dfxtp_4
X_15472_ cpuregs.regs\[12\]\[22\] cpuregs.regs\[13\]\[22\] cpuregs.regs\[14\]\[22\]
+ cpuregs.regs\[15\]\[22\] _02074_ _02075_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__mux4_1
XFILLER_0_167_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12684_ _06157_ cpuregs.regs\[12\]\[8\] _06825_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__mux2_1
XANTENNA__14213__B1 _07901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17211_ clknet_leaf_12_clk _00385_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14423_ reg_next_pc\[9\] _07948_ _08081_ _08091_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__a22o_1
X_11635_ reg_pc\[13\] _06187_ _06075_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__o21ai_1
X_18191_ clknet_leaf_29_clk _01262_ VGND VGND VPWR VPWR instr_lh sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12707__S _06836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11578__A1 _06116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17142_ clknet_leaf_126_clk _00316_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_14354_ _08017_ _08023_ _08026_ VGND VGND VPWR VPWR _08028_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11566_ reg_out\[6\] alu_out_q\[6\] latched_stalu VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13305_ _07180_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10250__B2 _03253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10517_ instr_or instr_ori VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__nor2_4
X_17073_ clknet_leaf_162_clk _00247_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_14285_ reg_pc\[27\] _07953_ _07966_ _07960_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11497_ irq_state\[0\] VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16024_ _02715_ decoded_imm_j\[3\] _02716_ mem_rdata_q\[10\] _02633_ VGND VGND VPWR
+ VPWR _02722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13236_ _06991_ cpuregs.regs\[8\]\[23\] _07140_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10448_ cpuregs.regs\[16\]\[30\] cpuregs.regs\[17\]\[30\] cpuregs.regs\[18\]\[30\]
+ cpuregs.regs\[19\]\[30\] _04472_ _04473_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09943__B2 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13167_ _07107_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__clkbuf_1
X_10379_ net53 _04811_ _04667_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12118_ _06232_ cpuregs.regs\[23\]\[17\] _06507_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17975_ clknet_leaf_44_clk _01112_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dfxtp_2
X_13098_ _06989_ cpuregs.regs\[7\]\[22\] _07068_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12049_ _06478_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__clkbuf_1
X_16926_ clknet_leaf_149_clk _00107_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16857_ _03172_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14596__C _07992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15808_ _02586_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__buf_2
X_16788_ _06571_ cpuregs.regs\[13\]\[18\] _03127_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14452__B1 _07947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15739_ _02540_ _02541_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__nand2_1
X_18527_ clknet_leaf_126_clk _01592_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09260_ _03892_ _03894_ _03998_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18458_ clknet_leaf_171_clk _01523_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16744__A2 _07274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08891__A _00067_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17409_ clknet_leaf_15_clk _00578_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_09191_ _03838_ _03934_ _03939_ _03888_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12617__S _06788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18389_ clknet_leaf_14_clk _01454_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09857__S1 _04284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12518__A0 _06312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08975_ _03736_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__16759__S _03116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09698__B1 _04425_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14691__B1 _07675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09793__S0 _04282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08785__B net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11492__A _06065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09527_ reg_pc\[5\] decoded_imm\[5\] VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_27_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16494__S _02979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15618__S0 _02046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09458_ _04010_ _04167_ _04190_ _04150_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08409_ _03194_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15943__B1 _02665_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09389_ _00069_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__buf_6
XFILLER_0_163_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14308__A _03379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11420_ _06006_ _03763_ _05995_ _06023_ _06025_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__a41o_1
XFILLER_0_117_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14027__B _07778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11351_ _03948_ _05964_ _05965_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10302_ net84 VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_130_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14070_ _03304_ VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__clkbuf_4
X_11282_ _05908_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13021_ cpuregs.regs\[3\]\[18\] _06571_ _07021_ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__mux2_1
X_10233_ net48 _04745_ _04666_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15459__C1 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10164_ _04821_ _04824_ _04877_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__nand3_1
XANTENNA__09137__A _03891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16669__S _03062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14978__A _04142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16671__A1 _06335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10095_ net43 _04811_ _04667_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__a21o_1
X_17760_ clknet_leaf_90_clk _00929_ VGND VGND VPWR VPWR count_instr\[31\] sky130_fd_sc_hd__dfxtp_1
X_14972_ _01863_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08976__A _03229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14682__B1 _08050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11496__A0 reg_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13923_ _07713_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__clkbuf_1
X_16711_ _03094_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10299__B2 _04187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09784__S0 _04282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17691_ clknet_leaf_105_clk _00860_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10394__S1 _04124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16642_ cpuregs.regs\[1\]\[16\] _06223_ _03051_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__mux2_1
X_13854_ _07666_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11248__A0 reg_next_pc\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12805_ cpuregs.regs\[9\]\[28\] _06592_ _06891_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__mux2_1
XANTENNA_output200_A net200 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16573_ _03021_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__clkbuf_1
X_13785_ _07611_ _07622_ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__nand2_1
X_10997_ _03472_ _05678_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11799__A1 _06116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15524_ _02012_ _02358_ _02017_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__o21a_1
X_18312_ clknet_leaf_35_clk _01380_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12736_ _03309_ _03384_ _06053_ _06861_ VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_123_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18243_ clknet_leaf_22_clk _01314_ VGND VGND VPWR VPWR decoded_imm\[1\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__10471__B2 _05176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15455_ cpuregs.regs\[28\]\[21\] cpuregs.regs\[29\]\[21\] cpuregs.regs\[30\]\[21\]
+ cpuregs.regs\[31\]\[21\] _01999_ _02000_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12667_ _06824_ VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12437__S _06700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14406_ _07921_ _07924_ _08048_ VGND VGND VPWR VPWR _08076_ sky130_fd_sc_hd__and3_1
X_11618_ irq_state\[1\] _03335_ _06065_ _06180_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__a22o_1
XANTENNA__09613__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18174_ clknet_leaf_31_clk _01245_ VGND VGND VPWR VPWR decoded_imm_j\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_170_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15386_ cpuregs.regs\[28\]\[17\] cpuregs.regs\[29\]\[17\] cpuregs.regs\[30\]\[17\]
+ cpuregs.regs\[31\]\[17\] _01908_ _01909_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__mux4_1
X_12598_ _06787_ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17125_ clknet_leaf_148_clk _00299_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14337_ _08010_ _08011_ _08012_ VGND VGND VPWR VPWR _08013_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_170_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11549_ _06072_ _03327_ _06098_ _06117_ _06118_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12961__A _06296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15698__C1 _06026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17056_ clknet_leaf_186_clk _00230_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_94_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14268_ _05909_ _06271_ VGND VGND VPWR VPWR _07955_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09916__A1 _03638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13268__S _07154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16007_ cpuregs.raddr2\[2\] _05974_ _05980_ _05982_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__a22o_1
X_13219_ _06974_ cpuregs.regs\[8\]\[15\] _07129_ VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__mux2_1
XANTENNA__15049__A _03671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09916__B2 _03226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14199_ _07899_ _07902_ _07906_ reg_pc\[1\] VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__a22o_1
XANTENNA__11296__B _05915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14888__A _05205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08760_ _03523_ _03525_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__and2_1
XANTENNA__12900__S _06943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17958_ clknet_leaf_191_clk _01095_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dfxtp_1
XANTENNA__14673__B1 _07969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16909_ clknet_leaf_6_clk _00054_ VGND VGND VPWR VPWR mem_rdata_q\[28\] sky130_fd_sc_hd__dfxtp_2
X_08691_ net115 net83 VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__nor2_1
X_17889_ clknet_leaf_92_clk _01058_ VGND VGND VPWR VPWR count_cycle\[34\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__14400__B _03378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12201__A _06223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16608__A _03039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09312_ cpu_state\[3\] cpu_state\[6\] _03410_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__nor3_2
XFILLER_0_87_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10462__A1 _04070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09243_ _03891_ _03862_ _03810_ _03867_ _03844_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__a32o_1
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15925__B1 _02623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12347__S _06652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14128__A _07778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09174_ _03864_ _03868_ _03781_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13400__A1 _07209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10375__B decoded_imm\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15153__A1 _01969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13164__A0 _06987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09368__C1 _04027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13178__S _07104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09907__A1 _04328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_149_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_149_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10073__S0 _04512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16489__S _02968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11190__A2 _05829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16653__A1 _06265_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08958_ cpuregs.regs\[20\]\[4\] cpuregs.regs\[21\]\[4\] cpuregs.regs\[22\]\[4\] cpuregs.regs\[23\]\[4\]
+ _03661_ _03662_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11478__B1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08889_ _00067_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_162_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14310__B _07986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10920_ _03618_ _05582_ _03617_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_86_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10851_ _04566_ _04532_ _05264_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__mux2_1
XANTENNA__14967__A1 _07679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08777__A_N net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13570_ _07420_ _07421_ _03275_ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_140_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_160_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10782_ _05434_ _05477_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__or2_2
XFILLER_0_137_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12521_ _06746_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12257__S _06604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18733__A net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15240_ _01984_ _02090_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__or2_1
X_12452_ _06709_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_175_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11403_ _06009_ _06010_ _06011_ _03750_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__a31o_1
X_15171_ _02021_ _02024_ _01984_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__mux2_1
XANTENNA__11402__B1 _03867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12383_ _06672_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14122_ _07851_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11334_ reg_next_pc\[30\] _05928_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16341__A0 _06947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11397__A _03635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14053_ count_instr\[21\] _07801_ _07790_ VGND VGND VPWR VPWR _07804_ sky130_fd_sc_hd__o21ai_1
X_11265_ _05891_ _05894_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13004_ _07009_ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__clkbuf_8
X_10216_ cpuregs.regs\[0\]\[23\] cpuregs.regs\[1\]\[23\] cpuregs.regs\[2\]\[23\] cpuregs.regs\[3\]\[23\]
+ _04472_ _04473_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__mux4_1
X_11196_ _04251_ _05838_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__and2_1
XANTENNA__16399__S _02895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output248_A net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16644__A1 _06231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17812_ clknet_leaf_62_clk _00981_ VGND VGND VPWR VPWR reg_pc\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11505__A_N cpuregs.waddr\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12720__S _06847_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10147_ _04215_ _04861_ _04296_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13458__A1 _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14955_ net212 net181 _01846_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__mux2_1
X_17743_ clknet_leaf_94_clk _00912_ VGND VGND VPWR VPWR count_instr\[14\] sky130_fd_sc_hd__dfxtp_1
X_10078_ _04793_ _04794_ _04575_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13906_ _07701_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__clkbuf_1
X_14886_ instr_sra instr_srai VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__nor2_1
X_17674_ clknet_leaf_126_clk _00843_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16625_ cpuregs.regs\[1\]\[8\] _06156_ _03040_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__mux2_1
X_13837_ cpuregs.regs\[0\]\[15\] VGND VGND VPWR VPWR _07658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10119__S1 _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_128_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16556_ _03012_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13768_ net86 decoded_imm\[27\] _07606_ VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13630__B2 _07217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09330__A _04064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15507_ cpuregs.regs\[0\]\[24\] cpuregs.regs\[1\]\[24\] cpuregs.regs\[2\]\[24\] cpuregs.regs\[3\]\[24\]
+ _02013_ _02014_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__mux4_1
X_12719_ _06852_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16487_ cpuregs.regs\[17\]\[7\] _06548_ _02968_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_13699_ net82 decoded_imm\[23\] VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18226_ clknet_leaf_104_clk _01297_ VGND VGND VPWR VPWR instr_timer sky130_fd_sc_hd__dfxtp_4
X_15438_ cpuregs.regs\[28\]\[20\] cpuregs.regs\[29\]\[20\] cpuregs.regs\[30\]\[20\]
+ cpuregs.regs\[31\]\[20\] _02030_ _02031_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18157_ clknet_leaf_72_clk alu_out\[31\] VGND VGND VPWR VPWR alu_out_q\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12736__A3 _06053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15369_ _02211_ _02212_ _02002_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__mux2_1
XANTENNA__09062__A1 mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10747__A2 _05367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16332__A0 _07007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17108_ clknet_leaf_112_clk _00282_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_471 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18088_ clknet_leaf_102_clk _01192_ VGND VGND VPWR VPWR timer\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09930_ cpuregs.regs\[4\]\[15\] cpuregs.regs\[5\]\[15\] cpuregs.regs\[6\]\[15\] cpuregs.regs\[7\]\[15\]
+ _04232_ _04233_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__mux4_1
X_17039_ clknet_leaf_124_clk _00213_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10055__S0 _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09861_ _04369_ _04583_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11172__A2 _05254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ net113 net81 VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__and2b_1
XANTENNA__12630__S _06799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09792_ _04272_ _04510_ _04516_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10380__B1 instr_rdinstr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14411__A _07998_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08743_ net129 net97 VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__or2_2
XANTENNA__09748__S0 _04472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09505__A _00073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10150__S _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08674_ net119 net87 VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_970 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14949__A1 net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15297__S1 _02075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10435__A1 _04010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11632__A0 _06193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16772__S _03127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10986__A2 _05398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09226_ _03957_ _03749_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__or2b_1
XANTENNA__15374__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15896__B _03940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15388__S _02110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09157_ mem_rdata_q\[16\] _03910_ _03846_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12805__S _06891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10294__S0 _04325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09088_ _03842_ _03737_ _03845_ _03847_ _03848_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_169_Right_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15221__S1 _01997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13688__A1 _04945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11050_ _05514_ _05700_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__nor2_1
XANTENNA__10046__S0 _04472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10001_ _03384_ _04718_ _04719_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__and3_1
XANTENNA__15417__A _03666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14637__B1 _08232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09415__A _03301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11156__S _04668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18728__A net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10349__S1 _04208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ count_cycle\[16\] _08365_ count_cycle\[17\] VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__a21o_1
X_11952_ _06427_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10903_ _05399_ _05591_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__and2_1
XANTENNA__15288__S1 _01974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14671_ _08309_ _08315_ _08318_ VGND VGND VPWR VPWR _08319_ sky130_fd_sc_hd__a21oi_1
X_11883_ _06390_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16410_ _02935_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__clkbuf_1
X_13622_ _07281_ _04777_ _07282_ reg_pc\[18\] VGND VGND VPWR VPWR _07471_ sky130_fd_sc_hd__a22o_1
X_10834_ net69 net68 net98 _03510_ _05236_ _05309_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__mux4_1
X_17390_ clknet_leaf_140_clk _00559_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16341_ _06947_ cpuregs.regs\[16\]\[2\] _02896_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__mux2_1
X_13553_ net71 decoded_imm\[13\] VGND VGND VPWR VPWR _07407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10765_ _03613_ _05221_ _05215_ _03615_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09292__A1 _04010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14991__A _03240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12504_ _06257_ cpuregs.regs\[28\]\[20\] _06737_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16272_ _06947_ cpuregs.regs\[15\]\[2\] _02859_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__mux2_1
X_13484_ _07191_ _07341_ _07342_ VGND VGND VPWR VPWR _07343_ sky130_fd_sc_hd__o21a_1
X_10696_ _05234_ _05267_ _05241_ _05233_ _05395_ _05287_ VGND VGND VPWR VPWR _05396_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13376__A0 _04040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output198_A net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18011_ clknet_leaf_79_clk _01148_ VGND VGND VPWR VPWR irq_mask\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15298__S _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15223_ _01937_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__buf_6
XFILLER_0_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12435_ cpuregs.regs\[27\]\[20\] _06575_ _06700_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15154_ _01933_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12366_ cpuregs.regs\[26\]\[20\] _06575_ _06663_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14105_ count_instr\[38\] count_instr\[37\] count_instr\[36\] VGND VGND VPWR VPWR
+ _07839_ sky130_fd_sc_hd__and3_1
XANTENNA__15668__A2 _02486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11317_ reg_next_pc\[27\] reg_out\[27\] _05928_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__mux2_2
XANTENNA__15212__S1 _01980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09309__B decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15085_ _01942_ _01943_ _03713_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__mux2_1
X_12297_ cpuregs.regs\[25\]\[20\] _06575_ _06626_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__mux2_1
XANTENNA__14876__B1 _07675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output75_A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14036_ count_instr\[16\] count_instr\[15\] _07787_ VGND VGND VPWR VPWR _07792_ sky130_fd_sc_hd__and3_1
X_11248_ reg_next_pc\[14\] reg_out\[14\] _05876_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__mux2_2
XFILLER_0_129_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09978__S0 _04487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16617__A1 _06124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11179_ net123 _04710_ _05824_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__a21o_2
XANTENNA__09325__A _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16093__A2 _03636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15987_ _03767_ _03788_ _03864_ _03880_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__a22o_1
XANTENNA__13300__A0 _06987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17726_ clknet_leaf_82_clk _00895_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14938_ net204 net173 _01835_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17657_ clknet_leaf_71_clk _00826_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_159_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14869_ count_cycle\[58\] _01798_ _01714_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__a21oi_1
XANTENNA__16158__A _02770_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13281__S _07165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15062__A _03666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16608_ _03039_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__buf_6
X_17588_ clknet_leaf_152_clk _00757_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16539_ _06080_ _02894_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__nand2_4
XFILLER_0_161_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09283__B2 _04014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13367__B1 _07210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12321__B_N cpuregs.waddr\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09011_ _03771_ _03772_ _03231_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18209_ clknet_leaf_39_clk _01280_ VGND VGND VPWR VPWR instr_slt sky130_fd_sc_hd__dfxtp_1
XANTENNA__15451__S1 _01997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16305__A0 _06980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10653__B net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08404__A reg_next_pc\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14867__B1 _07675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09913_ _04017_ count_cycle\[46\] _03252_ _04634_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__a211o_1
XFILLER_0_112_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_694 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11145__A2 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11765__A _06311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09844_ _04420_ _04567_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__or2_1
XANTENNA__15237__A _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16084__A2 _03935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ irq_pending\[10\] _04049_ _04465_ _03385_ _04500_ VGND VGND VPWR VPWR _08370_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__16767__S _03116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13980__A _07737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08726_ net104 net72 VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09510__A2 _04021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08657_ timer\[29\] timer\[28\] timer\[30\] VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__or3_1
XANTENNA__08944__S1 _03643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14398__A2 _07947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08588_ instr_waitirq decoder_trigger VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__or2b_2
XFILLER_0_49_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11605__B1 _06098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10959__A2 _04744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_1006 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15700__A _01881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10550_ _05226_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09209_ mem_rdata_q\[11\] _03763_ _03951_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10481_ _05184_ _05185_ _04223_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__mux2_1
XANTENNA__12535__S _06752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12220_ _06273_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12581__A1 _06584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12151_ cpuregs.waddr\[1\] cpuregs.waddr\[0\] _06532_ VGND VGND VPWR VPWR _06533_
+ sky130_fd_sc_hd__nor3_4
XANTENNA__14858__B1 _01723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11102_ _05776_ _05713_ _05413_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__mux2_1
X_12082_ _06495_ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__buf_6
XANTENNA__11675__A _06231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11033_ _05481_ _05621_ _05707_ _05712_ VGND VGND VPWR VPWR alu_out\[24\] sky130_fd_sc_hd__a211o_1
X_15910_ instr_slli _02635_ _02648_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__a21o_1
XANTENNA__15147__A _03653_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16890_ clknet_leaf_33_clk _00060_ VGND VGND VPWR VPWR mem_rdata_q\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11394__B _06003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15841_ _03634_ _02602_ _02603_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__and3_1
XANTENNA__16677__S _03076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14986__A _01872_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12097__A0 _06150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18560_ clknet_leaf_157_clk _01625_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15772_ _05139_ _02486_ _02566_ _02545_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__o211a_1
X_12984_ cpuregs.regs\[3\]\[0\] _06531_ _07010_ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17511_ clknet_leaf_178_clk _00680_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11844__A0 _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14723_ _08356_ _08350_ _08357_ VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__and3b_1
XANTENNA__08935__S1 _03659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11935_ _06417_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output113_A net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18491_ clknet_leaf_181_clk _01556_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17442_ clknet_leaf_188_clk _00611_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_14654_ _08303_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__clkbuf_1
X_11866_ _06379_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13605_ _07452_ _07454_ _07455_ _07283_ VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__o22a_1
X_10817_ _05510_ _05479_ _05235_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17373_ clknet_leaf_163_clk _00542_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14585_ _08212_ _07958_ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__or2_1
X_11797_ reg_out\[31\] alu_out_q\[31\] _06069_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13536_ _07190_ _07388_ _07390_ VGND VGND VPWR VPWR _07391_ sky130_fd_sc_hd__or3_1
XFILLER_0_137_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16324_ _06999_ cpuregs.regs\[15\]\[27\] _02881_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__mux2_1
X_10748_ _03520_ _05440_ _05400_ _05444_ _05445_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__o221a_1
XFILLER_0_153_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_615 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15433__S1 _02086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16255_ mem_rdata_q\[4\] _03885_ _03914_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__mux2_1
XANTENNA__15889__A2 _02635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13467_ _07310_ VGND VGND VPWR VPWR _07327_ sky130_fd_sc_hd__inv_2
XANTENNA__12445__S _06700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10679_ _05308_ _05312_ _05239_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12021__A0 _06114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15206_ _01959_ _02050_ _02058_ _01933_ decoded_imm\[7\] VGND VGND VPWR VPWR _02059_
+ sky130_fd_sc_hd__a32o_1
X_12418_ cpuregs.regs\[27\]\[12\] _06559_ _06689_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__mux2_1
X_16186_ _02811_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14561__A2 _07954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13398_ _07259_ _07260_ _07261_ VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__nand3_1
Xoutput206 net206 VGND VGND VPWR VPWR mem_la_addr[22] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput217 net217 VGND VGND VPWR VPWR mem_la_addr[3] sky130_fd_sc_hd__buf_1
X_15137_ _01991_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__buf_8
XFILLER_0_105_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput228 net228 VGND VGND VPWR VPWR mem_la_wdata[12] sky130_fd_sc_hd__buf_1
X_12349_ cpuregs.regs\[26\]\[12\] _06559_ _06652_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__mux2_1
Xoutput239 net239 VGND VGND VPWR VPWR mem_la_wdata[22] sky130_fd_sc_hd__buf_1
XFILLER_0_121_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14849__B1 _01723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15068_ _01913_ _01917_ _01923_ _01927_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__o22a_1
XANTENNA__14313__A2 _07988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14019_ _07780_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12180__S _06534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16066__A2 _08232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16587__S _03026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15491__S _03713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10904__A2_N _05301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09560_ _04290_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08894__A _00065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08511_ _03293_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__buf_4
X_17709_ clknet_leaf_75_clk _00878_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09491_ _04222_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__buf_6
XANTENNA__08926__S1 _03659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11524__S _06086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08442_ _03225_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_65_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09256__A1 _03994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10271__C1 _04982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12355__S _06652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11479__B _03428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15188__S0 _03670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11118__A2 _05221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14302__C irq_pending\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09827_ _04549_ _04550_ _04222_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09758_ cpuregs.regs\[4\]\[10\] cpuregs.regs\[5\]\[10\] cpuregs.regs\[6\]\[10\] cpuregs.regs\[7\]\[10\]
+ _04232_ _04233_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__mux4_1
XANTENNA__15360__S0 _02022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08709_ net77 VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__inv_2
X_09689_ _04271_ _04415_ _04416_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_159_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _06252_ _03320_ _06253_ _06271_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_159_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15032__A3 _05009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11651_ reg_pc\[15\] reg_pc\[14\] _06195_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__and3_1
XFILLER_0_167_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10602_ net77 net79 _05263_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11054__A1 _05277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10488__S0 _04325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14370_ _08024_ _08028_ _08040_ _08042_ VGND VGND VPWR VPWR _08043_ sky130_fd_sc_hd__a31o_1
X_11582_ _06145_ _06148_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__nor2_2
XFILLER_0_37_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13321_ _07188_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10533_ _05236_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12265__S _06604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12003__A0 _06312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16040_ _02715_ decoded_imm_j\[9\] _02726_ mem_rdata_q\[29\] _02634_ VGND VGND VPWR
+ VPWR _02732_ sky130_fd_sc_hd__a221o_1
X_13252_ _07007_ cpuregs.regs\[8\]\[31\] _07117_ VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__mux2_1
X_10464_ _05169_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__inv_2
XANTENNA__15740__A1 _04871_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11389__B _03994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12203_ _06568_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10565__A0 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13183_ _07115_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16261__A _07737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10395_ _05101_ _05102_ _04077_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12134_ _06523_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17991_ clknet_leaf_104_clk _01128_ VGND VGND VPWR VPWR irq_mask\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08698__B net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13096__S _07068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12065_ _06289_ cpuregs.regs\[22\]\[24\] _06482_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__mux2_1
X_16942_ clknet_leaf_119_clk _00123_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16048__A2 decoded_imm_j\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11016_ _05363_ _03473_ _05675_ _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__o31ai_1
XANTENNA__09722__A2 _04448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output230_A net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16873_ _06588_ cpuregs.regs\[14\]\[26\] _03174_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__mux2_1
X_18612_ clknet_leaf_117_clk _01677_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_15824_ _02595_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11817__A0 _06132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18543_ clknet_leaf_58_clk _01608_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_15755_ _05009_ _02486_ _02553_ _02545_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12967_ _06311_ VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__buf_2
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10096__A2 _04810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14706_ count_cycle\[4\] count_cycle\[5\] count_cycle\[6\] _08340_ VGND VGND VPWR
+ VPWR _08346_ sky130_fd_sc_hd__and4_2
X_11918_ _06408_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15559__A1 _02066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18474_ clknet_leaf_123_clk _01539_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12898_ _06952_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__clkbuf_1
X_15686_ _02477_ _02499_ _02501_ _02502_ _06026_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__o311a_1
XFILLER_0_157_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17425_ clknet_leaf_136_clk _00594_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14637_ _08268_ _07964_ _08232_ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__o21ai_2
X_11849_ _06257_ cpuregs.regs\[11\]\[20\] _06370_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12964__A _06303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15978__C mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09749__S _04430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17356_ clknet_leaf_147_clk _00525_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10479__S0 _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14568_ _08180_ _08189_ _08220_ _08224_ VGND VGND VPWR VPWR _08225_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_60_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08997__A0 mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12793__A1 _06580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16307_ _06982_ cpuregs.regs\[15\]\[19\] _02870_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__mux2_1
X_13519_ _07375_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__clkbuf_1
X_17287_ clknet_leaf_157_clk _00461_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14499_ _08160_ _08156_ VGND VGND VPWR VPWR _08161_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16238_ _02843_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09410__A1 irq_mask\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12903__S _06943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16169_ net278 net240 _02797_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__mux2_1
XANTENNA__09410__B2 _04024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08889__A _00067_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10020__A2 _04448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08991_ mem_la_secondword VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15495__A0 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12204__A _06231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15590__S0 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08871__A1_N _03630_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09174__B1 _03781_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16039__A2 _02711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09612_ net95 VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15342__S0 _02111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09513__A reg_pc\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09543_ _04273_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14470__A1 _07898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09474_ _04053_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09572__S1 _04219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_526 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08425_ _03209_ _03210_ _03203_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12784__A1 _06571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12085__S _06496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16780__S _03127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10795__B1 _05357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13733__B1 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08799__A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10180_ _04483_ _04893_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__nand2_1
XANTENNA__14289__A1 reg_pc\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14289__B2 _07960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15789__A1 _03385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13870_ _07674_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15789__B2 _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12821_ _06909_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09468__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09468__B2 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12752_ _06872_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12472__A0 _06132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15540_ cpuregs.regs\[24\]\[26\] cpuregs.regs\[25\]\[26\] cpuregs.regs\[26\]\[26\]
+ cpuregs.regs\[27\]\[26\] _03645_ _01991_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__mux4_1
XANTENNA__09563__S1 _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11703_ _06256_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__buf_2
XFILLER_0_139_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15471_ cpuregs.regs\[8\]\[22\] cpuregs.regs\[9\]\[22\] cpuregs.regs\[10\]\[22\]
+ cpuregs.regs\[11\]\[22\] _01999_ _02000_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__mux4_1
X_12683_ _06833_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17210_ clknet_leaf_188_clk _00384_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15160__A _03643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14422_ _08012_ _08089_ _08090_ VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11634_ reg_pc\[13\] _06187_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__and2_1
X_18190_ clknet_leaf_41_clk _01261_ VGND VGND VPWR VPWR instr_lb sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08979__A0 mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17141_ clknet_leaf_116_clk _00315_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_14353_ _08017_ _08023_ _08026_ VGND VGND VPWR VPWR _08027_ sky130_fd_sc_hd__or3_1
X_11565_ _06133_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13304_ _06991_ cpuregs.regs\[5\]\[23\] _07176_ VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__mux2_1
X_10516_ _05215_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17072_ clknet_leaf_164_clk _00246_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10250__A2 _04145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14284_ reg_next_pc\[27\] _05928_ _07944_ _07965_ VGND VGND VPWR VPWR _07966_ sky130_fd_sc_hd__o211a_2
XANTENNA__15713__A1 _04631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11496_ reg_out\[0\] alu_out_q\[0\] _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__mux2_1
XANTENNA_output180_A net180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13235_ _07143_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__clkbuf_1
X_16023_ mem_rdata_q\[23\] _02712_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__and2_1
X_10447_ cpuregs.regs\[20\]\[30\] cpuregs.regs\[21\]\[30\] cpuregs.regs\[22\]\[30\]
+ cpuregs.regs\[23\]\[30\] _04472_ _04473_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__mux4_1
XFILLER_0_150_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13166_ _06989_ cpuregs.regs\[4\]\[22\] _07104_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__mux2_1
X_10378_ net87 VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__buf_4
XANTENNA__08502__A _03239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15477__B1 _02313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12117_ _06514_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17974_ clknet_leaf_43_clk _01111_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dfxtp_2
XANTENNA__15572__S0 _01918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13097_ _07070_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__clkbuf_1
X_12048_ _06224_ cpuregs.regs\[22\]\[16\] _06471_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__mux2_1
X_16925_ clknet_leaf_115_clk _00106_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15229__B1 _02079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16856_ _06571_ cpuregs.regs\[14\]\[18\] _03163_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__mux2_1
XANTENNA__15324__S0 _01976_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15807_ _05960_ _05970_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__nor2_1
X_16787_ _03135_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16865__S _03174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14452__A1 _07898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13999_ _07765_ _07766_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18526_ clknet_leaf_175_clk _01591_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15738_ timer\[21\] _02538_ _02488_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_29_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18457_ clknet_leaf_1_clk _01522_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15669_ timer\[3\] timer\[2\] _02483_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__or3_1
XFILLER_0_158_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17408_ clknet_leaf_169_clk _00577_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_09190_ _03935_ _03938_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__or2_1
XANTENNA__13412__C1 _07274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18388_ clknet_leaf_168_clk _01453_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17339_ clknet_leaf_17_clk _00086_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10777__B1 _05357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15165__C1 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10529__A0 _04419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16105__S _03635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10153__S _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08974_ _03728_ _03732_ _03734_ _03735_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__a31oi_4
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09698__A1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09698__B2 _03225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10701__A0 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15315__S0 _02022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09793__S1 _04285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14979__C1 _08335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15640__B1 _03364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09526_ _04256_ _04248_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10465__C1 _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09457_ _04168_ _04186_ _04189_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__a21o_1
XANTENNA__15618__S1 _02047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08408_ irq_state\[1\] irq_state\[0\] VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__or2_1
XANTENNA__16334__B_N _06082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15943__A1 _04018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09388_ cpuregs.regs\[20\]\[2\] cpuregs.regs\[21\]\[2\] cpuregs.regs\[22\]\[2\] cpuregs.regs\[23\]\[2\]
+ _04072_ _04074_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__mux4_1
XANTENNA__15943__B2 _02667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_778 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14308__B _07984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_812 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11350_ _03787_ _03762_ _03770_ _03736_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10301_ _04010_ _04992_ _05011_ _04150_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_130_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11281_ _04848_ _05907_ _05827_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__mux2_1
XANTENNA__12543__S _06752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13020_ _07029_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__clkbuf_1
X_10232_ net82 VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10163_ _04821_ _04824_ _04877_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_167_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16120__B2 _02771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15554__S0 _02085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14978__B _01865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10094_ _04668_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__buf_2
X_14971_ _01862_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09689__A1 _04271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14682__A1 _03195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08976__B _03237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16710_ _06976_ cpuregs.regs\[19\]\[16\] _03087_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__mux2_1
X_13922_ _07691_ _07712_ VGND VGND VPWR VPWR _07713_ sky130_fd_sc_hd__and2_1
XANTENNA__10299__A2 _04448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11496__A1 alu_out_q\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12693__A0 _06193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09784__S1 _04285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17690_ clknet_leaf_20_clk _00859_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16641_ _03057_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__clkbuf_1
X_13853_ cpuregs.regs\[0\]\[23\] VGND VGND VPWR VPWR _07666_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16685__S _03076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14434__A1 _07899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12804_ _06899_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__clkbuf_1
X_16572_ _06974_ cpuregs.regs\[18\]\[15\] _03015_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__mux2_1
X_10996_ _05675_ _05677_ _05323_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__mux2_1
X_13784_ _07620_ _07621_ VGND VGND VPWR VPWR _07622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18311_ clknet_leaf_35_clk _01379_ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15523_ cpuregs.regs\[12\]\[25\] cpuregs.regs\[13\]\[25\] cpuregs.regs\[14\]\[25\]
+ cpuregs.regs\[15\]\[25\] _02069_ _02070_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12735_ cpu_state\[3\] _06860_ VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12718__S _06847_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11622__S _06176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18242_ clknet_leaf_22_clk _01313_ VGND VGND VPWR VPWR decoded_imm\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12666_ _06383_ _06823_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__nand2_2
X_15454_ _02012_ _02292_ _02005_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11617_ reg_out\[11\] alu_out_q\[11\] _06067_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__mux2_1
X_14405_ _08072_ _08073_ _08060_ _08064_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_26_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18173_ clknet_leaf_24_clk _01244_ VGND VGND VPWR VPWR decoded_imm_j\[14\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_136_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09613__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15385_ _02226_ _02227_ _02110_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__mux2_1
X_12597_ _06080_ _06713_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__nand2_4
XFILLER_0_136_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17124_ clknet_leaf_143_clk _00298_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11548_ _06074_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__buf_2
X_14336_ _07972_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13549__S _07374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14267_ reg_pc\[21\] _07953_ _07954_ _07935_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__a22o_1
X_17055_ clknet_leaf_181_clk _00229_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12453__S _06700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11479_ irq_mask\[27\] _03428_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13218_ _07134_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__clkbuf_1
X_16006_ cpuregs.raddr2\[1\] _05974_ _05975_ _05978_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__a22o_1
XANTENNA__09916__A2 _04611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09328__A _00071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14198_ _07905_ VGND VGND VPWR VPWR _07906_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13149_ _06972_ cpuregs.regs\[4\]\[14\] _07093_ VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11296__C _05918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14888__B decoded_imm\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ clknet_leaf_191_clk _01094_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dfxtp_1
XANTENNA__13476__A2 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14673__A1 _07968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16908_ clknet_leaf_7_clk _00053_ VGND VGND VPWR VPWR mem_rdata_q\[27\] sky130_fd_sc_hd__dfxtp_4
X_08690_ _03454_ _03455_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__nor2_2
X_17888_ clknet_leaf_90_clk _01057_ VGND VGND VPWR VPWR count_cycle\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16839_ _03151_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__buf_6
XANTENNA__16595__S _03026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09311_ cpu_state\[3\] _04044_ _04045_ _04037_ _04046_ VGND VGND VPWR VPWR _04047_
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_24_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18509_ clknet_leaf_162_clk _01574_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12628__S _06799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09242_ _03749_ _03978_ _03982_ _03739_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_924 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10656__B _05357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09173_ _03781_ _03768_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__nor2_2
XANTENNA__08592__C_N _03364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09604__A1 _04289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13400__A2 _04186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11411__A1 _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11768__A reg_pc\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12363__S _06652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11487__B _03428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10073__S1 _04513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16102__A1 _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15536__S0 _02046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10922__B1 _05218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09672__S _04078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08957_ _03717_ _03718_ _03719_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__mux2_1
XANTENNA__13194__S _07118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11478__A1 _06054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08888_ _03652_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_162_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_162_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10850_ _03499_ _05357_ _05478_ _05540_ _05541_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10438__C1 _04202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16169__A1 net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09509_ _04240_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__inv_2
X_10781_ _05244_ _05334_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09843__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09843__B2 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14319__A _06860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12520_ _06320_ cpuregs.regs\[28\]\[28\] _06737_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09420__B decoded_imm\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12451_ cpuregs.regs\[27\]\[28\] _06592_ _06700_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11402_ _03844_ _03923_ _03867_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15170_ cpuregs.regs\[24\]\[6\] cpuregs.regs\[25\]\[6\] cpuregs.regs\[26\]\[6\] cpuregs.regs\[27\]\[6\]
+ _02022_ _02023_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12382_ cpuregs.regs\[26\]\[28\] _06592_ _06663_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_90 net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14121_ _07849_ _07815_ _07850_ VGND VGND VPWR VPWR _07851_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_169_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11333_ _05950_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__buf_2
XANTENNA__11678__A reg_pc\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12273__S _06604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14052_ count_instr\[21\] count_instr\[20\] _07799_ VGND VGND VPWR VPWR _07803_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11264_ reg_out\[17\] _05857_ _05893_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11166__B1 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13003_ _07020_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_37_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10215_ cpuregs.regs\[4\]\[23\] cpuregs.regs\[5\]\[23\] cpuregs.regs\[6\]\[23\] cpuregs.regs\[7\]\[23\]
+ _04472_ _04473_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__mux4_1
X_11195_ _03841_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__buf_4
XANTENNA__08987__A _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17811_ clknet_leaf_62_clk _00980_ VGND VGND VPWR VPWR reg_pc\[19\] sky130_fd_sc_hd__dfxtp_2
X_10146_ _04859_ _04860_ _04211_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__mux2_1
XANTENNA__13458__A2 _05227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17742_ clknet_leaf_95_clk _00911_ VGND VGND VPWR VPWR count_instr\[13\] sky130_fd_sc_hd__dfxtp_1
X_14954_ _01852_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__clkbuf_1
X_10077_ cpuregs.regs\[24\]\[19\] cpuregs.regs\[25\]\[19\] cpuregs.regs\[26\]\[19\]
+ cpuregs.regs\[27\]\[19\] _04579_ _04284_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13905_ _07691_ _07700_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17673_ clknet_leaf_176_clk _00842_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_14885_ count_cycle\[63\] _01807_ _01810_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__o21a_1
XFILLER_0_159_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16624_ _03048_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13836_ _07657_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16555_ _06957_ cpuregs.regs\[18\]\[7\] _03004_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__mux2_1
X_10979_ _03465_ _05651_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__and2_1
X_13767_ net86 decoded_imm\[27\] decoded_imm\[26\] net85 VGND VGND VPWR VPWR _07606_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15506_ _01984_ _02341_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12718_ _06289_ cpuregs.regs\[12\]\[24\] _06847_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__mux2_1
X_16486_ _02975_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__clkbuf_1
X_13698_ net82 decoded_imm\[23\] VGND VGND VPWR VPWR _07542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18225_ clknet_leaf_29_clk _01296_ VGND VGND VPWR VPWR instr_waitirq sky130_fd_sc_hd__dfxtp_2
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15437_ _02275_ _02276_ _01907_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__mux2_1
X_12649_ _06289_ cpuregs.regs\[30\]\[24\] _06810_ VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_154_Left_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18156_ clknet_leaf_47_clk alu_out\[30\] VGND VGND VPWR VPWR alu_out_q\[30\] sky130_fd_sc_hd__dfxtp_1
X_15368_ cpuregs.regs\[0\]\[16\] cpuregs.regs\[1\]\[16\] cpuregs.regs\[2\]\[16\] cpuregs.regs\[3\]\[16\]
+ _01985_ _01986_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13279__S _07165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17107_ clknet_leaf_19_clk _00281_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18081__D _01186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14319_ _06860_ _07995_ VGND VGND VPWR VPWR _07996_ sky130_fd_sc_hd__nor2_1
X_18087_ clknet_leaf_102_clk _01191_ VGND VGND VPWR VPWR timer\[2\] sky130_fd_sc_hd__dfxtp_1
X_15299_ _02141_ _02143_ _02146_ _02088_ _02018_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17038_ clknet_leaf_123_clk _00212_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09445__S0 _04084_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09860_ cpuregs.regs\[0\]\[13\] cpuregs.regs\[1\]\[13\] cpuregs.regs\[2\]\[13\] cpuregs.regs\[3\]\[13\]
+ _04487_ _04469_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__mux4_1
XANTENNA__10055__S1 _04478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15518__S0 _01973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10904__B1 _05356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08897__A _00065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09492__S _04223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08811_ _03573_ net79 _03574_ _03576_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__a31o_1
XANTENNA__09770__B1 instr_rdinstr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09791_ _04289_ _04515_ _04296_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_163_Left_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14646__A1 _08232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08742_ _03507_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__inv_2
XANTENNA__12657__A0 _06320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09748__S1 _04473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08673_ _03434_ _03438_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_186_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_186_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_1015 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_982 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09521__A _04036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_172_Left_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09225_ _03959_ _03966_ _03960_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12882__A _06077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09156_ _03849_ _03201_ _03202_ _03850_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12093__S _06496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09087_ _03783_ _03748_ _03835_ _03844_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_142_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10294__S1 _04277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_110_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11148__A0 _05324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09436__S0 _04056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10046__S1 _04473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15509__S0 _02022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_164_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10000_ _04716_ _04717_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__or2_1
XANTENNA__10371__A1 _04391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09989_ _03225_ _04672_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_125_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11320__A0 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_177_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_177_clk sky130_fd_sc_hd__clkbuf_2
X_11951_ _06105_ cpuregs.regs\[21\]\[2\] _06424_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__mux2_1
XANTENNA__11383__D _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10902_ _05461_ _05590_ _05244_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__mux2_1
X_11882_ _06105_ cpuregs.regs\[20\]\[2\] _06387_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14670_ _08316_ _08317_ VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13621_ _07470_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__clkbuf_1
X_10833_ _03501_ _05440_ _05522_ _03503_ _05525_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__o221a_1
XFILLER_0_168_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11680__B _06118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16340_ _02898_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12820__A0 _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13552_ net71 decoded_imm\[13\] VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__or2_1
X_10764_ _05460_ _05376_ _05242_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12503_ _06714_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__buf_6
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13483_ _07281_ _04415_ _07282_ reg_pc\[8\] _07284_ VGND VGND VPWR VPWR _07342_ sky130_fd_sc_hd__a221o_1
X_16271_ _02861_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10695_ _05246_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__16264__A reg_next_pc\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18010_ clknet_leaf_78_clk _01147_ VGND VGND VPWR VPWR irq_mask\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15222_ _01995_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__buf_8
X_12434_ _06677_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12365_ _06640_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__clkbuf_8
X_15153_ _01969_ _01983_ _02007_ _01960_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_101_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_101_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_91_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11316_ _05936_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_2
X_14104_ count_instr\[37\] _07836_ _07838_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__a21oi_1
X_15084_ cpuregs.regs\[0\]\[1\] cpuregs.regs\[1\]\[1\] cpuregs.regs\[2\]\[1\] cpuregs.regs\[3\]\[1\]
+ _03669_ _03646_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__mux4_1
XANTENNA_output260_A net260 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12296_ _06603_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__clkbuf_8
X_14035_ _07789_ _07791_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__nor2_1
X_11247_ _05829_ _05878_ _05879_ _05880_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__a31o_4
XTAP_TAPCELL_ROW_52_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09978__S1 _04469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output68_A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09606__A _04051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11178_ _04038_ net128 net105 _03297_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__a22o_1
XANTENNA__08510__A _03292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10362__B2 _04187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10129_ count_instr\[52\] _04104_ _04105_ count_cycle\[52\] VGND VGND VPWR VPWR _04845_
+ sky130_fd_sc_hd__a22o_1
X_15986_ _05990_ _02701_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17725_ clknet_leaf_83_clk _00894_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dfxtp_1
XANTENNA__11311__A0 reg_next_pc\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14937_ _01843_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_168_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_168_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__12967__A _06311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17656_ clknet_leaf_48_clk _00825_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfxtp_2
X_14868_ _01798_ _01799_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15053__A1 _01907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16607_ _06750_ cpuregs.waddr\[1\] cpuregs.waddr\[0\] VGND VGND VPWR VPWR _03039_
+ sky130_fd_sc_hd__nor3b_4
XFILLER_0_86_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13819_ cpuregs.regs\[0\]\[6\] VGND VGND VPWR VPWR _07649_ sky130_fd_sc_hd__clkbuf_1
X_17587_ clknet_leaf_153_clk _00756_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16873__S _03174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14799_ _03304_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16538_ _03002_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09283__A2 _04012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11090__A2 _05398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09995__B decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12906__S _06943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16469_ _07007_ cpuregs.regs\[29\]\[31\] _02931_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09010_ net34 mem_rdata_q\[10\] _03729_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__mux2_1
X_18208_ clknet_leaf_41_clk _01279_ VGND VGND VPWR VPWR instr_sll sky130_fd_sc_hd__dfxtp_2
XFILLER_0_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18139_ clknet_leaf_71_clk alu_out\[13\] VGND VGND VPWR VPWR alu_out_q\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15108__A2 _03703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12207__A _06239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09912_ count_instr\[46\] instr_rdinstrh instr_rdinstr count_instr\[14\] VGND VGND
+ VPWR VPWR _04634_ sky130_fd_sc_hd__a22o_1
XANTENNA__10519__A2_N _05221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12878__A0 _06336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12641__S _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09843_ net53 _04030_ _04034_ net36 _04423_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__o221a_1
X_09774_ _03638_ _04466_ _04468_ _03226_ _04499_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ net104 net72 VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_159_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_159_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_87_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_174_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ timer\[8\] _03417_ _03421_ _03422_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__or4_1
XANTENNA__16241__A0 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08587_ instr_jal VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_189_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10959__A3 _04708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15700__B _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_1018 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12816__S _06906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09208_ _03952_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10480_ cpuregs.regs\[16\]\[31\] cpuregs.regs\[17\]\[31\] cpuregs.regs\[18\]\[31\]
+ cpuregs.regs\[19\]\[31\] _04291_ _04292_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__mux4_1
XFILLER_0_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14316__B _07983_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09139_ _03883_ _03894_ _03895_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_118_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09982__B1 _04100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12150_ cpuregs.waddr\[2\] _06081_ _06082_ _06083_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_20_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11101_ _05143_ _05086_ _05076_ _05044_ _05324_ _05286_ VGND VGND VPWR VPWR _05776_
+ sky130_fd_sc_hd__mux4_1
X_12081_ _06346_ _06385_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__nand2_4
XANTENNA_clkbuf_leaf_127_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11032_ _05219_ _05711_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__nor2_1
XANTENNA__13530__A1 _03276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09426__A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15840_ _03215_ _03979_ _03864_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__and3_1
XANTENNA__15283__B2 _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15771_ timer\[29\] _02561_ _02565_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__a21o_1
X_12983_ _07009_ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__buf_6
XFILLER_0_19_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17510_ clknet_leaf_18_clk _00679_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14722_ count_cycle\[10\] _08353_ count_cycle\[11\] VGND VGND VPWR VPWR _08357_ sky130_fd_sc_hd__a21o_1
XANTENNA__15163__A _03674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18490_ clknet_leaf_171_clk _01555_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11934_ _06312_ cpuregs.regs\[20\]\[27\] _06409_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17441_ clknet_leaf_15_clk _00610_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14653_ _08298_ _08299_ _08302_ VGND VGND VPWR VPWR _08303_ sky130_fd_sc_hd__or3b_1
XANTENNA__16693__S _03076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11865_ _06320_ cpuregs.regs\[11\]\[28\] _06370_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__mux2_1
XANTENNA_output106_A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13604_ _03387_ _04702_ _07210_ reg_pc\[16\] VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__a2bb2o_1
X_10816_ net68 net98 _05229_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__mux2_1
X_17372_ clknet_leaf_163_clk _00541_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_11796_ reg_pc\[31\] _06330_ _06338_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__a21oi_1
X_14584_ _08212_ _07958_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09896__S0 _04216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16323_ _02888_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11072__A2 _05397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13535_ _04419_ _07315_ _07389_ _07216_ VGND VGND VPWR VPWR _07390_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_31_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10747_ _03519_ _05367_ _05356_ _03522_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__o22a_1
XANTENNA__12726__S _06847_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10280__B1 _04105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14546__B1 _07997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16254_ _02851_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__clkbuf_1
X_10678_ _05305_ _05307_ _05239_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__mux2_1
X_13466_ _04360_ decoded_imm\[7\] VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__nor2_1
XANTENNA__09648__S0 _04216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15205_ _02005_ _02053_ _02057_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__a21o_1
X_12417_ _06691_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__clkbuf_1
X_16185_ net287 net249 _02770_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__mux2_1
X_13397_ _07244_ _07246_ _07243_ VGND VGND VPWR VPWR _07261_ sky130_fd_sc_hd__a21bo_1
XANTENNA__16299__A0 _06974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput207 net207 VGND VGND VPWR VPWR mem_la_addr[23] sky130_fd_sc_hd__clkbuf_1
Xoutput218 net218 VGND VGND VPWR VPWR mem_la_addr[4] sky130_fd_sc_hd__clkbuf_1
XANTENNA__09973__B1 _04082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15136_ _03642_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__buf_6
Xoutput229 net229 VGND VGND VPWR VPWR mem_la_wdata[13] sky130_fd_sc_hd__clkbuf_1
X_12348_ _06654_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13557__S _05227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10770__A net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12279_ _06617_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__clkbuf_1
X_15067_ _03657_ _01926_ _03675_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__a21o_1
X_14018_ _07777_ _07778_ _07779_ VGND VGND VPWR VPWR _07780_ sky130_fd_sc_hd__and3b_1
XANTENNA__10335__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10886__A2 _05398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15969_ _04168_ _03636_ _06003_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08510_ _03292_ _03196_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__nor2_4
XFILLER_0_172_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17708_ clknet_leaf_76_clk _00877_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dfxtp_1
XANTENNA__15073__A _01932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09490_ _04063_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__buf_6
XFILLER_0_78_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16223__A0 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08441_ cpu_state\[6\] VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__clkbuf_4
X_17639_ clknet_leaf_51_clk _00808_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_65_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13588__A1 _07217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_985 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12636__S _06799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09639__S0 _04290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10023__B1 _04009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15188__S1 _03671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13512__A1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10326__A1 _04052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16778__S _03127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14302__D irq_pending\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09826_ cpuregs.regs\[0\]\[12\] cpuregs.regs\[1\]\[12\] cpuregs.regs\[2\]\[12\] cpuregs.regs\[3\]\[12\]
+ _04216_ _04376_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__mux4_1
XANTENNA__09680__S _04078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09757_ _04069_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__buf_4
XANTENNA__15360__S1 _02023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08708_ _03463_ _03466_ _03469_ _03473_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__or4_1
X_09688_ irq_mask\[8\] _04308_ timer\[8\] _04023_ _04026_ VGND VGND VPWR VPWR _04416_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__10185__S0 _04056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _03258_ _03291_ _03287_ instr_sb VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11650_ _06209_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10601_ _04744_ net76 _05229_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16517__A1 _06578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11581_ _06146_ _06147_ _06075_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__o21a_1
XFILLER_0_153_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10488__S1 _04277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10532_ _03609_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__clkbuf_4
X_13320_ _07007_ cpuregs.regs\[5\]\[31\] _07153_ VGND VGND VPWR VPWR _07188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15725__C1 _06026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10463_ _05156_ _05160_ net300 _05168_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__a211o_2
X_13251_ _07151_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11389__C _04000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12202_ cpuregs.regs\[24\]\[16\] _06567_ _06555_ VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__mux2_1
X_13182_ _07005_ cpuregs.regs\[4\]\[30\] _07081_ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__mux2_1
X_10394_ cpuregs.regs\[8\]\[28\] cpuregs.regs\[9\]\[28\] cpuregs.regs\[10\]\[28\]
+ cpuregs.regs\[11\]\[28\] _04123_ _04124_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__mux4_1
XANTENNA__10565__A1 _04945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12133_ _06289_ cpuregs.regs\[23\]\[24\] _06518_ VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15158__A _03653_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17990_ clknet_leaf_105_clk _01127_ VGND VGND VPWR VPWR irq_mask\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09707__B1 _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14700__B1 _07826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12064_ _06486_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__clkbuf_1
X_16941_ clknet_leaf_105_clk _00122_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__14997__A _04493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11015_ _05323_ _03470_ _05677_ _05695_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__a31o_1
X_16872_ _03180_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08995__A _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16453__A0 _06991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08930__A1 _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18611_ clknet_leaf_113_clk _01676_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_15823_ decoded_imm_j\[12\] _03737_ _03635_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__mux2_1
XANTENNA_output223_A net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18542_ clknet_leaf_110_clk _01607_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15754_ _02476_ _02551_ _02552_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__or3b_1
X_12966_ _06998_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _08345_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__clkbuf_1
X_11917_ _06248_ cpuregs.regs\[20\]\[19\] _06398_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18473_ clknet_leaf_121_clk _01538_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15685_ _04382_ _02479_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__nand2_1
X_12897_ _06951_ cpuregs.regs\[31\]\[4\] _06943_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17424_ clknet_leaf_159_clk _00593_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14767__B1 _01717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14636_ _08221_ _07966_ VGND VGND VPWR VPWR _08287_ sky130_fd_sc_hd__xnor2_1
X_11848_ _06347_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17355_ clknet_leaf_139_clk _00524_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16508__A1 _06569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10479__S1 _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14567_ _08187_ _08199_ _08220_ _08223_ VGND VGND VPWR VPWR _08224_ sky130_fd_sc_hd__o31a_1
XFILLER_0_144_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11779_ _06322_ _06323_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16306_ _02879_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08997__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13518_ _04466_ _07373_ _07374_ VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17286_ clknet_leaf_136_clk _00460_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_14498_ _07941_ VGND VGND VPWR VPWR _08160_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16237_ net52 mem_16bit_buffer\[11\] _02830_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__mux2_1
XANTENNA__15192__B1 _00067_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13449_ net95 decoded_imm\[6\] VGND VGND VPWR VPWR _07310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16168_ _02802_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09410__A2 _04022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13287__S _07165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15119_ _01919_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__buf_8
XANTENNA__10704__S _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16099_ _03854_ _02760_ _02761_ _05993_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__o211a_1
X_08990_ mem_rdata_q\[31\] net57 _03227_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__mux2_1
XANTENNA__15495__A1 _02331_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15590__S1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09174__A1 _03864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10005__A _04483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15247__A1 _02020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09611_ _04336_ _04337_ _04340_ _04149_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__o211a_1
XANTENNA__15342__S1 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09513__B decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09542_ _04055_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__buf_8
XANTENNA__12220__A _06273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14470__A2 _07934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09473_ _04018_ count_cycle\[36\] _04165_ count_cycle\[4\] _04204_ VGND VGND VPWR
+ VPWR _04205_ sky130_fd_sc_hd__a221o_1
XANTENNA__13750__S _07224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_90_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__14758__B1 _01717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08424_ mem_rdata_q\[17\] net41 _03207_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12366__S _06663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12233__A1 _06588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13430__B1 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13051__A _07045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_835 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12890__A _06104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09675__S _00071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13733__A1 _07304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14930__A0 net200 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13733__B2 reg_pc\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16683__A0 _06949_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10950__A2_N _05397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15706__A _08335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16301__S _02870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08912__A1 _03639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09809_ irq_pending\[11\] _04049_ _04507_ _04533_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__a211o_1
XANTENNA__15789__A2 _03292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12820_ _06105_ cpuregs.regs\[6\]\[2\] _06906_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__mux2_1
XANTENNA__09468__A2 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11275__A2 _05899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12751_ cpuregs.regs\[9\]\[2\] _06538_ _06869_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09873__C1 _04150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_579 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_81_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_2
X_11702_ _06226_ reg_next_pc\[20\] _06251_ _06255_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__a211o_2
XANTENNA__15441__A _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15470_ _02066_ _02307_ _03692_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12682_ _06150_ cpuregs.regs\[12\]\[7\] _06825_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14421_ _07925_ _07988_ _08076_ VGND VGND VPWR VPWR _08090_ sky130_fd_sc_hd__and3_1
XFILLER_0_166_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11633_ _06194_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12224__A1 _06582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10585__A _05287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12276__S _06615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08979__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17140_ clknet_leaf_120_clk _00314_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14352_ _08024_ _08025_ VGND VGND VPWR VPWR _08026_ sky130_fd_sc_hd__and2_1
X_11564_ _06132_ cpuregs.regs\[10\]\[5\] _06086_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13303_ _07179_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__clkbuf_1
X_10515_ _05218_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__clkbuf_8
X_17071_ clknet_leaf_122_clk _00245_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11495_ _06068_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__buf_4
X_14283_ _05941_ _06309_ VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__or2_1
XANTENNA__15713__A2 _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09585__S _04223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16022_ _02611_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__clkbuf_4
X_10446_ count_instr\[30\] _04012_ count_cycle\[30\] _04013_ _05151_ VGND VGND VPWR
+ VPWR _05152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13234_ _06989_ cpuregs.regs\[8\]\[22\] _07140_ VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10377_ _05082_ _05083_ _04156_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__a21o_1
X_13165_ _07106_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15477__A1 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12116_ _06224_ cpuregs.regs\[23\]\[16\] _06507_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__mux2_1
X_17973_ clknet_leaf_44_clk _01110_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dfxtp_2
X_13096_ _06987_ cpuregs.regs\[7\]\[21\] _07068_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__mux2_1
XANTENNA__15572__S1 _01919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12047_ _06477_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__clkbuf_1
X_16924_ clknet_leaf_130_clk _00105_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15229__A1 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09614__A _04036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16855_ _03171_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15324__S1 _01977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15806_ decoded_imm_j\[4\] _06006_ _02585_ _05988_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__o22a_1
X_16786_ _06569_ cpuregs.regs\[13\]\[17\] _03127_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10149__S0 _04758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13998_ count_instr\[4\] _07763_ _07759_ VGND VGND VPWR VPWR _07766_ sky130_fd_sc_hd__o21ai_1
X_18525_ clknet_leaf_186_clk _01590_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_15737_ timer\[21\] _02538_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12949_ _06265_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_29_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_72_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_153_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15088__S0 _03669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18456_ clknet_leaf_11_clk _01521_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_15668_ _07250_ _02486_ _02487_ _02489_ _06026_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17407_ clknet_leaf_163_clk _00576_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12215__A1 _06575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14619_ _08267_ _08271_ VGND VGND VPWR VPWR _08272_ sky130_fd_sc_hd__or2_2
XANTENNA__15070__B _01929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18387_ clknet_leaf_163_clk _01452_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15599_ cpuregs.regs\[0\]\[30\] cpuregs.regs\[1\]\[30\] cpuregs.regs\[2\]\[30\] cpuregs.regs\[3\]\[30\]
+ _01908_ _01909_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17338_ clknet_leaf_17_clk _00085_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__dfxtp_2
XANTENNA__09092__A0 mem_rdata_q\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17269_ clknet_leaf_115_clk _00443_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10529__A1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08973_ mem_16bit_buffer\[12\] _03728_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__nor2_1
XANTENNA__16121__S _02771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09698__A2 _04419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10701__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15315__S1 _02023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13326__S0 _04758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15640__A1 _03379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09525_ _04245_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_63_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__15079__S0 _01936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16357__A _02895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15261__A _02110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09456_ irq_mask\[3\] _04021_ timer\[3\] _04187_ _04188_ VGND VGND VPWR VPWR _04189_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08407_ _03191_ _03192_ _03187_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__and3b_1
XFILLER_0_163_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09607__C1 _04188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09387_ _04077_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__buf_6
XANTENNA__15943__A2 _02650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13954__B2 net146 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10768__A1 _05255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11965__A0 _06166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10312__S0 _04084_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12824__S _06906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10300_ _04168_ _05009_ _05010_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15200__S _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15251__S0 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14903__A0 net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11280_ _05904_ _05906_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_130_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_991 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11717__B1 _06101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10231_ _04268_ _04923_ _04943_ _04149_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__o211a_1
XANTENNA__09386__B2 _04120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09418__B decoded_imm\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15459__A1 _02020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10162_ _04875_ _04876_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_167_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10940__A1 _05361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_58_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15554__S1 _02086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10093_ net77 VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__clkbuf_4
X_14970_ _03301_ _04448_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__nand2_1
XANTENNA__09689__A2 _04415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13921_ _03352_ _07704_ _07705_ net135 VGND VGND VPWR VPWR _07712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16640_ cpuregs.regs\[1\]\[15\] _06215_ _03051_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13852_ _07665_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12803_ cpuregs.regs\[9\]\[27\] _06590_ _06891_ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__mux2_1
X_16571_ _03020_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12445__A1 _06586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13783_ net88 decoded_imm\[29\] VGND VGND VPWR VPWR _07621_ sky130_fd_sc_hd__or2_1
X_10995_ _05676_ _03464_ _05662_ _03462_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__o31ai_2
Xclkbuf_leaf_54_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__11903__S _06398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18310_ clknet_leaf_35_clk _01378_ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dfxtp_1
X_15522_ _03687_ _02356_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__or2_1
X_12734_ _03298_ _03277_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_26_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_67_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18241_ clknet_leaf_16_clk _01312_ VGND VGND VPWR VPWR cpuregs.raddr2\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15395__B1 _00068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15453_ cpuregs.regs\[20\]\[21\] cpuregs.regs\[21\]\[21\] cpuregs.regs\[22\]\[21\]
+ cpuregs.regs\[23\]\[21\] _02069_ _02070_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__mux4_1
XFILLER_0_167_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12665_ _06081_ _06082_ _06384_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__and3b_2
XFILLER_0_155_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15490__S0 _03640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14404_ _08060_ _08064_ _08072_ _08073_ VGND VGND VPWR VPWR _08074_ sky130_fd_sc_hd__a211o_1
X_11616_ reg_pc\[11\] _06171_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__or2_1
X_18172_ clknet_leaf_24_clk _01243_ VGND VGND VPWR VPWR decoded_imm_j\[13\] sky130_fd_sc_hd__dfxtp_2
X_15384_ cpuregs.regs\[16\]\[17\] cpuregs.regs\[17\]\[17\] cpuregs.regs\[18\]\[17\]
+ cpuregs.regs\[19\]\[17\] _02221_ _02222_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__mux4_1
X_12596_ _06786_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17123_ clknet_leaf_134_clk _00297_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14335_ decoded_imm_j\[1\] _07902_ _08009_ VGND VGND VPWR VPWR _08011_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11420__A2 _03763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11547_ reg_out\[4\] alu_out_q\[4\] latched_stalu VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15698__A1 _07371_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17054_ clknet_leaf_172_clk _00228_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_output98_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14266_ _05909_ _06263_ _07942_ _05910_ VGND VGND VPWR VPWR _07954_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_94_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11478_ _06054_ irq_pending\[26\] _06058_ net19 VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09377__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16005_ cpuregs.raddr2\[0\] _06006_ _05968_ _05972_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__o22a_1
XANTENNA__09377__B2 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13217_ _06972_ cpuregs.regs\[8\]\[14\] _07129_ VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__mux2_1
X_10429_ _04069_ _05135_ _04095_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14197_ _07904_ VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13148_ _07097_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09129__A1 _03878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11874__A cpuregs.waddr\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17956_ clknet_leaf_191_clk _01093_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dfxtp_1
X_13079_ _06970_ cpuregs.regs\[7\]\[13\] _07057_ VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__mux2_1
X_16907_ clknet_leaf_7_clk _00052_ VGND VGND VPWR VPWR mem_rdata_q\[26\] sky130_fd_sc_hd__dfxtp_4
X_17887_ clknet_leaf_90_clk _01056_ VGND VGND VPWR VPWR count_cycle\[32\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11085__S _05363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16838_ _03162_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13633__A0 _04754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16769_ _06552_ cpuregs.regs\[13\]\[9\] _03116_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09837__C1 net300 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12909__S _06943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_2
X_09310_ _03312_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__buf_4
XANTENNA__15081__A _03713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11813__S _06348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18508_ clknet_leaf_109_clk _01573_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09241_ _03878_ _03844_ _03968_ _03981_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__a211o_1
XFILLER_0_158_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18439_ clknet_leaf_151_clk _01504_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15925__A2 _02617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12739__A2 _06863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09172_ mem_rdata_q\[12\] _03736_ _03757_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11947__A0 _06078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11411__A2 _06016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15233__S0 _01976_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09519__A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09368__A1 irq_mask\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09368__B2 _04024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14361__A1 _07960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11175__A1 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13983__B _07754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15536__S1 _02047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15310__B1 _02006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08956_ _03713_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10135__C1 _04850_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16786__S _03127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08887_ _00066_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_162_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_36_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__11723__S _06258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09508_ _04213_ _04226_ _04227_ _04239_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__a211o_4
XFILLER_0_78_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10780_ _05278_ _05475_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10989__A1 _05281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09439_ _04053_ _04171_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11024__A _05288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15472__S0 _02074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12450_ _06708_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11938__A0 _06328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11401_ _03770_ _05989_ _03867_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__or3b_1
XANTENNA__10863__A _05414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12554__S _06763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12381_ _06671_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_80 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10610__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15224__S0 _02074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14120_ count_instr\[41\] count_instr\[40\] _07843_ count_instr\[42\] VGND VGND VPWR
+ VPWR _07850_ sky130_fd_sc_hd__a31o_1
X_11332_ _05143_ _05949_ _03219_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14051_ _07801_ _07802_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__nor2_1
XANTENNA__10074__S _04321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11263_ reg_next_pc\[17\] _05876_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__or2_1
XANTENNA__11166__A1 _04038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11166__B2 _03297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13002_ cpuregs.regs\[3\]\[9\] _06552_ _07010_ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10214_ _04206_ _04926_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__nand2_1
X_11194_ _05831_ _05835_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15301__B1 _01963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15166__A _03639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10145_ cpuregs.regs\[0\]\[21\] cpuregs.regs\[1\]\[21\] cpuregs.regs\[2\]\[21\] cpuregs.regs\[3\]\[21\]
+ _04758_ _04759_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__mux4_1
X_17810_ clknet_leaf_61_clk _00979_ VGND VGND VPWR VPWR reg_pc\[18\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__14070__A _03304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17741_ clknet_leaf_94_clk _00910_ VGND VGND VPWR VPWR count_instr\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09164__A _03916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14953_ net211 net180 _01846_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__mux2_1
X_10076_ cpuregs.regs\[28\]\[19\] cpuregs.regs\[29\]\[19\] cpuregs.regs\[30\]\[19\]
+ cpuregs.regs\[31\]\[19\] _04579_ _04284_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__mux4_1
XANTENNA__10126__C1 _04227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13904_ _03359_ _07678_ _07682_ net161 VGND VGND VPWR VPWR _07700_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17672_ clknet_leaf_185_clk _00841_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_14884_ count_cycle\[63\] _01807_ _01714_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16801__A0 _06584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16623_ cpuregs.regs\[1\]\[7\] _06149_ _03040_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13835_ cpuregs.regs\[0\]\[14\] VGND VGND VPWR VPWR _07657_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_43_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10429__B1 _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_471 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16554_ _03011_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__clkbuf_1
X_13766_ _07568_ _07604_ _07603_ VGND VGND VPWR VPWR _07605_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10978_ _05225_ _05654_ _05655_ _05661_ VGND VGND VPWR VPWR alu_out\[20\] sky130_fd_sc_hd__a211o_1
XANTENNA__08508__A _03239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15505_ cpuregs.regs\[4\]\[24\] cpuregs.regs\[5\]\[24\] cpuregs.regs\[6\]\[24\] cpuregs.regs\[7\]\[24\]
+ _01990_ _01992_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__mux4_1
X_12717_ _06851_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__clkbuf_1
X_16485_ cpuregs.regs\[17\]\[6\] _06546_ _02968_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13697_ _07537_ _07539_ _07540_ _07284_ VGND VGND VPWR VPWR _07541_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13918__A1 _03357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18224_ clknet_leaf_65_clk _01295_ VGND VGND VPWR VPWR instr_maskirq sky130_fd_sc_hd__dfxtp_2
XANTENNA__15463__S0 _02030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15436_ cpuregs.regs\[16\]\[20\] cpuregs.regs\[17\]\[20\] cpuregs.regs\[18\]\[20\]
+ cpuregs.regs\[19\]\[20\] _01918_ _01919_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12648_ _06814_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18155_ clknet_leaf_46_clk alu_out\[29\] VGND VGND VPWR VPWR alu_out_q\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15367_ cpuregs.regs\[4\]\[16\] cpuregs.regs\[5\]\[16\] cpuregs.regs\[6\]\[16\] cpuregs.regs\[7\]\[16\]
+ _02022_ _02023_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__mux4_1
XANTENNA__12464__S _06715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12579_ cpuregs.regs\[2\]\[23\] _06582_ _06774_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__mux2_1
XANTENNA__10601__A0 _04744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15215__S0 _01985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17106_ clknet_leaf_111_clk _00280_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09339__A _04073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14318_ _07992_ _07994_ VGND VGND VPWR VPWR _07995_ sky130_fd_sc_hd__or2_2
X_18086_ clknet_leaf_102_clk _01190_ VGND VGND VPWR VPWR timer\[1\] sky130_fd_sc_hd__dfxtp_1
X_15298_ _02144_ _02145_ _02002_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17037_ clknet_leaf_120_clk _00211_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_14249_ reg_pc\[16\] _07926_ _07941_ _07935_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09445__S1 _04086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15518__S1 _01974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13295__S _07165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16096__A1 _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08810_ net112 _03575_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__nor2_1
XANTENNA__12106__A0 _06184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09790_ _04511_ _04514_ _04321_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__mux2_1
XANTENNA__10380__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14646__A2 _07966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08741_ _03505_ _03506_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__nor2b_2
X_17939_ clknet_leaf_68_clk _08379_ VGND VGND VPWR VPWR reg_out\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09522__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10668__B1 _05220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09522__B2 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08672_ _03437_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_105_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10667__B _05367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09224_ mem_rdata_q\[26\] _03965_ _03757_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__mux2_2
XANTENNA__16020__B2 mem_rdata_q\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12374__S _06663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09155_ _03909_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09086_ mem_rdata_q\[7\] _03822_ _03846_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15531__B1 _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11148__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09436__S1 _04091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09683__S _04064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15509__S1 _02023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09988_ net74 VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__14098__B1 _07834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14637__A2 _07964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08939_ _03679_ _03694_ _03702_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _06426_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10901_ _05589_ _05527_ _05242_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__mux2_1
XANTENNA__12549__S _06752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11881_ _06389_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13620_ _04744_ _07469_ _07374_ VGND VGND VPWR VPWR _07470_ sky130_fd_sc_hd__mux2_1
X_10832_ _05288_ _05381_ _05524_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14270__B1 _07956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13551_ _07281_ _04593_ _07282_ reg_pc\[13\] VGND VGND VPWR VPWR _07405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10763_ _03518_ net95 _03524_ net93 _05236_ _05309_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09858__S _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12502_ _06736_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09029__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16270_ _06945_ cpuregs.regs\[15\]\[1\] _02859_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13482_ _07274_ _07294_ _07339_ _07340_ VGND VGND VPWR VPWR _07341_ sky130_fd_sc_hd__a31o_1
X_10694_ _05270_ _05273_ _05276_ _05334_ _05277_ _05278_ VGND VGND VPWR VPWR _05394_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_152_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16264__B _07778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15221_ cpuregs.regs\[24\]\[8\] cpuregs.regs\[25\]\[8\] cpuregs.regs\[26\]\[8\] cpuregs.regs\[27\]\[8\]
+ _01996_ _01997_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__mux4_1
X_12433_ _06699_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14573__A1 _08012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12284__S _06615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15152_ _01988_ _01994_ _02003_ _02004_ _02006_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__a221o_1
X_12364_ _06662_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14103_ count_instr\[37\] _07836_ _07675_ VGND VGND VPWR VPWR _07838_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11315_ _05044_ _05838_ _05935_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__a21bo_1
X_15083_ cpuregs.regs\[4\]\[1\] cpuregs.regs\[5\]\[1\] cpuregs.regs\[6\]\[1\] cpuregs.regs\[7\]\[1\]
+ _03669_ _03646_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__mux4_1
XANTENNA__11139__A1 _04040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12295_ _06625_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14034_ count_instr\[15\] _07787_ _07790_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11246_ _04602_ _03841_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16078__A1 decoded_imm\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16078__B2 mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13409__A _04419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_690 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11177_ net122 _04710_ _05823_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__a21o_2
XANTENNA__09606__B _04335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10362__A2 _04448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08510__B _03196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10128_ _04168_ _04842_ _04843_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__a21o_1
X_15985_ _03228_ _02697_ _02700_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17724_ clknet_leaf_82_clk _00893_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dfxtp_1
X_10059_ _04776_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__inv_2
X_14936_ net203 net172 _01835_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17655_ clknet_leaf_72_clk _00824_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfxtp_4
X_14867_ count_cycle\[57\] _01795_ _07675_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16606_ _03038_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__clkbuf_1
X_13818_ _07648_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17586_ clknet_leaf_141_clk _00755_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__14261__B1 _07950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14798_ count_cycle\[34\] count_cycle\[35\] _01748_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16537_ cpuregs.regs\[17\]\[31\] _06598_ _02967_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__mux2_1
X_13749_ _03276_ _07581_ _07582_ _07589_ VGND VGND VPWR VPWR _07590_ sky130_fd_sc_hd__a31o_1
XANTENNA__12811__A1 _06598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12983__A _07009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16002__A1 _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15436__S0 _01918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16468_ _02965_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14013__B1 _07775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18207_ clknet_leaf_41_clk _01278_ VGND VGND VPWR VPWR instr_sub sky130_fd_sc_hd__dfxtp_2
X_15419_ cpuregs.regs\[20\]\[19\] cpuregs.regs\[21\]\[19\] cpuregs.regs\[22\]\[19\]
+ cpuregs.regs\[23\]\[19\] _03649_ _01991_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_947 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16399_ _07005_ cpuregs.regs\[16\]\[30\] _02895_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18138_ clknet_leaf_41_clk alu_out\[12\] VGND VGND VPWR VPWR alu_out_q\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18069_ clknet_leaf_73_clk _01174_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfxtp_4
XANTENNA__09991__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15513__B1 _02027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12922__S _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09911_ irq_mask\[14\] _04021_ timer\[14\] _04187_ _04188_ VGND VGND VPWR VPWR _04633_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08701__A net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16069__A1 decoded_imm\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16069__B2 mem_rdata_q\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09842_ net70 VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12223__A _06280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15816__A1 _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11550__A1 _06116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10984__S0 _05264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15816__B2 _03987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09773_ _04494_ _04495_ _04498_ _04149_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_107_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08724_ net73 net105 VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_87_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ timer\[9\] timer\[11\] timer\[10\] VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__or3_1
XANTENNA__15044__A2 _01865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09259__B1 _03737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _03298_ _03319_ _03364_ _03308_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14252__B1 _07943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09354__S0 _04085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11605__A2 _03333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12893__A _06113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14004__B1 _07759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09207_ mem_rdata_q\[10\] _03892_ _03951_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11369__A1 _03885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09138_ _03794_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__buf_4
XANTENNA__09431__B1 _04008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15504__B1 _02006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12832__S _06906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09069_ _03828_ _03830_ _03231_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__mux2_1
X_11100_ _05564_ _05602_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12080_ _06494_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10329__C1 _04027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08611__A _03277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11031_ _03459_ _05710_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09734__B2 _04460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15770_ _02484_ _02564_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__nand2_1
X_12982_ _06676_ _06750_ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__nor2_4
XFILLER_0_19_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14721_ count_cycle\[10\] count_cycle\[11\] _08353_ VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__and3_1
X_11933_ _06416_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17440_ clknet_leaf_170_clk _00609_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_14652_ _08300_ _08301_ _08121_ VGND VGND VPWR VPWR _08302_ sky130_fd_sc_hd__or3b_1
XFILLER_0_68_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11864_ _06378_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13603_ _07254_ _07412_ _07453_ _07189_ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__a31o_1
X_10815_ _03506_ _05440_ _05367_ _03505_ _05508_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17371_ clknet_leaf_128_clk _00540_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14583_ _08071_ _08234_ _08235_ _08238_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__a211o_1
XANTENNA__10100__B decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11795_ reg_pc\[31\] _06330_ _06101_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11911__S _06398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09896__S1 _04376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16322_ _06997_ cpuregs.regs\[15\]\[26\] _02881_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__mux2_1
X_13534_ _04708_ _07276_ VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10746_ _05443_ _05344_ _05246_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16253_ mem_rdata_q\[3\] _03810_ _03914_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__mux2_1
XANTENNA__14546__A1 _07898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13465_ _03518_ decoded_imm\[7\] VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10677_ _05228_ _05375_ _05377_ _05251_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09648__S1 _04376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15204_ _03654_ _02056_ _03675_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13754__C1 _07274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12416_ cpuregs.regs\[27\]\[11\] _06557_ _06689_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__mux2_1
X_16184_ _02810_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__clkbuf_1
X_13396_ net92 decoded_imm\[3\] VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput208 net208 VGND VGND VPWR VPWR mem_la_addr[24] sky130_fd_sc_hd__buf_1
XANTENNA__08776__A2 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09973__A1 _04070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15135_ _01936_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__buf_8
XFILLER_0_50_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12347_ cpuregs.regs\[26\]\[11\] _06557_ _06652_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput219 net219 VGND VGND VPWR VPWR mem_la_addr[5] sky130_fd_sc_hd__buf_1
XFILLER_0_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11780__A1 alu_out_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15066_ _01924_ _01925_ _03664_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12278_ cpuregs.regs\[25\]\[11\] _06557_ _06615_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__mux2_1
XANTENNA__10770__B net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14017_ count_instr\[9\] _07773_ count_instr\[10\] VGND VGND VPWR VPWR _07779_ sky130_fd_sc_hd__a21o_1
X_11229_ _05862_ _05864_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11532__B2 _06093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15968_ net262 _02684_ _02688_ _01821_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09352__A _04086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17707_ clknet_leaf_75_clk _00876_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09584__S0 _04217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14919_ net195 net164 _01824_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15899_ instr_slti _02618_ _02641_ _02643_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08440_ _03197_ VGND VGND VPWR VPWR clear_prefetched_high_word sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17638_ clknet_leaf_51_clk _00807_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_172_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17569_ clknet_leaf_17_clk _00738_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11821__S _06348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13602__A _04642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09498__S _04211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09661__B1 _04389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10271__A1 _03638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10271__B2 _04960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09639__S1 _04276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09413__B1 _04009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10023__A1 _04018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13512__A2 _05259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09825_ cpuregs.regs\[4\]\[12\] cpuregs.regs\[5\]\[12\] cpuregs.regs\[6\]\[12\] cpuregs.regs\[7\]\[12\]
+ _04216_ _04376_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__mux4_1
XANTENNA__11792__A _06335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09756_ _04070_ _04481_ _04082_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__a21oi_1
X_08707_ _03472_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12099__S _06496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09687_ _04414_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__inv_2
XANTENNA__10185__S1 _04091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08638_ mem_wordsize\[1\] VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13028__A1 _06578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11039__B1 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09327__S0 _04057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08569_ irq_mask\[17\] irq_pending\[17\] VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__and2b_2
XANTENNA__15973__B1 _02650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11731__S _06258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10600_ _04040_ _05286_ _05222_ _05299_ _05302_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__a311o_1
XANTENNA__15203__S _03666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11580_ reg_pc\[7\] _06137_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10531_ _05231_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_137_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11032__A _05219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13250_ _07005_ cpuregs.regs\[8\]\[30\] _07117_ VGND VGND VPWR VPWR _07151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10462_ _04070_ _05163_ _05167_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12201_ _06223_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_40_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09955__A1 irq_pending\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09955__B2 _03385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12562__S _06763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13181_ _07114_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10393_ cpuregs.regs\[12\]\[28\] cpuregs.regs\[13\]\[28\] cpuregs.regs\[14\]\[28\]
+ cpuregs.regs\[15\]\[28\] _04123_ _04124_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__mux4_1
XANTENNA__11762__A1 alu_out_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09108__B_N _03867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12132_ _06522_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14062__B _07778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09707__A1 _04211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10082__S _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16940_ clknet_leaf_166_clk _00121_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_12063_ _06281_ cpuregs.regs\[22\]\[23\] _06482_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__mux2_1
X_11014_ instr_sub _04913_ _03578_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__o21ba_1
X_16871_ _06586_ cpuregs.regs\[14\]\[25\] _03174_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__mux2_1
XANTENNA__13393__S _07225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18610_ clknet_leaf_106_clk _01675_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10810__S _05363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ _05971_ _02594_ decoded_imm_j\[11\] _03636_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__o2bb2a_1
X_15753_ timer\[25\] timer\[24\] _02547_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__or3_1
X_18541_ clknet_leaf_114_clk _01606_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12965_ _06997_ cpuregs.regs\[31\]\[26\] _06985_ VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__mux2_1
XANTENNA_output216_A net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14704_ _08343_ _07815_ _08344_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__and3b_1
X_11916_ _06407_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_47_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15684_ _02500_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__inv_2
XANTENNA__13019__A1 _06569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18472_ clknet_leaf_149_clk _01537_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_47_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _06124_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__buf_2
XANTENNA__14216__B1 _07901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17423_ clknet_leaf_145_clk _00592_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14635_ _03294_ _07966_ _07997_ _08285_ VGND VGND VPWR VPWR _08286_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11847_ _06369_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_783 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11641__S _06176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17354_ clknet_leaf_148_clk _00523_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_14566_ _08221_ _07952_ _08222_ VGND VGND VPWR VPWR _08223_ sky130_fd_sc_hd__o21ai_1
X_11778_ reg_pc\[29\] _06314_ _06101_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13517_ _07223_ VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__buf_4
X_16305_ _06980_ cpuregs.regs\[15\]\[18\] _02870_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10729_ _05361_ _05411_ _05412_ _05427_ VGND VGND VPWR VPWR alu_out\[5\] sky130_fd_sc_hd__a31o_1
XANTENNA__11450__B1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17285_ clknet_leaf_153_clk _00459_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10257__S _04222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14497_ _07899_ _07939_ _07992_ _08159_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__a31o_1
XFILLER_0_141_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16236_ _02842_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__clkbuf_1
X_13448_ _03524_ decoded_imm\[5\] _07291_ _07289_ _07287_ VGND VGND VPWR VPWR _07309_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__15192__A1 _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_173_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12472__S _06715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16167_ net277 net239 _02797_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__mux2_1
XANTENNA__10781__A _05244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13379_ net89 decoded_imm\[2\] VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__or2_1
XANTENNA__14253__A _07942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11753__A1 alu_out_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12950__A0 _06987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15118_ _01918_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09347__A _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16098_ _03799_ _03833_ _03916_ _03893_ _03891_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__a311o_1
XFILLER_0_121_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16879__S _03174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11088__S _05237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15049_ _03671_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__buf_6
XFILLER_0_76_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_188_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09610_ count_cycle\[6\] _04165_ _04339_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09082__A _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09541_ _04054_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09472_ count_instr\[36\] _04104_ _04145_ count_instr\[4\] VGND VGND VPWR VPWR _04204_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09882__B1 _04604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08423_ mem_rdata_q\[1\] net44 _03208_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12647__S _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_126_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13430__A1 _03631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15707__B1 _02488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10795__A2 _05367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13194__A0 _06949_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13478__S _07225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09937__A1 _04483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13733__A2 _05009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15259__A _02066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12382__S _06663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09257__A _03891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09796__S0 _04325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13507__A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09808_ _04149_ _04528_ _04531_ _04046_ _04532_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__a32o_1
XANTENNA__09548__S0 _04275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09739_ _04463_ _04464_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12750_ _06871_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11701_ _06252_ _03332_ _06253_ _06254_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__a22o_1
XANTENNA__09720__A _04133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15946__B1 _02659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12681_ _06832_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14420_ _08087_ _08088_ VGND VGND VPWR VPWR _08089_ sky130_fd_sc_hd__nand2_1
X_11632_ _06193_ cpuregs.regs\[10\]\[12\] _06176_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10235__B2 _04947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11432__B1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14351_ decoded_imm_j\[4\] _07915_ VGND VGND VPWR VPWR _08025_ sky130_fd_sc_hd__or2_1
X_11563_ _06131_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__buf_2
XFILLER_0_37_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09866__S _04064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13302_ _06989_ cpuregs.regs\[5\]\[22\] _07176_ VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__mux2_1
X_10514_ _05217_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17070_ clknet_leaf_123_clk _00244_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_14282_ reg_pc\[26\] _07953_ _07964_ _07960_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__a22o_1
X_11494_ _06067_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16021_ decoded_imm\[2\] _02711_ _02718_ _02719_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__o22a_1
XANTENNA__15169__A _03647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13233_ _07142_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__clkbuf_1
X_10445_ count_instr\[62\] _04104_ _04017_ count_cycle\[62\] VGND VGND VPWR VPWR _05151_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12292__S _06615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13164_ _06987_ cpuregs.regs\[4\]\[21\] _07104_ VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__mux2_1
X_10376_ _05082_ _05083_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15477__A2 _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12115_ _06513_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__clkbuf_1
X_17972_ clknet_leaf_44_clk _01109_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dfxtp_2
X_13095_ _07069_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14685__B1 _08097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11499__B1 _03338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16923_ clknet_leaf_183_clk _00104_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12046_ _06216_ cpuregs.regs\[22\]\[15\] _06471_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15229__A2 _01906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16854_ _06569_ cpuregs.regs\[14\]\[17\] _03163_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__mux2_1
XANTENNA__12321__A cpuregs.waddr\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15805_ _05960_ _03763_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__and2_1
X_16785_ _03134_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__clkbuf_1
X_13997_ count_instr\[4\] count_instr\[3\] _07761_ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__and3_1
XANTENNA__10149__S1 _04759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15632__A _04271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18524_ clknet_leaf_172_clk _01589_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__14452__A3 _08050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15736_ _04842_ _02506_ _02539_ _02481_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__o211a_1
X_12948_ _06986_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15088__S1 _03646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18455_ clknet_leaf_12_clk _01520_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10776__A _03509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15667_ timer\[2\] _02483_ _02488_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__a21o_1
X_12879_ _06939_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17406_ clknet_leaf_128_clk _00575_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14618_ _08269_ _08270_ VGND VGND VPWR VPWR _08271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13412__A1 _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09616__B1 _04345_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15598_ cpuregs.regs\[4\]\[30\] cpuregs.regs\[5\]\[30\] cpuregs.regs\[6\]\[30\] cpuregs.regs\[7\]\[30\]
+ _01908_ _01909_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__mux4_1
X_18386_ clknet_leaf_128_clk _01451_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10226__A1 _04054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17337_ clknet_leaf_17_clk _00084_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__dfxtp_2
X_14549_ _08203_ _08205_ _08207_ _07905_ reg_next_pc\[19\] VGND VGND VPWR VPWR _01011_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_154_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10777__A2 _05440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16362__A0 _06968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15165__A1 _01989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17268_ clknet_leaf_113_clk _00442_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13176__A0 _06999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13298__S _07176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16219_ net42 mem_16bit_buffer\[2\] _02831_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17199_ clknet_leaf_124_clk _00373_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10529__A2 _04466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16665__A1 _06311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08972_ _03203_ _03733_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_110_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14676__B1 _07904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14979__A1 irq_mask\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13326__S1 _04759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13100__A0 _06991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15640__A2 _07994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09524_ _04244_ _04250_ _04255_ _04008_ irq_pending\[4\] VGND VGND VPWR VPWR _08395_
+ sky130_fd_sc_hd__o32a_2
XFILLER_0_78_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09540__A instr_retirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15079__S1 _01937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10465__B2 _04023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09455_ _04025_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14158__A _06053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08406_ mem_do_rinst mem_do_prefetch VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09386_ irq_pending\[1\] _04008_ _04109_ _04120_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10768__A2 _05261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10312__S1 _04086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15156__A1 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15251__S1 _02014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10230_ _04271_ _04941_ _04942_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__a21o_1
XANTENNA__09386__A2 _04008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10076__S0 _04579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16105__A0 is_alu_reg_reg VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10161_ reg_pc\[21\] decoded_imm\[21\] VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__or2_1
XANTENNA__16312__S _02881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10092_ _04268_ _04788_ _04808_ _03302_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__o211a_1
X_13920_ _07711_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14682__A3 _07971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13851_ cpuregs.regs\[0\]\[22\] VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_145_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12802_ _06898_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15452__A _02066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14434__A3 _08050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13782_ net88 decoded_imm\[29\] VGND VGND VPWR VPWR _07620_ sky130_fd_sc_hd__nand2_1
X_16570_ _06972_ cpuregs.regs\[18\]\[14\] _03015_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__mux2_1
X_10994_ net112 _04880_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__nor2_1
X_12733_ _06859_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__clkbuf_1
X_15521_ cpuregs.regs\[8\]\[25\] cpuregs.regs\[9\]\[25\] cpuregs.regs\[10\]\[25\]
+ cpuregs.regs\[11\]\[25\] _01996_ _01997_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15452_ _02066_ _02290_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__or2_1
X_18240_ clknet_leaf_24_clk _01311_ VGND VGND VPWR VPWR cpuregs.raddr2\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15395__A1 _03709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12664_ _06822_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14403_ decoded_imm_j\[8\] _07924_ VGND VGND VPWR VPWR _08073_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11615_ reg_pc\[11\] _06171_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__nand2_1
X_15383_ cpuregs.regs\[20\]\[17\] cpuregs.regs\[21\]\[17\] cpuregs.regs\[22\]\[17\]
+ cpuregs.regs\[23\]\[17\] _02221_ _02222_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15490__S1 _03642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18171_ clknet_leaf_24_clk _01242_ VGND VGND VPWR VPWR decoded_imm_j\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12595_ cpuregs.regs\[2\]\[31\] _06598_ _06751_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17122_ clknet_leaf_185_clk _00296_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_14334_ decoded_imm_j\[1\] _07902_ _08009_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11546_ _06071_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08821__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15698__A2 _02486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17053_ clknet_leaf_1_clk _00227_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14265_ _07905_ VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11477_ irq_mask\[26\] _03428_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16004_ _03635_ _03763_ _05995_ _06023_ _06025_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_94_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13216_ _07133_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09377__A2 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10428_ _05133_ _05134_ _04320_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_164_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14196_ _07903_ VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13147_ _06970_ cpuregs.regs\[4\]\[13\] _07093_ VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _04215_ _05063_ _05067_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14658__B1 _08232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09129__A2 _03880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09625__A _04341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11874__B _06083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17955_ clknet_leaf_191_clk _01092_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dfxtp_1
X_13078_ _07060_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12029_ _06150_ cpuregs.regs\[22\]\[7\] _06460_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__mux2_1
X_16906_ clknet_leaf_35_clk _00051_ VGND VGND VPWR VPWR mem_rdata_q\[25\] sky130_fd_sc_hd__dfxtp_2
X_17886_ clknet_leaf_90_clk _01055_ VGND VGND VPWR VPWR count_cycle\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11892__A0 _06150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16837_ _06552_ cpuregs.regs\[14\]\[9\] _03152_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16768_ _03125_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09360__A _00073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18507_ clknet_leaf_122_clk _01572_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_15719_ timer\[16\] _02524_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16699_ _03088_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09240_ _03979_ _03902_ _03927_ _03980_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_118_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18438_ clknet_leaf_147_clk _01503_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16583__A0 _06984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09171_ _03908_ _03921_ _03917_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12925__S _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18369_ clknet_leaf_149_clk _01434_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13610__A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08704__A net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15233__S1 _01977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12226__A _06288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09368__A2 _04022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11175__A2 _04710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16638__A1 _06207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12372__A1 _06582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09773__C1 _04149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14649__B1 _07904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15310__A1 _02037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08955_ cpuregs.regs\[24\]\[4\] cpuregs.regs\[25\]\[4\] cpuregs.regs\[26\]\[4\] cpuregs.regs\[27\]\[4\]
+ _03649_ _03643_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__mux4_1
X_08886_ cpuregs.regs\[8\]\[2\] cpuregs.regs\[9\]\[2\] cpuregs.regs\[10\]\[2\] cpuregs.regs\[11\]\[2\]
+ _03649_ _03643_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_162_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12896__A _06124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09828__B1 _04237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10438__A1 _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09270__A _04006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09507_ _04215_ _04230_ _04238_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10438__B2 _05144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09923__S0 _04472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09438_ _04169_ _04170_ _04064_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15472__S1 _02075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09369_ instr_rdinstrh VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__buf_4
XANTENNA__16307__S _02870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13520__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11400_ _03816_ _03916_ _03902_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__a21o_1
X_12380_ cpuregs.regs\[26\]\[27\] _06590_ _06663_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_70 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_81 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10610__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11331_ _05946_ _05948_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__xor2_1
XANTENNA_92 _00001_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15224__S1 _02075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14050_ count_instr\[20\] _07799_ _07790_ VGND VGND VPWR VPWR _07802_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11262_ _05838_ _05890_ _05891_ _05892_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__o31ai_4
XFILLER_0_104_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11166__A2 _05286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13001_ _07019_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__clkbuf_1
X_10213_ _04924_ _04925_ _04575_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__mux2_1
XANTENNA__12570__S _06763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11193_ _05831_ _05835_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15301__A1 decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10144_ cpuregs.regs\[4\]\[21\] cpuregs.regs\[5\]\[21\] cpuregs.regs\[6\]\[21\] cpuregs.regs\[7\]\[21\]
+ _04758_ _04759_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__mux4_1
XANTENNA__13312__A0 _06999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17740_ clknet_leaf_95_clk _00909_ VGND VGND VPWR VPWR count_instr\[11\] sky130_fd_sc_hd__dfxtp_1
X_14952_ _01851_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__clkbuf_1
X_10075_ _04289_ _04791_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ _07699_ VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10677__B2 _05251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17671_ clknet_leaf_172_clk _00840_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_14883_ _01809_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output129_A net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16622_ _03047_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13834_ _07656_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09819__B1 _04017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10429__A1 _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13765_ _07555_ _07567_ VGND VGND VPWR VPWR _07604_ sky130_fd_sc_hd__or2b_1
X_16553_ _06955_ cpuregs.regs\[18\]\[6\] _03004_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10977_ _05544_ _05601_ _05657_ _05660_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15504_ _02037_ _02339_ _02006_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12716_ _06281_ cpuregs.regs\[12\]\[23\] _06847_ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__mux2_1
X_13696_ _07281_ _04941_ _07282_ reg_pc\[23\] VGND VGND VPWR VPWR _07540_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16484_ _02974_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18223_ clknet_leaf_25_clk _01294_ VGND VGND VPWR VPWR instr_retirq sky130_fd_sc_hd__dfxtp_4
XFILLER_0_155_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12647_ _06281_ cpuregs.regs\[30\]\[23\] _06810_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__mux2_1
XANTENNA__15463__S1 _02031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15435_ cpuregs.regs\[20\]\[20\] cpuregs.regs\[21\]\[20\] cpuregs.regs\[22\]\[20\]
+ cpuregs.regs\[23\]\[20\] _01918_ _01919_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18154_ clknet_leaf_73_clk alu_out\[28\] VGND VGND VPWR VPWR alu_out_q\[28\] sky130_fd_sc_hd__dfxtp_1
X_15366_ _02012_ _02209_ _01968_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12578_ _06777_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08524__A _03277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10601__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10062__C1 _03302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15215__S1 _01986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17105_ clknet_leaf_162_clk _00279_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_11529_ _06074_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__buf_2
X_14317_ _07993_ VGND VGND VPWR VPWR _07994_ sky130_fd_sc_hd__inv_2
X_18085_ clknet_leaf_102_clk _01189_ VGND VGND VPWR VPWR timer\[0\] sky130_fd_sc_hd__dfxtp_1
X_15297_ cpuregs.regs\[16\]\[12\] cpuregs.regs\[17\]\[12\] cpuregs.regs\[18\]\[12\]
+ cpuregs.regs\[19\]\[12\] _02074_ _02075_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14248_ reg_next_pc\[16\] _05858_ _07922_ _07940_ VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__o211a_2
X_17036_ clknet_leaf_180_clk _00210_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15357__A _01989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14179_ count_instr\[59\] _07887_ count_instr\[60\] VGND VGND VPWR VPWR _07891_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12480__S _06715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16096__A2 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08740_ net100 net68 VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__nand2_1
X_17938_ clknet_leaf_69_clk _08378_ VGND VGND VPWR VPWR reg_out\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10117__B1 _04296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09522__A2 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10212__S0 _04512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11865__A0 _06320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08671_ _03435_ _03436_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__or2_1
X_17869_ clknet_leaf_94_clk _01038_ VGND VGND VPWR VPWR count_cycle\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13606__A1 _03276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09905__S0 _04290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11125__A _05517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09223_ _03754_ _03771_ _03772_ _03753_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__a22o_2
XANTENNA__12655__S _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16127__S _02771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09154_ _03906_ _03895_ _03908_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11396__A2 _03636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09249__B _03885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09085_ _03757_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15531__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12345__A1 _06554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16087__A2 _02650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10451__S0 _04085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09987_ _04703_ _04704_ _04706_ _04010_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__o22a_1
XANTENNA__16797__S _03138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15295__B1 _03654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08938_ _03683_ _03697_ _03701_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__a21o_1
XANTENNA__10659__A1 _05255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08869_ _03634_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10900_ _04642_ net72 net71 net70 _05236_ _05309_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__mux4_1
X_11880_ _06096_ cpuregs.regs\[20\]\[1\] _06387_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__mux2_1
XANTENNA__16795__A0 _06578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10831_ _05278_ _05523_ _05228_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__o21a_1
XFILLER_0_168_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13550_ _07404_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16547__A0 _06949_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10762_ _05372_ _05379_ _05374_ _05370_ _05395_ _05287_ VGND VGND VPWR VPWR _05459_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12501_ _06248_ cpuregs.regs\[28\]\[19\] _06726_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13481_ _04360_ _05260_ _07301_ _07279_ VGND VGND VPWR VPWR _07340_ sky130_fd_sc_hd__o211a_1
XANTENNA__09029__A1 mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10693_ _03529_ _05391_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15220_ _02012_ _02071_ _02017_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__o21a_1
XANTENNA__12033__A0 _06166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12432_ cpuregs.regs\[27\]\[19\] _06573_ _06689_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15151_ _02005_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_152_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10085__S _04320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12363_ cpuregs.regs\[26\]\[19\] _06573_ _06652_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16561__A _03003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08883__S0 _03645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14102_ _07836_ _07837_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__nor2_1
X_11314_ _03841_ _05933_ _05934_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_91_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15082_ _03709_ _01938_ _01940_ _00067_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__o211a_1
X_12294_ cpuregs.regs\[25\]\[19\] _06573_ _06615_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11139__A2 _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14033_ _06053_ VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11909__S _06398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11245_ _05872_ _05877_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__or2_1
XANTENNA__15177__A _03684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09175__A _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11176_ _04038_ net127 net104 _03297_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output246_A net246 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15286__B1 _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10127_ irq_mask\[20\] _04448_ timer\[20\] _04024_ _04027_ VGND VGND VPWR VPWR _04843_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__15381__S0 _03641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16500__S _02979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15984_ _03856_ _02698_ _02699_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__a21bo_1
X_17723_ clknet_leaf_76_clk _00892_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dfxtp_1
XANTENNA__09903__A _04070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10058_ _04763_ _04767_ _04133_ _04775_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__o211ai_4
X_14935_ _01842_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13425__A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17654_ clknet_leaf_47_clk _00823_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfxtp_2
XANTENNA__09622__B decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16786__A0 _06569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14866_ count_cycle\[57\] _01795_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16605_ _07007_ cpuregs.regs\[18\]\[31\] _03003_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__mux2_1
X_13817_ cpuregs.regs\[0\]\[5\] VGND VGND VPWR VPWR _07648_ sky130_fd_sc_hd__clkbuf_1
X_17585_ clknet_leaf_131_clk _00754_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_14797_ count_cycle\[34\] _01748_ _01751_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16536_ _03001_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__clkbuf_1
X_13748_ _07586_ _07588_ _07190_ VGND VGND VPWR VPWR _07589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16002__A2 _06016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15436__S1 _01919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16467_ _07005_ cpuregs.regs\[29\]\[30\] _02931_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13679_ net81 decoded_imm\[22\] VGND VGND VPWR VPWR _07524_ sky130_fd_sc_hd__nand2_1
XANTENNA__14256__A _07904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18206_ clknet_leaf_42_clk _01277_ VGND VGND VPWR VPWR instr_add sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15418_ _02005_ _02254_ _02256_ _02258_ _03692_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__a221o_2
XFILLER_0_26_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_959 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16398_ _02928_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11378__A2 _03636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12575__A1 _06578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18137_ clknet_leaf_47_clk alu_out\[11\] VGND VGND VPWR VPWR alu_out_q\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10586__A0 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15349_ _02192_ _02193_ _02002_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18068_ clknet_leaf_73_clk _01173_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_151_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09991__A2 _04710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11819__S _06348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09910_ _04051_ _04631_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__nor2_1
X_17019_ clknet_leaf_2_clk _00193_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08701__B net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16069__A2 _02650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09841_ _04268_ _04544_ _04564_ _04149_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__o211a_1
XANTENNA__09085__A _03757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10984__S1 _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15816__A2 _06016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09772_ count_cycle\[10\] _04013_ _04497_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__a21o_1
XANTENNA__15815__A decoded_imm_j\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _03479_ _03482_ _03485_ _03488_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__or4_1
XANTENNA__11838__A0 _06216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15029__B1 _01714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08654_ _03418_ _03419_ _03420_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_87_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _03195_ _03363_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_120_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09354__S1 _04087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10813__A1 _05288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_946 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12015__A0 _06078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09206_ _03730_ _03848_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12566__A1 _06569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11302__B _05923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09137_ _03891_ _03893_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__nor2_2
XFILLER_0_115_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10672__S0 _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15504__A1 _02037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09068_ net63 _03730_ _03829_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11030_ _03581_ _05709_ _05390_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__mux2_1
XANTENNA__09734__A2 _04008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10424__S0 _04057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15268__B1 _02027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15363__S0 _01990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16320__S _02881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12981_ _07008_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14720_ count_cycle\[10\] _08353_ _08355_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11932_ _06304_ cpuregs.regs\[20\]\[26\] _06409_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11863_ _06312_ cpuregs.regs\[11\]\[27\] _06370_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__mux2_1
X_14651_ _07966_ _07967_ _08277_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__and3_1
XFILLER_0_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10814_ _03507_ _05220_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13602_ _04642_ _05258_ VGND VGND VPWR VPWR _07453_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17370_ clknet_leaf_119_clk _00539_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_11794_ _06337_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__clkbuf_1
X_14582_ _08236_ _08121_ _08237_ VGND VGND VPWR VPWR _08238_ sky130_fd_sc_hd__and3b_1
XFILLER_0_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16321_ _02887_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13533_ _04532_ _07315_ _07358_ _07254_ VGND VGND VPWR VPWR _07388_ sky130_fd_sc_hd__o211a_1
X_10745_ _05442_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10280__A2 _04016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13464_ _07324_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__clkbuf_1
X_16252_ _02850_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__clkbuf_1
X_10676_ _05243_ _05376_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_49 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14546__A2 _07950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output196_A net196 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15203_ _02054_ _02055_ _03666_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__mux2_1
X_12415_ _06690_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10568__A0 _05044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13395_ net92 decoded_imm\[3\] VGND VGND VPWR VPWR _07259_ sky130_fd_sc_hd__nand2_1
X_16183_ net286 net248 _02770_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12346_ _06653_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__clkbuf_1
X_15134_ _03666_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__buf_4
Xoutput209 net209 VGND VGND VPWR VPWR mem_la_addr[25] sky130_fd_sc_hd__buf_1
XFILLER_0_51_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12309__A1 _06588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15065_ cpuregs.regs\[16\]\[0\] cpuregs.regs\[17\]\[0\] cpuregs.regs\[18\]\[0\] cpuregs.regs\[19\]\[0\]
+ _03670_ _03671_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__mux4_1
XANTENNA__09617__B decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12277_ _06616_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14016_ _03304_ VGND VGND VPWR VPWR _07778_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_output73_A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11228_ _05862_ _05864_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__nand2_1
XANTENNA__10415__S0 _04579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11159_ _05814_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15967_ _02686_ _02687_ _02684_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_69_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14482__B2 _06863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17706_ clknet_leaf_75_clk _00875_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14918_ _01833_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12493__A0 _06216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09584__S1 _04219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15898_ _02642_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_172_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17637_ clknet_leaf_50_clk _00806_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfxtp_4
X_14849_ count_cycle\[51\] _01783_ _01723_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_102_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17568_ clknet_leaf_170_clk _00737_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15982__A1 _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16519_ cpuregs.regs\[17\]\[22\] _06580_ _02990_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17499_ clknet_leaf_20_clk _00668_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10271__A2 _04959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10019__A _04737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16405__S _02932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_1019 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10961__B _05334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10453__S _04078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09527__B decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15593__S0 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09824_ _04231_ _04547_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__nand2_1
XANTENNA__15345__S0 _02069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09543__A _04273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09755_ _04479_ _04480_ _04078_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__mux2_1
X_08706_ _03470_ _03471_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09686_ _04099_ _04405_ _04413_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__or3_4
XPHY_EDGE_ROW_169_Left_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08637_ _03406_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_159_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08568_ irq_mask\[25\] irq_pending\[25\] VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__and2b_1
XANTENNA__09327__S1 _04060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15973__A1 mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15973__B2 _04022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08499_ _03218_ _03278_ cpu_state\[6\] VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__or3b_2
XANTENNA__09652__A1 _04206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10798__B1 _05322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10530_ _04566_ _04602_ _04611_ _04642_ _05230_ _05232_ VGND VGND VPWR VPWR _05234_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_172_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15725__A1 _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10461_ _04053_ _05166_ _04095_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__a21o_1
XANTENNA__12843__S _06917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12200_ _06566_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09955__A2 _04049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13180_ _07003_ cpuregs.regs\[4\]\[29\] _07104_ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__mux2_1
X_10392_ _05098_ _05099_ _04222_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12131_ _06281_ cpuregs.regs\[23\]\[23\] _06518_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__mux2_1
XANTENNA__16150__A1 net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15584__S0 _01908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12062_ _06485_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11013_ _05590_ _05601_ _05690_ _05281_ _05693_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__a221o_1
X_16870_ _03179_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ _05960_ _03737_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__nand2_1
XANTENNA__15110__C1 _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09453__A _04185_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11278__A1 _03475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18540_ clknet_leaf_164_clk _01605_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_15752_ timer\[24\] _02547_ timer\[25\] VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__o21a_1
X_12964_ _06303_ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__buf_2
XANTENNA__13672__C1 _07217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16205__A2 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14703_ count_cycle\[4\] _08340_ count_cycle\[5\] VGND VGND VPWR VPWR _08344_ sky130_fd_sc_hd__a21o_1
X_11915_ _06240_ cpuregs.regs\[20\]\[18\] _06398_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__mux2_1
X_18471_ clknet_leaf_156_clk _01536_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_output111_A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15683_ timer\[0\] _03416_ _03427_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_47_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _06950_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output209_A net209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11922__S _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17422_ clknet_leaf_137_clk _00591_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ _07998_ _08277_ VGND VGND VPWR VPWR _08285_ sky130_fd_sc_hd__or2_1
X_11846_ _06248_ cpuregs.regs\[11\]\[19\] _06359_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__mux2_1
XANTENNA__12778__A1 _06565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17353_ clknet_leaf_159_clk _00522_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11777_ reg_pc\[29\] reg_pc\[28\] _06306_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09643__A1 _04289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14565_ decoded_imm_j\[19\] _07950_ _07952_ _08212_ VGND VGND VPWR VPWR _08222_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16304_ _02878_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10728_ _05298_ _05415_ _05421_ _05426_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__a211o_1
X_13516_ _07367_ _07370_ _07372_ _07284_ VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_60_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17284_ clknet_leaf_160_clk _00458_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14496_ reg_next_pc\[15\] _07947_ _08158_ _08033_ VGND VGND VPWR VPWR _08159_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16235_ net51 mem_16bit_buffer\[10\] _02830_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10659_ _05255_ _05261_ _05337_ _05360_ VGND VGND VPWR VPWR alu_out\[2\] sky130_fd_sc_hd__a31o_1
X_13447_ _07308_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12753__S _06869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14534__A _03293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13378_ net89 decoded_imm\[2\] VGND VGND VPWR VPWR _07243_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16166_ _02801_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10781__B _05334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15117_ cpuregs.regs\[4\]\[5\] cpuregs.regs\[5\]\[5\] cpuregs.regs\[6\]\[5\] cpuregs.regs\[7\]\[5\]
+ _01970_ _01971_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__mux4_1
X_12329_ _06644_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15575__S0 _02030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16097_ _03747_ _03781_ _03768_ _02759_ _06009_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__o221a_1
XANTENNA__14152__B1 _07834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15048_ _03670_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__buf_6
XANTENNA__15327__S0 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16999_ clknet_leaf_147_clk _00173_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_09540_ instr_retirq VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__buf_4
XANTENNA__12466__A0 _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09082__B _03781_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10302__A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09471_ _04191_ _04197_ _04203_ _04008_ irq_pending\[3\] VGND VGND VPWR VPWR _08394_
+ sky130_fd_sc_hd__o32a_2
XFILLER_0_78_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12928__S _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09882__B2 _03225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11832__S _06359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08422_ _03207_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10229__C1 _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09634__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08437__A2 _03215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12229__A _06296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09634__B2 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16135__S _02771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08442__A _03225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10183__S _04065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09972__S _04121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12899__A _06131_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15891__B1 _02623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09796__S1 _04277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09273__A _04009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09807_ net69 VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__buf_4
XANTENNA__13507__B decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14446__A1 _07899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09738_ _04453_ _04454_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09548__S1 _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09873__A1 _04010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09669_ _04105_ count_cycle\[40\] _04013_ count_cycle\[8\] _04396_ VGND VGND VPWR
+ VPWR _04397_ sky130_fd_sc_hd__a221o_1
XFILLER_0_173_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11700_ reg_out\[20\] alu_out_q\[20\] _06068_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15946__A1 _04012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12680_ _06141_ cpuregs.regs\[12\]\[6\] _06825_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10866__B _05227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15946__B2 _02669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09212__S _03757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11631_ _06192_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10235__A2 _04006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14350_ decoded_imm_j\[4\] _07915_ VGND VGND VPWR VPWR _08024_ sky130_fd_sc_hd__nand2_1
X_11562_ _06075_ _06127_ _06130_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_147_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10513_ _05211_ _05216_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__or2_1
X_13301_ _07178_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14281_ reg_next_pc\[26\] _05928_ _07942_ _07963_ VGND VGND VPWR VPWR _07964_ sky130_fd_sc_hd__o211a_2
X_11493_ latched_stalu VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12573__S _06774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16020_ _02715_ decoded_imm_j\[2\] _02716_ mem_rdata_q\[9\] _02633_ VGND VGND VPWR
+ VPWR _02719_ sky130_fd_sc_hd__a221o_1
X_13232_ _06987_ cpuregs.regs\[8\]\[21\] _07140_ VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__mux2_1
X_10444_ _05148_ _05149_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_1002 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13163_ _07105_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__clkbuf_1
X_10375_ reg_pc\[28\] decoded_imm\[28\] VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16123__A1 _05286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12114_ _06216_ cpuregs.regs\[23\]\[15\] _06507_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__mux2_1
X_17971_ clknet_leaf_4_clk _01108_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dfxtp_1
X_13094_ _06984_ cpuregs.regs\[7\]\[20\] _07068_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__mux2_1
XANTENNA__10106__B decoded_imm\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14801__B _01753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11917__S _06398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16922_ clknet_leaf_183_clk _00103_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12045_ _06476_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11499__B2 _06072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16853_ _03170_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__clkbuf_1
X_15804_ decoded_imm_j\[3\] _05983_ _03895_ _06016_ _05985_ VGND VGND VPWR VPWR _01233_
+ sky130_fd_sc_hd__a221o_1
X_16784_ _06567_ cpuregs.regs\[13\]\[16\] _03127_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13996_ _07763_ _07764_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__nor2_1
X_18523_ clknet_leaf_178_clk _01588_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_15735_ _02476_ _02537_ _02538_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__or3b_1
XFILLER_0_133_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15632__B instr_jalr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12947_ _06984_ cpuregs.regs\[31\]\[20\] _06985_ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18454_ clknet_leaf_189_clk _01519_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15666_ _02475_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12878_ _06336_ cpuregs.regs\[6\]\[30\] _06905_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__mux2_1
XANTENNA__10776__B _05301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17405_ clknet_leaf_119_clk _00574_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_14617_ _08221_ _08268_ VGND VGND VPWR VPWR _08270_ sky130_fd_sc_hd__or2_1
XANTENNA__09616__A1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14963__S _07755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11829_ _06360_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__clkbuf_1
X_18385_ clknet_leaf_113_clk _01450_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15597_ net120 _01906_ _02427_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__o21a_1
XANTENNA__13412__A2 _05260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09616__B2 _03225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17336_ clknet_leaf_176_clk _00510_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14548_ _07988_ _08206_ VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12483__S _06726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17267_ clknet_leaf_165_clk _00441_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14479_ _08128_ _08131_ _08141_ VGND VGND VPWR VPWR _08143_ sky130_fd_sc_hd__or3b_1
XFILLER_0_153_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16218_ _02833_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09919__A2 decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17198_ clknet_leaf_123_clk _00372_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10529__A3 _04532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16114__A1 _03199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16149_ _02792_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08971_ net53 mem_rdata_q\[28\] _03730_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14676__A1 _07898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14676__B2 reg_next_pc\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11034__S0 _05264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09093__A _03767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09523_ _03680_ _04251_ _04254_ _03226_ _04202_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__a221o_2
XFILLER_0_79_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13343__A instr_lui VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09454_ instr_timer VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10465__A2 _04308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08405_ reg_out\[1\] _03188_ _03190_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__o21ai_2
X_09385_ _03226_ _04112_ _04119_ _04049_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__a211o_1
XANTENNA__13403__A2 _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09607__B2 _04187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10768__A3 _05458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12393__S _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_140_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_140_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__15156__A2 _01906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11178__B1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10076__S1 _04284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14116__B1 _07675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10160_ reg_pc\[21\] decoded_imm\[21\] VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_7_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09791__B1 _04296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15864__B1 _02620_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12678__A0 _06132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10091_ _04271_ _04806_ _04807_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15616__B1 _00068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13850_ _07664_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_145_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12801_ cpuregs.regs\[9\]\[26\] _06588_ _06891_ VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__mux2_1
X_13781_ _07619_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__clkbuf_1
X_10993_ _03574_ _05663_ _03577_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12568__S _06763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_172_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09846__B2 _04569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15520_ _02351_ _02352_ _02353_ _02354_ _02111_ _03639_ VGND VGND VPWR VPWR _02355_
+ sky130_fd_sc_hd__mux4_1
X_12732_ _06343_ cpuregs.regs\[12\]\[31\] _06824_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15451_ cpuregs.regs\[16\]\[21\] cpuregs.regs\[17\]\[21\] cpuregs.regs\[18\]\[21\]
+ cpuregs.regs\[19\]\[21\] _01996_ _01997_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12663_ _06343_ cpuregs.regs\[30\]\[31\] _06787_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14402_ decoded_imm_j\[8\] _07924_ VGND VGND VPWR VPWR _08072_ sky130_fd_sc_hd__and2_1
X_11614_ _06177_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11405__A1 _03867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18170_ clknet_leaf_24_clk _01241_ VGND VGND VPWR VPWR decoded_imm_j\[11\] sky130_fd_sc_hd__dfxtp_1
X_15382_ _02223_ _02224_ _02110_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_187_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12594_ _06785_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17121_ clknet_leaf_184_clk _00295_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[8\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14333_ _08007_ _08008_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__nor2_1
X_11545_ _06115_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_131_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_131_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17052_ clknet_leaf_3_clk _00226_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11476_ _06054_ irq_pending\[25\] _06057_ net18 VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__a31o_1
X_14264_ reg_pc\[20\] _07926_ _07952_ _07935_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16003_ cpuregs.raddr1\[3\] _06006_ _06020_ _06022_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_94_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13215_ _06970_ cpuregs.regs\[8\]\[13\] _07129_ VGND VGND VPWR VPWR _07133_ sky130_fd_sc_hd__mux2_1
X_10427_ cpuregs.regs\[0\]\[29\] cpuregs.regs\[1\]\[29\] cpuregs.regs\[2\]\[29\] cpuregs.regs\[3\]\[29\]
+ _04487_ _04469_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14195_ _03298_ _03196_ VGND VGND VPWR VPWR _07903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09782__B1 _03225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13146_ _07096_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__clkbuf_1
X_10358_ _04231_ _05066_ _04237_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__a21o_1
XANTENNA__08810__A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_115_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14658__A1 _07966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17954_ clknet_leaf_191_clk _01091_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__dfxtp_1
X_13077_ _06968_ cpuregs.regs\[7\]\[12\] _07057_ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_125_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _04206_ _04999_ _04225_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12028_ _06467_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__clkbuf_1
X_16905_ clknet_leaf_34_clk _00050_ VGND VGND VPWR VPWR mem_rdata_q\[24\] sky130_fd_sc_hd__dfxtp_2
X_17885_ clknet_leaf_89_clk _01054_ VGND VGND VPWR VPWR count_cycle\[30\] sky130_fd_sc_hd__dfxtp_1
X_16836_ _03161_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13618__C1 _07283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13094__A0 _06984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16767_ _06550_ cpuregs.regs\[13\]\[8\] _03116_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__mux2_1
XANTENNA__12478__S _06715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13979_ _03331_ _07677_ _07681_ net155 VGND VGND VPWR VPWR _07752_ sky130_fd_sc_hd__a22o_1
X_18506_ clknet_leaf_121_clk _01571_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_15718_ timer\[16\] _02524_ _02488_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__a21o_1
XANTENNA__12841__A0 _06193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16698_ _06963_ cpuregs.regs\[19\]\[10\] _03087_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_124_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18437_ clknet_leaf_135_clk _01502_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15649_ mem_do_wdata _03278_ _04006_ _07904_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__or4b_1
XFILLER_0_118_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09170_ mem_rdata_q\[19\] _03920_ _03914_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__mux2_1
X_18368_ clknet_leaf_160_clk _01433_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17319_ clknet_leaf_145_clk _00493_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13610__B decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09470__C1 _04202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_122_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_122_clk sky130_fd_sc_hd__clkbuf_2
X_18299_ clknet_leaf_5_clk _01367_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08704__B net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13102__S _07068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09448__S0 _04055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16413__S _02932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14361__A3 _07992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08720__A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14649__A1 _03293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14649__B2 reg_next_pc\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08954_ cpuregs.regs\[28\]\[4\] cpuregs.regs\[29\]\[4\] cpuregs.regs\[30\]\[4\] cpuregs.regs\[31\]\[4\]
+ _03649_ _03643_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11332__A0 _05143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_189_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_189_clk sky130_fd_sc_hd__clkbuf_2
X_08885_ cpuregs.regs\[12\]\[2\] cpuregs.regs\[13\]\[2\] cpuregs.regs\[14\]\[2\] cpuregs.regs\[15\]\[2\]
+ _03649_ _03643_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10135__B2 irq_pending\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09551__A _04281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09828__A1 _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12388__S _06640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11292__S _03219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09506_ _04231_ _04236_ _04237_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10438__A2 _05143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09923__S1 _04473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09437_ cpuregs.regs\[24\]\[3\] cpuregs.regs\[25\]\[3\] cpuregs.regs\[26\]\[3\] cpuregs.regs\[27\]\[3\]
+ _04056_ _04086_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09368_ irq_mask\[1\] _04022_ timer\[1\] _04024_ _04027_ VGND VGND VPWR VPWR _04103_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13520__B decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09299_ _04033_ mem_wordsize\[2\] _04034_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__o21a_2
XFILLER_0_7_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_113_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_113_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA_60 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08614__B _03254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10071__B1 _04013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ reg_out\[29\] _05941_ _05947_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_10_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_82 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14337__B1 _08012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 _01908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15728__A _02476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11261_ _04708_ _05838_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12851__S _06917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13000_ cpuregs.regs\[3\]\[8\] _06550_ _07010_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__mux2_1
X_10212_ cpuregs.regs\[8\]\[23\] cpuregs.regs\[9\]\[23\] cpuregs.regs\[10\]\[23\]
+ cpuregs.regs\[11\]\[23\] _04512_ _04513_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__mux4_1
X_11192_ reg_next_pc\[4\] reg_out\[4\] _05834_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_37_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08630__A instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10143_ _04272_ _04857_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__nand2_1
XANTENNA__15301__A2 _02009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12152__A _06533_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14951_ net210 net179 _01846_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__mux2_1
X_10074_ _04789_ _04790_ _04321_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__mux2_1
X_13902_ _07691_ _07698_ VGND VGND VPWR VPWR _07699_ sky130_fd_sc_hd__and2_1
X_17670_ clknet_leaf_177_clk _00839_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14882_ _01807_ _01753_ _01808_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_50_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16621_ cpuregs.regs\[1\]\[6\] _06140_ _03040_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__mux2_1
X_13833_ cpuregs.regs\[0\]\[13\] VGND VGND VPWR VPWR _07656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16552_ _03010_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__clkbuf_1
X_13764_ _07602_ VGND VGND VPWR VPWR _07603_ sky130_fd_sc_hd__inv_2
X_10976_ _05404_ _05622_ _05659_ _05251_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__a2bb2o_1
X_15503_ _02337_ _02338_ _01984_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12715_ _06850_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__clkbuf_1
X_16483_ cpuregs.regs\[17\]\[5\] _06544_ _02968_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__mux2_1
X_13695_ _07274_ _07538_ _07191_ VGND VGND VPWR VPWR _07539_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11930__S _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18222_ clknet_leaf_38_clk _01293_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dfxtp_4
XANTENNA__15402__S _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15434_ _02270_ _02271_ _02272_ _02273_ _02111_ _02088_ VGND VGND VPWR VPWR _02274_
+ sky130_fd_sc_hd__mux4_1
X_12646_ _06813_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09678__S0 _04085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18153_ clknet_leaf_45_clk alu_out\[27\] VGND VGND VPWR VPWR alu_out_q\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15365_ cpuregs.regs\[12\]\[16\] cpuregs.regs\[13\]\[16\] cpuregs.regs\[14\]\[16\]
+ cpuregs.regs\[15\]\[16\] _02013_ _02014_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_104_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_104_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_136_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12577_ cpuregs.regs\[2\]\[22\] _06580_ _06774_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_943 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17104_ clknet_leaf_164_clk _00278_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14316_ _03369_ _07983_ VGND VGND VPWR VPWR _07993_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18084_ clknet_leaf_27_clk _00000_ VGND VGND VPWR VPWR decoder_trigger sky130_fd_sc_hd__dfxtp_4
X_11528_ _06098_ _06099_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__and2_1
X_15296_ cpuregs.regs\[20\]\[12\] cpuregs.regs\[21\]\[12\] cpuregs.regs\[22\]\[12\]
+ cpuregs.regs\[23\]\[12\] _01999_ _02000_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17035_ clknet_leaf_177_clk _00209_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_14247_ _05856_ _06221_ VGND VGND VPWR VPWR _07940_ sky130_fd_sc_hd__or2_1
XANTENNA__12761__S _06869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11459_ irq_mask\[18\] _06042_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_74_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14178_ count_instr\[60\] count_instr\[59\] _07887_ VGND VGND VPWR VPWR _07890_ sky130_fd_sc_hd__and3_1
XANTENNA__09850__S0 _04512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15828__B1 _03781_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13129_ _07087_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__clkbuf_1
X_17937_ clknet_leaf_66_clk _08377_ VGND VGND VPWR VPWR reg_out\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10117__A1 _04215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13592__S _07374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08670_ net122 net90 VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__and2_1
XANTENNA__10668__A2 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17868_ clknet_leaf_94_clk _01037_ VGND VGND VPWR VPWR count_cycle\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10212__S1 _04513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16819_ _06531_ cpuregs.regs\[14\]\[0\] _03152_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_132_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17799_ clknet_leaf_57_clk _00968_ VGND VGND VPWR VPWR reg_pc\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_88_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11617__A1 alu_out_q\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12001__S _06446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09905__S1 _04276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12290__A1 _06569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11840__S _06359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09222_ _03838_ _03955_ _03964_ _03888_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08715__A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09153_ _03907_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_90_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10053__B1 _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09994__B1 _04707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09084_ _03739_ _03844_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__and2_2
XFILLER_0_4_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_141_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_662 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15531__A2 _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13542__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09546__A _04276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14171__B _07815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10191__S _04064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09986_ count_instr\[48\] _04016_ count_cycle\[16\] _04014_ _04705_ VGND VGND VPWR
+ VPWR _04706_ sky130_fd_sc_hd__a221o_1
XANTENNA__10451__S1 _04087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15295__A1 _02066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08937_ _03657_ _03700_ _03675_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__a21o_1
XANTENNA__10204__B decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10659__A2 _05261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08868_ _03633_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_150_Left_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09281__A _04017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13058__A0 _06949_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12528__D_N _06083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_637 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08799_ net106 net74 VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__or2b_1
XANTENNA__13007__S _07021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10830_ _05370_ _05372_ _05331_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10761_ _05455_ _05457_ _05278_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__mux2_1
XANTENNA__16318__S _02881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14627__A _08050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12500_ _06735_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10692_ _03529_ _05391_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__nand2_1
X_13480_ _04566_ _07276_ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__or2_1
X_12431_ _06698_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13230__A0 _06984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09985__B1 _04105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15150_ _03656_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__clkbuf_8
X_12362_ _06661_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13677__S _07374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14101_ count_instr\[36\] _07833_ _07834_ VGND VGND VPWR VPWR _07837_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08883__S1 _03647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11313_ _05925_ _05929_ _05932_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__and3_1
XANTENNA__10890__A _05414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15081_ _03713_ _01939_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__or2_1
X_12293_ _06624_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12581__S _06774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14362__A _03379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13533__A1 _04532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14032_ count_instr\[15\] _07787_ VGND VGND VPWR VPWR _07789_ sky130_fd_sc_hd__and2_1
X_11244_ _05872_ _05877_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11544__A0 _06114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14081__B _07815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09832__S0 _04084_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11175_ net120 _04710_ _05822_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_52_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09175__B _03892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15286__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10126_ _04829_ _04833_ _04841_ _04227_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__a211oi_4
X_15983_ _03844_ _05963_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__nor2_1
XANTENNA__15381__S1 _03684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output239_A net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17722_ clknet_leaf_77_clk _00891_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dfxtp_1
XANTENNA__15193__A _03669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13706__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10057_ _04769_ _04771_ _04774_ _04231_ _04237_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__a221o_1
X_14934_ net202 net171 _01835_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__mux2_1
XANTENNA__16235__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08803__B_N net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17653_ clknet_leaf_48_clk _00822_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dfxtp_2
X_14865_ _01797_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13425__B decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16604_ _03037_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__clkbuf_1
X_13816_ _07647_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__clkbuf_1
X_17584_ clknet_leaf_129_clk _00753_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14796_ count_cycle\[34\] _01748_ _01717_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_67_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16535_ cpuregs.regs\[17\]\[30\] _06596_ _02967_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13747_ _07209_ _07587_ _07210_ reg_pc\[26\] VGND VGND VPWR VPWR _07588_ sky130_fd_sc_hd__a22o_1
X_10959_ _04810_ _04754_ _04744_ _04708_ _05237_ _05240_ VGND VGND VPWR VPWR _05644_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_128_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14537__A decoded_imm_j\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14549__B1 _07905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16466_ _02964_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__clkbuf_1
X_13678_ _07523_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18205_ clknet_leaf_41_clk _01276_ VGND VGND VPWR VPWR instr_srli sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15417_ _03666_ _02257_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__or2_1
XANTENNA__15974__D_N _03977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12629_ _06804_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__clkbuf_1
X_16397_ _07003_ cpuregs.regs\[16\]\[29\] _02918_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18136_ clknet_leaf_48_clk alu_out\[10\] VGND VGND VPWR VPWR alu_out_q\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15348_ cpuregs.regs\[24\]\[15\] cpuregs.regs\[25\]\[15\] cpuregs.regs\[26\]\[15\]
+ cpuregs.regs\[27\]\[15\] _02074_ _02075_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10586__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_693 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18067_ clknet_leaf_72_clk _01172_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_170_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12491__S _06726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15279_ _02012_ _02127_ _02005_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17018_ clknet_leaf_190_clk _00192_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10338__A1 _04391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09840_ _04271_ _04562_ _04563_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09771_ _04017_ count_cycle\[42\] _03252_ _04496_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__a211o_1
X_08722_ _03486_ _03487_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_107_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09305__S _04040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08653_ timer\[17\] timer\[16\] timer\[19\] timer\[18\] VGND VGND VPWR VPWR _03420_
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_87_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10040__A _04232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08584_ _03340_ _03361_ _03362_ decoder_trigger VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__o211a_2
XFILLER_0_49_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16529__A1 _06590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14447__A decoded_imm_j\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08445__A _03199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09040__S _03730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09205_ _03848_ _03946_ _03950_ _03888_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09136_ _03862_ _03879_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__nand2_1
XANTENNA__09431__A2 _04159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10121__S0 _04282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09067_ mem_rdata_q\[8\] _03208_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10672__S1 _05324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15060__S0 _01918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09276__A _03253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10329__B2 _04187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16601__S _03026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10424__S1 _04060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08942__A1 _03638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09969_ _04054_ _04688_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__nand2_1
XANTENNA__15363__S1 _01992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11745__S _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13526__A _04642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12980_ _07007_ cpuregs.regs\[31\]\[31\] _06942_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__mux2_1
XANTENNA__16217__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11931_ _06415_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10501__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14650_ _07966_ _08277_ _07967_ VGND VGND VPWR VPWR _08300_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11862_ _06377_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__clkbuf_1
X_13601_ _04566_ _05259_ _07451_ _07217_ VGND VGND VPWR VPWR _07452_ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10813_ _05288_ _05332_ _05506_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _07952_ _07954_ _08206_ _07956_ VGND VGND VPWR VPWR _08237_ sky130_fd_sc_hd__a31o_1
XANTENNA__09655__C1 _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11793_ _06336_ cpuregs.regs\[10\]\[30\] _06085_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10265__B1 _04080_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16320_ _06995_ cpuregs.regs\[15\]\[25\] _02881_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__mux2_1
X_13532_ _07387_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10744_ _05441_ _05401_ _05231_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16251_ mem_rdata_q\[2\] _03864_ _03914_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13463_ _04342_ _07323_ _07225_ VGND VGND VPWR VPWR _07324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09407__C1 _00073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10675_ _04198_ _04160_ _04039_ _04036_ _05236_ _05239_ VGND VGND VPWR VPWR _05376_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15202_ cpuregs.regs\[28\]\[7\] cpuregs.regs\[29\]\[7\] cpuregs.regs\[30\]\[7\] cpuregs.regs\[31\]\[7\]
+ _03640_ _03642_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__mux4_1
XANTENNA__13754__A1 _04945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14951__A0 net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12414_ cpuregs.regs\[27\]\[10\] _06554_ _06689_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__mux2_1
X_16182_ _02809_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10568__A1 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13394_ _07258_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15133_ _01984_ _01987_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__or2_1
X_12345_ cpuregs.regs\[26\]\[10\] _06554_ _06652_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_1006 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13200__S _07118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15051__S0 _03658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09186__A _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15064_ cpuregs.regs\[20\]\[0\] cpuregs.regs\[21\]\[0\] cpuregs.regs\[22\]\[0\] cpuregs.regs\[23\]\[0\]
+ _03670_ _03671_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__mux4_1
X_12276_ cpuregs.regs\[25\]\[10\] _06554_ _06615_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__mux2_1
X_14015_ count_instr\[10\] count_instr\[9\] _07773_ VGND VGND VPWR VPWR _07777_ sky130_fd_sc_hd__and3_1
X_11227_ reg_next_pc\[10\] reg_out\[10\] _05858_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__mux2_2
XANTENNA__10415__S1 _04284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11158_ net126 net112 _04668_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10109_ _04820_ _04823_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__nand2_1
XANTENNA__13436__A _04262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11089_ _05764_ _05729_ _05702_ _05682_ _05266_ _05331_ VGND VGND VPWR VPWR _05765_
+ sky130_fd_sc_hd__mux4_1
X_15966_ _03286_ _03198_ _03233_ _02674_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14482__A2 _07992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17705_ clknet_leaf_75_clk _00874_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dfxtp_1
X_14917_ net194 net163 _01824_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15897_ _03304_ is_alu_reg_imm _02610_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_19_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15651__A _03301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17636_ clknet_leaf_51_clk _00805_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfxtp_4
X_14848_ count_cycle\[49\] count_cycle\[50\] count_cycle\[51\] _01780_ VGND VGND VPWR
+ VPWR _01786_ sky130_fd_sc_hd__and4_2
XFILLER_0_81_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17567_ clknet_leaf_162_clk _00736_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14779_ count_cycle\[28\] _01736_ count_cycle\[29\] VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_82_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15982__A2 _03916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16518_ _02992_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17498_ clknet_leaf_109_clk _00667_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09661__A2 _04049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16449_ _06987_ cpuregs.regs\[29\]\[21\] _02954_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15290__S0 _02085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09795__S _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09413__A2 _04145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14714__B _08350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18119_ clknet_leaf_53_clk _01223_ VGND VGND VPWR VPWR latched_store sky130_fd_sc_hd__dfxtp_2
XFILLER_0_143_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13110__S _07068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15593__S1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16421__S _02932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16447__A0 _06984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09824__A _04231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09823_ _04545_ _04546_ _04369_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__mux2_1
XANTENNA__10192__C1 _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15345__S1 _02070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13991__D _07755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09754_ cpuregs.regs\[16\]\[10\] cpuregs.regs\[17\]\[10\] cpuregs.regs\[18\]\[10\]
+ cpuregs.regs\[19\]\[10\] _04085_ _04087_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__mux4_1
XANTENNA__12250__A _06083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08705_ net113 net81 VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__nand2_1
X_09685_ _04231_ _04408_ _04412_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13780__S _07224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_93_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10495__B1 _04100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08636_ instr_sltu instr_sltiu instr_bltu VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__or3_1
XFILLER_0_96_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10590__S0 _05239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12236__A1 _06590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08567_ irq_mask\[21\] irq_pending\[21\] VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08498_ _03277_ _03279_ _03280_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11313__B _05929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15186__B1 _01963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15281__S0 _02074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10460_ _05164_ _05165_ _04064_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08903__A _03666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09119_ mem_rdata_q\[22\] _03876_ _03846_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10391_ cpuregs.regs\[0\]\[28\] cpuregs.regs\[1\]\[28\] cpuregs.regs\[2\]\[28\] cpuregs.regs\[3\]\[28\]
+ _04273_ _04283_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12130_ _06521_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15584__S1 _01909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12061_ _06274_ cpuregs.regs\[22\]\[22\] _06482_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11012_ _05461_ _05603_ _05691_ _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__a211o_1
XANTENNA__10722__A1 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15820_ decoded_imm_j\[10\] _05974_ _02593_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__a21o_1
XANTENNA__15110__B1 decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _04979_ _02506_ _02550_ _02545_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__o211a_1
XANTENNA__11278__A2 _05829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12963_ _06996_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_84_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_2
X_14702_ count_cycle\[4\] count_cycle\[5\] _08340_ VGND VGND VPWR VPWR _08343_ sky130_fd_sc_hd__and3_1
XANTENNA__16205__A3 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18470_ clknet_leaf_140_clk _01535_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_11914_ _06406_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10486__B1 _04225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15682_ timer\[6\] _02495_ timer\[7\] VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_47_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _06949_ cpuregs.regs\[31\]\[3\] _06943_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17421_ clknet_leaf_149_clk _00590_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_47_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12227__A1 _06584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14633_ _07899_ _07964_ _08279_ _08284_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__a31o_1
XFILLER_0_158_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11845_ _06368_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_64_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output104_A net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10819__S _05287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17352_ clknet_leaf_133_clk _00521_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11504__A _06077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14564_ _08212_ VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__clkbuf_4
X_11776_ _06321_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10789__A1 _05416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16303_ _06978_ cpuregs.regs\[15\]\[17\] _02870_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13515_ _07281_ _07371_ _07282_ reg_pc\[10\] VGND VGND VPWR VPWR _07372_ sky130_fd_sc_hd__a22o_1
XANTENNA__11223__B _05860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10727_ _05254_ _05261_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__and3_1
X_17283_ clknet_leaf_126_clk _00457_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16506__S _02979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14495_ _03368_ _08153_ _08154_ _08157_ VGND VGND VPWR VPWR _08158_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15272__S0 _01973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14924__A0 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16234_ _02841_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__clkbuf_1
X_13446_ _04262_ _07307_ _07225_ VGND VGND VPWR VPWR _07308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09909__A _04227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10658_ _05225_ _05341_ _05354_ _05359_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14534__B _07944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16165_ net276 net238 _02797_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__mux2_1
X_13377_ _07242_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09628__B decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10589_ _03530_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08532__B _03311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16677__A0 _06941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15116_ _01919_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__buf_8
XFILLER_0_11_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12328_ cpuregs.regs\[26\]\[2\] _06538_ _06641_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__mux2_1
X_16096_ _03762_ _03736_ _03776_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15575__S1 _02031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15047_ _03664_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__buf_8
XFILLER_0_76_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12259_ cpuregs.regs\[25\]\[2\] _06538_ _06604_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__mux2_1
XANTENNA__14550__A _07952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15327__S1 _01997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16998_ clknet_leaf_139_clk _00172_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09867__C1 _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15949_ _02661_ _02670_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_75_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__10477__B1 _04105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09470_ _03680_ _04198_ _04201_ _03226_ _04202_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14207__A2 _07906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09882__A2 _04602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08421_ net262 net65 _03198_ mem_do_rinst VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17619_ clknet_leaf_154_clk _00788_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12218__A1 _06578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18599_ clknet_leaf_131_clk _01664_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11414__A _03215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09634__A2 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13718__A1 _04945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14915__A0 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14460__A decoded_imm_j\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13351__C1 _05260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09554__A _04284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11901__A0 _06184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09806_ count_cycle\[11\] _04165_ _04530_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__a21o_1
XANTENNA__13329__S0 _04207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15643__A1 mem_do_prefetch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16840__A0 _06554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15643__B2 _03301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11308__B _05929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09737_ _04461_ _04462_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__nand2_1
XANTENNA__12457__A1 _06598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_66_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__17921__D _08380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09668_ count_instr\[40\] _04104_ _04011_ count_instr\[8\] VGND VGND VPWR VPWR _04396_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_19_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13406__A0 _04198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08619_ irq_mask\[2\] irq_active _03248_ _03245_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__nor4b_4
XANTENNA__15946__A2 _02650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09599_ _04123_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_167_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13015__S _07021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11630_ _06186_ reg_next_pc\[12\] _06189_ _06191_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__a211o_2
XANTENNA__09086__A0 mem_rdata_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10315__S0 _04123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ _06071_ reg_next_pc\[5\] _06129_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_42_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16326__S _02881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10640__A0 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15254__S0 _01990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13300_ _06987_ cpuregs.regs\[5\]\[21\] _07176_ VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10512_ is_compare _05212_ _05213_ _05215_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__or4_1
XANTENNA__09729__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14280_ _05909_ _06301_ VGND VGND VPWR VPWR _07963_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_21_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11492_ _06065_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_21_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13231_ _07141_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__clkbuf_1
X_10443_ _05113_ _05117_ _05118_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12155__A _06095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_1014 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13162_ _06984_ cpuregs.regs\[4\]\[20\] _07104_ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__mux2_1
X_10374_ _05016_ _05019_ _05080_ _05081_ _05049_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__a311o_1
XFILLER_0_131_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12113_ _06512_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12145__A0 _06336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17970_ clknet_leaf_4_clk _01107_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dfxtp_1
X_13093_ _07045_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09010__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12044_ _06208_ cpuregs.regs\[22\]\[14\] _06471_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__mux2_1
X_16921_ clknet_leaf_172_clk _00102_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11499__A2 latched_compr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10156__C1 _04227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16852_ _06567_ cpuregs.regs\[14\]\[16\] _03163_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__mux2_1
X_15803_ decoded_imm_j\[2\] _05974_ _05982_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__a21o_1
XANTENNA_output221_A net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16783_ _03133_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13645__B1 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13995_ count_instr\[3\] _07761_ _07759_ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_57_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__15405__S _03713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15734_ timer\[19\] timer\[20\] _02533_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__or3_1
X_18522_ clknet_leaf_19_clk _01587_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12946_ _06942_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__buf_6
XANTENNA__11120__B2 _05281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15665_ timer\[2\] _02483_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_29_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18453_ clknet_leaf_14_clk _01518_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_150 net203 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12877_ _06938_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13948__A1 _03346_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17404_ clknet_leaf_100_clk _00573_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_14616_ _08221_ _08268_ VGND VGND VPWR VPWR _08269_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11828_ _06175_ cpuregs.regs\[11\]\[10\] _06359_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18384_ clknet_leaf_106_clk _01449_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15596_ decoded_imm\[29\] _02216_ _01959_ _02426_ _01934_ VGND VGND VPWR VPWR _02427_
+ sky130_fd_sc_hd__a221o_2
XANTENNA__09616__A2 _04342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17335_ clknet_leaf_177_clk _00509_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_14547_ _07943_ _07946_ _07950_ _08162_ VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__and4_1
XFILLER_0_138_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11759_ reg_pc\[27\] reg_pc\[26\] _06291_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17266_ clknet_leaf_113_clk _00440_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14478_ _08128_ _08131_ _08141_ VGND VGND VPWR VPWR _08142_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_125_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16217_ net41 mem_16bit_buffer\[1\] _02831_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13429_ _07287_ _07291_ _07289_ VGND VGND VPWR VPWR _07292_ sky130_fd_sc_hd__and3b_1
XFILLER_0_153_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17197_ clknet_leaf_121_clk _00371_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__14373__B2 _08033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16148_ net267 net229 _02786_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08970_ _03231_ _03731_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__nand2_1
X_16079_ decoded_imm\[29\] _02750_ _02746_ mem_rdata_q\[29\] _02749_ VGND VGND VPWR
+ VPWR _01342_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14676__A2 _07969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11128__B _05301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13636__A0 _04642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput1 irq[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12439__A1 _06580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__13624__A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09522_ net59 net258 _04035_ net45 _04253_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__a221o_1
XANTENNA__08718__A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08512__C1 _03294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13343__B _07209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09453_ _04185_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__inv_2
XANTENNA__15928__A2 _02617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10870__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16050__B2 _02613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08404_ reg_next_pc\[1\] _03189_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09384_ _03384_ _04116_ _04117_ _04118_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09607__A2 _04021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13403__A3 _05259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12674__S _06825_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14455__A _06860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15236__S0 _02085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09549__A _04055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11178__A1 _04038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11178__B2 _03297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09791__A1 _04289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12127__A0 _06266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14190__A _03293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09284__A instr_maskirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10090_ irq_mask\[19\] _04021_ timer\[19\] _04023_ _04026_ VGND VGND VPWR VPWR _04807_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__15616__A1 _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12849__S _06917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11753__S _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15225__S _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12800_ _06897_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13534__A _04708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13780_ _05086_ _07618_ _07224_ VGND VGND VPWR VPWR _07619_ sky130_fd_sc_hd__mux2_1
X_10992_ _05255_ _05439_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__or2b_1
X_12731_ _06858_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16041__A1 decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15450_ _02285_ _02286_ _02287_ _02288_ _02111_ _03683_ VGND VGND VPWR VPWR _02289_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12662_ _06821_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14401_ _08070_ VGND VGND VPWR VPWR _08071_ sky130_fd_sc_hd__buf_2
X_11613_ _06175_ cpuregs.regs\[10\]\[10\] _06176_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15381_ cpuregs.regs\[8\]\[17\] cpuregs.regs\[9\]\[17\] cpuregs.regs\[10\]\[17\]
+ cpuregs.regs\[11\]\[17\] _03641_ _03684_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12593_ cpuregs.regs\[2\]\[30\] _06596_ _06751_ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17120_ clknet_leaf_174_clk _00294_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10613__B1 _05205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14332_ _07901_ _07907_ decoded_imm_j\[2\] VGND VGND VPWR VPWR _08008_ sky130_fd_sc_hd__a21oi_1
X_11544_ _06114_ cpuregs.regs\[10\]\[3\] _06086_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_36_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17051_ clknet_leaf_3_clk _00225_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14263_ reg_next_pc\[20\] _05876_ _07922_ _07951_ VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__o211a_2
X_11475_ irq_mask\[25\] _03428_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__or2_1
XANTENNA__11169__A1 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16002_ _03826_ _06016_ _05996_ _06018_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__a31o_1
X_13214_ _07132_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10426_ cpuregs.regs\[4\]\[29\] cpuregs.regs\[5\]\[29\] cpuregs.regs\[6\]\[29\] cpuregs.regs\[7\]\[29\]
+ _04273_ _04469_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14194_ _03188_ _06088_ _07901_ _03190_ VGND VGND VPWR VPWR _07902_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15196__A _03709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11928__S _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13145_ _06968_ cpuregs.regs\[4\]\[12\] _07093_ VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10357_ _05064_ _05065_ _04065_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08810__B _03575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14658__A2 _07967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17953_ clknet_leaf_191_clk _01090_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dfxtp_1
X_13076_ _07059_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _04997_ _04998_ _04223_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09534__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09534__B2 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12027_ _06141_ cpuregs.regs\[22\]\[6\] _06460_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__mux2_1
X_16904_ clknet_leaf_33_clk _00049_ VGND VGND VPWR VPWR mem_rdata_q\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_100_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17884_ clknet_leaf_81_clk _01053_ VGND VGND VPWR VPWR count_cycle\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10775__S0 _05413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16835_ _06550_ cpuregs.regs\[14\]\[8\] _03152_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__mux2_1
XANTENNA__13618__B1 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12759__S _06869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13978_ _07751_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__clkbuf_1
X_16766_ _03124_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14291__B1 _07969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18505_ clknet_leaf_99_clk _01570_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15717_ _07441_ _02506_ _02525_ _02481_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__o211a_1
X_12929_ _06973_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10301__C1 _04150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16697_ _03075_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16032__A1 decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15466__S0 _02111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18436_ clknet_leaf_133_clk _01501_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15648_ _03218_ _02472_ _03291_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__a21o_1
XANTENNA__14594__A1 _07958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14594__B2 _07984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18367_ clknet_leaf_127_clk _01432_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_15579_ _02088_ _02406_ _02408_ _02410_ _02004_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__a221o_1
XANTENNA__14275__A _03294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10604__A0 _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17318_ clknet_leaf_138_clk _00492_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09470__B1 _04201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18298_ clknet_leaf_5_clk _01366_ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17249_ clknet_leaf_183_clk _00423_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_955 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09448__S1 _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10907__A1 _05361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11838__S _06359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08720__B net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14649__A2 _07967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08953_ _03683_ _03710_ _03715_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08959__S0 _03661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08884_ _03640_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10135__A2 _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14282__B1 _07964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09043__S _03730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09505_ _00073_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__buf_6
XANTENNA__11096__B1 _05390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09436_ cpuregs.regs\[28\]\[3\] cpuregs.regs\[29\]\[3\] cpuregs.regs\[30\]\[3\] cpuregs.regs\[31\]\[3\]
+ _04056_ _04091_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_502 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14034__B1 _07790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09367_ _04051_ _04101_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__nor2_1
XANTENNA__15209__S0 _01970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11399__A1 _03767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09279__A _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_50 decoded_imm\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09298_ mem_wordsize\[2\] mem_wordsize\[1\] _03242_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__o21a_2
XFILLER_0_118_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_61 net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10071__A1 _04018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_83 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 _01968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11260_ _05878_ _05881_ _05885_ _05889_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__and4b_1
XFILLER_0_105_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11020__B1 _05334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10211_ cpuregs.regs\[12\]\[23\] cpuregs.regs\[13\]\[23\] cpuregs.regs\[14\]\[23\]
+ cpuregs.regs\[15\]\[23\] _04512_ _04513_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09726__B decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11191_ _03189_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_37_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10142_ _04855_ _04856_ _04430_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__mux2_1
Xoutput190 net190 VGND VGND VPWR VPWR mem_addr[7] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14950_ _01850_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__clkbuf_1
X_10073_ cpuregs.regs\[16\]\[19\] cpuregs.regs\[17\]\[19\] cpuregs.regs\[18\]\[19\]
+ cpuregs.regs\[19\]\[19\] _04512_ _04513_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__mux4_1
XANTENNA__12520__A0 _06320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13901_ _03349_ _07678_ _07682_ net160 VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__a22o_1
X_14881_ count_cycle\[60\] count_cycle\[61\] _01801_ count_cycle\[62\] VGND VGND VPWR
+ VPWR _01808_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_50_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12579__S _06774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13832_ _07655_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__clkbuf_1
X_16620_ _03046_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14273__B1 _07958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09819__A2 _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16551_ _06953_ cpuregs.regs\[18\]\[5\] _03004_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__mux2_1
X_13763_ _07580_ _07598_ VGND VGND VPWR VPWR _07602_ sky130_fd_sc_hd__nor2_1
X_10975_ _05658_ _05633_ _05598_ _05571_ _05266_ _05395_ VGND VGND VPWR VPWR _05659_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10834__A0 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15448__S0 _01976_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15502_ cpuregs.regs\[24\]\[24\] cpuregs.regs\[25\]\[24\] cpuregs.regs\[26\]\[24\]
+ cpuregs.regs\[27\]\[24\] _02022_ _02023_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__mux4_1
X_12714_ _06274_ cpuregs.regs\[12\]\[22\] _06847_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__mux2_1
X_16482_ _02973_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__clkbuf_1
X_13694_ _05076_ _04810_ _07277_ VGND VGND VPWR VPWR _07538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18221_ clknet_leaf_41_clk _01292_ VGND VGND VPWR VPWR instr_fence sky130_fd_sc_hd__dfxtp_1
X_15433_ cpuregs.regs\[0\]\[20\] cpuregs.regs\[1\]\[20\] cpuregs.regs\[2\]\[20\] cpuregs.regs\[3\]\[20\]
+ _02085_ _02086_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12645_ _06274_ cpuregs.regs\[30\]\[22\] _06810_ VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09678__S1 _04087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18152_ clknet_leaf_45_clk alu_out\[26\] VGND VGND VPWR VPWR alu_out_q\[26\] sky130_fd_sc_hd__dfxtp_1
X_15364_ _02066_ _02207_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09452__B1 _04099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12576_ _06776_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10062__A1 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14315_ decoder_trigger _03319_ _03364_ VGND VGND VPWR VPWR _07992_ sky130_fd_sc_hd__o21ai_4
X_17103_ clknet_leaf_124_clk _00277_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_18083_ clknet_leaf_27_clk _01188_ VGND VGND VPWR VPWR mem_do_wdata sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11527_ reg_out\[2\] alu_out_q\[2\] latched_stalu VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15295_ _02066_ _02142_ _03654_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17034_ clknet_leaf_139_clk _00208_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_output96_A net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14246_ reg_pc\[15\] _07926_ _07939_ _07935_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11458_ _06041_ irq_pending\[17\] _06047_ net9 VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11658__S _06176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10409_ reg_pc\[28\] decoded_imm\[28\] _05084_ _05115_ VGND VGND VPWR VPWR _05116_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13439__A _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13551__A2 _04593_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14177_ count_instr\[59\] _07887_ _07889_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__o21a_1
X_11389_ _03756_ _03994_ _04000_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__or3_1
XANTENNA__10365__A2 _04165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15828__A1 decoded_imm_j\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09850__S1 _04513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13128_ _06951_ cpuregs.regs\[4\]\[4\] _07082_ VGND VGND VPWR VPWR _07087_ sky130_fd_sc_hd__mux2_1
XANTENNA__09507__A1 _04215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17936_ clknet_leaf_50_clk _08376_ VGND VGND VPWR VPWR reg_out\[16\] sky130_fd_sc_hd__dfxtp_1
X_13059_ _07050_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17867_ clknet_leaf_94_clk _01036_ VGND VGND VPWR VPWR count_cycle\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12489__S _06726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16253__A1 _03810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16818_ _03151_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__buf_6
XANTENNA__14264__B1 _07952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17798_ clknet_leaf_56_clk _00967_ VGND VGND VPWR VPWR reg_pc\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_105_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11406__B _03910_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16749_ _06422_ _06823_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_105_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09798__S _04321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09221_ _03786_ _03955_ _03956_ _03737_ _03963_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__a221o_1
X_18419_ clknet_leaf_162_clk _01484_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08715__B net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09152_ _03739_ _03842_ _03869_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09443__B1 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10053__A1 _04321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09994__A1 _03385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11250__B1 _05881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09994__B2 _03303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09083_ _03843_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_674 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08731__A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_171_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13542__A2 decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15819__A1 _03867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09106__C_N _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15819__B2 _04000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09985_ count_instr\[16\] _04145_ _04105_ count_cycle\[48\] VGND VGND VPWR VPWR _04705_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_129_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08936_ _03698_ _03699_ _03664_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_186_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12399__S _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08867_ _03199_ _03310_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_142_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08798_ _03490_ _03562_ _03563_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11069__A0 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09357__S0 _04056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10816__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15503__S _01984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10760_ _05456_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14007__B1 _07759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08906__A _03646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10911__S0 _05286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09419_ reg_pc\[2\] decoded_imm\[2\] VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__or2_1
X_10691_ _03542_ _05389_ _05390_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__mux2_1
XANTENNA__10647__S _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13023__S _07021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_124_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12430_ cpuregs.regs\[27\]\[18\] _06571_ _06689_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09434__B1 _04165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12361_ cpuregs.regs\[26\]\[18\] _06571_ _06652_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12862__S _06928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14100_ count_instr\[36\] count_instr\[35\] _07831_ VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__and3_1
X_11312_ _05925_ _05929_ _05932_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15602__S0 _03641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15080_ cpuregs.regs\[12\]\[1\] cpuregs.regs\[13\]\[1\] cpuregs.regs\[14\]\[1\] cpuregs.regs\[15\]\[1\]
+ _03669_ _03646_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__mux4_1
XFILLER_0_160_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12292_ cpuregs.regs\[25\]\[18\] _06571_ _06615_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_139_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14362__B _07984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14031_ _07787_ _07788_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__nor2_1
X_11243_ reg_next_pc\[13\] reg_out\[13\] _05876_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__mux2_2
XANTENNA__09832__S1 _04086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11174_ _04038_ net126 net103 _03297_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10125_ _04272_ _04836_ _04840_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__a21oi_1
X_15982_ _03743_ _03916_ _03862_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14494__B1 _07994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17721_ clknet_leaf_83_clk _00890_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dfxtp_1
XANTENNA__09596__S0 _04325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13706__B decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10056_ _04772_ _04773_ _04121_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__mux2_1
X_14933_ _01841_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15038__A2 _01865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17652_ clknet_leaf_49_clk _00821_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfxtp_2
X_14864_ _01795_ _01753_ _01796_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__and3b_1
XANTENNA__10411__A reg_pc\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15443__C1 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16603_ _07005_ cpuregs.regs\[18\]\[30\] _03003_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13815_ cpuregs.regs\[0\]\[4\] VGND VGND VPWR VPWR _07647_ sky130_fd_sc_hd__clkbuf_1
X_14795_ _01750_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__clkbuf_1
X_17583_ clknet_leaf_146_clk _00752_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15413__S _03664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13746_ _05037_ VGND VGND VPWR VPWR _07587_ sky130_fd_sc_hd__inv_2
X_16534_ _03000_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__clkbuf_1
X_10958_ _03479_ _05642_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_67_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14537__B _07950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11480__B1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13677_ _04880_ _07522_ _07374_ VGND VGND VPWR VPWR _07523_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16465_ _07003_ cpuregs.regs\[29\]\[29\] _02954_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10889_ _05348_ _05329_ _05413_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18204_ clknet_leaf_28_clk _01275_ VGND VGND VPWR VPWR instr_slli sky130_fd_sc_hd__dfxtp_2
XFILLER_0_54_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15416_ cpuregs.regs\[8\]\[19\] cpuregs.regs\[9\]\[19\] cpuregs.regs\[10\]\[19\]
+ cpuregs.regs\[11\]\[19\] _02046_ _02047_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__mux4_1
X_12628_ _06208_ cpuregs.regs\[30\]\[14\] _06799_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__mux2_1
X_16396_ _02927_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10035__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11232__A0 reg_next_pc\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18135_ clknet_leaf_50_clk alu_out\[9\] VGND VGND VPWR VPWR alu_out_q\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15649__A mem_do_wdata VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15347_ cpuregs.regs\[28\]\[15\] cpuregs.regs\[29\]\[15\] cpuregs.regs\[30\]\[15\]
+ cpuregs.regs\[31\]\[15\] _01999_ _02000_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__mux4_1
XANTENNA__12772__S _06880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12559_ _06767_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10586__A2 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12980__A0 _07007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09647__A _04124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18066_ clknet_leaf_72_clk _01171_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_2
X_15278_ cpuregs.regs\[20\]\[11\] cpuregs.regs\[21\]\[11\] cpuregs.regs\[22\]\[11\]
+ cpuregs.regs\[23\]\[11\] _02069_ _02070_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__mux4_1
XFILLER_0_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14229_ reg_next_pc\[10\] _05858_ _07922_ _07927_ VGND VGND VPWR VPWR _07928_ sky130_fd_sc_hd__o211a_2
XFILLER_0_1_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17017_ clknet_leaf_172_clk _00191_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09770_ count_instr\[42\] instr_rdinstrh instr_rdinstr count_instr\[10\] VGND VGND
+ VPWR VPWR _04496_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08721_ net107 net75 VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__and2_1
X_17919_ clknet_leaf_69_clk _01088_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_107_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15029__A2 _01863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11417__A _03215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13108__S _07068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08652_ timer\[13\] timer\[12\] timer\[15\] timer\[14\] VGND VGND VPWR VPWR _03419_
+ sky130_fd_sc_hd__or4_1
XANTENNA__15649__D_N _07904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08583_ irq_active irq_delay VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__nor2_1
XANTENNA__16419__S _02932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12947__S _06985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11851__S _06370_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08726__A net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08445__B mem_do_prefetch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09204_ _03885_ _03845_ _03948_ _03826_ _03949_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09135_ _03774_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_162_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12682__S _06825_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14463__A decoded_imm_j\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10577__A2 _05219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09431__A3 _04164_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10121__S1 _04285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09066_ mem_rdata_q\[24\] net49 _03227_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09719__A1 _04206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15060__S1 _01919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13515__A2 _07371_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10329__A2 _04448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__17924__D _08395_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08942__A2 _03703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09968_ _04686_ _04687_ _04575_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__mux2_1
X_08919_ _03654_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__buf_6
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09899_ _04328_ _04620_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11930_ _06297_ cpuregs.regs\[20\]\[25\] _06409_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15976__A0 instr_waitirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11861_ _06304_ cpuregs.regs\[11\]\[26\] _06370_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13600_ _04848_ _05227_ VGND VGND VPWR VPWR _07451_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10812_ _05278_ _05349_ _05228_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _07954_ _07956_ _08209_ VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _06335_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13531_ _04532_ _07386_ _07374_ VGND VGND VPWR VPWR _07387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10265__A1 _04068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10743_ net95 _03524_ _03609_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__mux2_1
XANTENNA__11462__B1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12158__A _06104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16250_ _02849_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__clkbuf_1
X_13462_ _07313_ _07314_ _07320_ _07322_ VGND VGND VPWR VPWR _07323_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_45_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10674_ _05370_ _05372_ _05373_ _05374_ _05243_ _05244_ VGND VGND VPWR VPWR _05375_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10017__A1 _04070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15201_ cpuregs.regs\[24\]\[7\] cpuregs.regs\[25\]\[7\] cpuregs.regs\[26\]\[7\] cpuregs.regs\[27\]\[7\]
+ _03661_ _03662_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_62_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11214__B1 _05851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12413_ _06677_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13754__A2 _05261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14951__A1 net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16181_ net284 net246 _02770_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__mux2_1
XANTENNA__09502__S0 _04232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13393_ _04160_ _07257_ _07225_ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15132_ cpuregs.regs\[28\]\[5\] cpuregs.regs\[29\]\[5\] cpuregs.regs\[30\]\[5\] cpuregs.regs\[31\]\[5\]
+ _01985_ _01986_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__mux4_1
XANTENNA__09467__A _04036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12344_ _06640_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__buf_6
XFILLER_0_105_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_1018 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15063_ _01907_ _01920_ _01922_ _03654_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__o211a_1
XANTENNA__15051__S1 _03659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12275_ _06603_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10406__A reg_pc\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14014_ count_instr\[9\] _07773_ _07776_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__o21a_1
X_11226_ _05838_ _05861_ _05862_ _05863_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__o31ai_4
XANTENNA__11936__S _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13717__A _05086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11157_ _05813_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10108_ _04820_ _04823_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__or2_1
XANTENNA__09569__S0 _04275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09406__S _04077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13436__B decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11088_ _05086_ _05076_ _05237_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__mux2_1
X_15965_ _02685_ _02678_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__or2_1
XANTENNA__16208__A1 _06082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17704_ clknet_leaf_75_clk _00873_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10039_ count_instr\[18\] _04012_ count_cycle\[18\] _04165_ _04756_ VGND VGND VPWR
+ VPWR _04757_ sky130_fd_sc_hd__a221o_1
X_14916_ _01832_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_69_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14219__B1 _07901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13690__A1 _07232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15896_ _02612_ _03940_ _02613_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_19_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17635_ clknet_leaf_51_clk _00804_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dfxtp_4
XANTENNA__15651__B _04187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14847_ _01785_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_102_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14548__A _07988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17566_ clknet_leaf_125_clk _00735_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_14778_ count_cycle\[28\] _01736_ _01738_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16517_ cpuregs.regs\[17\]\[21\] _06578_ _02990_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__mux2_1
X_13729_ _07555_ _07558_ _07569_ VGND VGND VPWR VPWR _07571_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17497_ clknet_leaf_114_clk _00666_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16448_ _02955_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_30_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09949__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15290__S1 _02086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15379__A _03659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16379_ _06984_ cpuregs.regs\[16\]\[20\] _02918_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18118_ clknet_leaf_63_clk _01222_ VGND VGND VPWR VPWR irq_state\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18049_ clknet_leaf_45_clk _01154_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_41_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16702__S _03087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12007__S _06446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12705__A0 _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11846__S _06359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09822_ cpuregs.regs\[12\]\[12\] cpuregs.regs\[13\]\[12\] cpuregs.regs\[14\]\[12\]
+ cpuregs.regs\[15\]\[12\] _04085_ _04087_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09753_ cpuregs.regs\[20\]\[10\] cpuregs.regs\[21\]\[10\] cpuregs.regs\[22\]\[10\]
+ cpuregs.regs\[23\]\[10\] _04477_ _04478_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__mux4_1
X_08704_ net113 net81 VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__or2_1
XANTENNA__10051__A _04430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09684_ _04069_ _04411_ _04081_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08635_ _03405_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13362__A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10590__S1 _05237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08566_ _03341_ _03342_ _03343_ _03344_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13433__A1 _04342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08456__A _03239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14630__B1 _08097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11444__B1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08497_ mem_do_wdata _03278_ cpu_state\[5\] VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10798__A2 _04419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15186__A1 decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11313__C _05932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15281__S1 _02075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09287__A _04023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09118_ _03850_ _03795_ _03796_ _03849_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10390_ cpuregs.regs\[4\]\[28\] cpuregs.regs\[5\]\[28\] cpuregs.regs\[6\]\[28\] cpuregs.regs\[7\]\[28\]
+ _04290_ _04283_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_40_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09049_ net42 mem_rdata_q\[18\] _03729_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__mux2_1
XANTENNA__14921__A _01823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12060_ _06484_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__clkbuf_1
X_11011_ _03468_ _05440_ _05646_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10722__A2 _04262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15110__B2 _01932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ timer\[24\] _02547_ _02549_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__o21ai_1
X_12962_ _06995_ cpuregs.regs\[31\]\[25\] _06985_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__mux2_1
XANTENNA__13672__A1 _04744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11132__C1 _05251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14701_ count_cycle\[4\] _08340_ _08342_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__o21a_1
X_11913_ _06232_ cpuregs.regs\[20\]\[17\] _06398_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__mux2_1
XANTENNA__09750__A _04054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10486__A1 _04206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09971__S0 _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12893_ _06113_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12587__S _06774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15681_ _02477_ _02497_ _02498_ _02481_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ clknet_leaf_162_clk _00589_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_47_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _06240_ cpuregs.regs\[11\]\[18\] _06359_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__mux2_1
X_14632_ reg_next_pc\[26\] _07947_ _08283_ _08033_ VGND VGND VPWR VPWR _08284_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17351_ clknet_leaf_182_clk _00520_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_14563_ _08198_ _08213_ VGND VGND VPWR VPWR _08220_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11775_ _06320_ cpuregs.regs\[10\]\[28\] _06258_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16302_ _02877_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10726_ _05422_ _05424_ _03530_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13514_ _04493_ VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__inv_2
XANTENNA__16374__A0 _06980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17282_ clknet_leaf_175_clk _00456_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_14494_ _07986_ _08155_ _08156_ _07994_ _07939_ VGND VGND VPWR VPWR _08157_ sky130_fd_sc_hd__a32o_1
XFILLER_0_138_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13188__A0 _06941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output299_A net299 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13445_ _07191_ _07295_ _07303_ _07306_ VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__o31a_1
XFILLER_0_36_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15272__S1 _01974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16233_ net50 mem_16bit_buffer\[9\] _02831_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__mux2_1
XANTENNA__10835__S _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10657_ _05355_ _05222_ _05301_ _03532_ _05358_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09909__B _04630_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13211__S _07129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13376_ _04040_ _07241_ _07225_ VGND VGND VPWR VPWR _07242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16164_ _02800_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__clkbuf_1
X_10588_ _05289_ _05290_ _05242_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12327_ _06643_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__clkbuf_1
X_15115_ _01918_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__buf_8
XFILLER_0_23_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16095_ _03309_ _06006_ _02758_ _06026_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__o211a_1
X_15046_ _01905_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__buf_4
XFILLER_0_121_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09925__A _04483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12258_ _06606_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11209_ _05844_ _05848_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12189_ _06192_ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__buf_2
XANTENNA__15637__C1 _03277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16997_ clknet_leaf_157_clk _00171_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_15948_ mem_rdata_q\[5\] mem_rdata_q\[4\] mem_rdata_q\[6\] mem_rdata_q\[3\] VGND
+ VGND VPWR VPWR _02670_ sky130_fd_sc_hd__or4b_1
XANTENNA__14860__B1 _01714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12497__S _06726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15879_ decoder_pseudo_trigger decoder_trigger VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__or2b_1
XANTENNA__14278__A _03293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08420_ mem_16bit_buffer\[0\] _03204_ _03205_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__mux2_2
X_17618_ clknet_leaf_140_clk _00787_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18598_ clknet_leaf_129_clk _01663_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10229__B2 instr_timer VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17549_ clknet_leaf_145_clk _00718_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16493__A _02967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13910__A _07677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10401__A1 instr_retirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16432__S _02943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14679__B1 _08033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13351__B1 _07217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15891__A2 _02635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13367__A1_N _03387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09805_ count_instr\[11\] _04011_ _03252_ _04529_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__a211o_1
XANTENNA__10260__S0 _04329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13329__S1 _04208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14446__A3 _08050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09736_ reg_pc\[10\] decoded_imm\[10\] VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__or2_1
XANTENNA__14851__B1 _01714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09667_ _04356_ _04359_ _04392_ _04393_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_173_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08618_ mem_do_wdata _03218_ _03244_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__o21ai_1
X_09598_ _04052_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__buf_4
XANTENNA__14603__B1 _07944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08549_ irq_mask\[30\] irq_pending\[30\] VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__and2b_1
XFILLER_0_65_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09086__A1 _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15511__S _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10315__S1 _04124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11560_ irq_state\[1\] _03322_ _06098_ _06128_ _06074_ VGND VGND VPWR VPWR _06129_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_42_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10511_ _05214_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15254__S1 _01992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11491_ latched_branch latched_store VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_80_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _06984_ cpuregs.regs\[8\]\[20\] _07140_ VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__mux2_1
X_10442_ _05146_ _05147_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16659__A1 _06288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15747__A _02476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13590__B1 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13161_ _07081_ VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__clkbuf_8
X_10373_ _05017_ _05050_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12870__S _06928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14651__A _07966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12112_ _06208_ cpuregs.regs\[23\]\[14\] _06507_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__mux2_1
X_13092_ _07067_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12043_ _06475_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__clkbuf_1
X_16920_ clknet_leaf_180_clk _00101_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09010__A1 mem_rdata_q\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16851_ _03169_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10251__S0 _04217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15802_ decoded_imm_j\[1\] _05974_ _05978_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__a21o_1
XANTENNA__13645__A1 _03631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16782_ _06565_ cpuregs.regs\[13\]\[15\] _03127_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09849__B1 _04014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13994_ count_instr\[3\] _07761_ VGND VGND VPWR VPWR _07763_ sky130_fd_sc_hd__and2_1
XANTENNA__14842__B1 _01714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10003__S0 _04057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18521_ clknet_leaf_2_clk _01586_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_15733_ timer\[19\] _02533_ timer\[20\] VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__o21a_1
X_12945_ _06256_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__buf_2
XANTENNA_output214_A net214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13206__S _07118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12110__S _06507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18452_ clknet_leaf_177_clk _01517_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_15664_ _02484_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12876_ _06328_ cpuregs.regs\[6\]\[29\] _06928_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_151 net203 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17403_ clknet_leaf_166_clk _00572_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_14615_ _07942_ _07961_ VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11827_ _06347_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__clkbuf_8
X_18383_ clknet_leaf_166_clk _01448_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15595_ _02416_ _02419_ _02422_ _02425_ _01968_ _02037_ VGND VGND VPWR VPWR _02426_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__16517__S _02990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13730__A _03275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15421__S _03653_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17334_ clknet_leaf_128_clk _00508_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08824__A1 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11758_ _06305_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__clkbuf_1
X_14546_ _07898_ _07950_ _07997_ _08204_ VGND VGND VPWR VPWR _08205_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10092__C1 _03302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10709_ _05361_ _05392_ _05393_ _05408_ VGND VGND VPWR VPWR alu_out\[4\] sky130_fd_sc_hd__a31o_1
XFILLER_0_71_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17265_ clknet_leaf_160_clk _00439_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08770__A_N net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11689_ _06242_ _06243_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__nor2_1
X_14477_ _08139_ _08140_ VGND VGND VPWR VPWR _08141_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16216_ _02832_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13428_ _07288_ VGND VGND VPWR VPWR _07291_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14373__A2 _07947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17196_ clknet_leaf_151_clk _00370_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15657__A _07778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13359_ _04037_ _07219_ _07225_ VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__mux2_1
XANTENNA__12780__S _06880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16147_ _02791_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10934__A2 instr_slli VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10490__S0 _04329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16078_ decoded_imm\[28\] _02750_ _02746_ mem_rdata_q\[28\] _02749_ VGND VGND VPWR
+ VPWR _01341_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_110_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14676__A3 _08050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15029_ irq_mask\[24\] _01863_ _01714_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__a21o_1
XANTENNA__10147__B1 _04296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15086__B1 _00068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15181__S0 _01985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput2 irq[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
XANTENNA__13636__A1 _04945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14833__B1 _01717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09521_ _04036_ mem_wordsize\[1\] _04252_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13624__B decoded_imm\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08718__B net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13116__S _07045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11425__A _03305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09452_ _04172_ _04176_ _04099_ _04184_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__a211o_4
XFILLER_0_149_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08403_ latched_branch latched_store VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__and2_2
XFILLER_0_137_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16050__A2 decoded_imm_j\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10870__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09383_ _04040_ _03312_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__and2_1
XANTENNA__09068__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13640__A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08815__A1 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08734__A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15236__S1 _02086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14665__A1_N _08012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11178__A2 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14471__A _07934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09565__A _04237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10138__B1 _04012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14824__B1 _01717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08909__A _00068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09504__S _04121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11638__B1 _06066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09719_ _04206_ _04441_ _04445_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__a21o_1
XANTENNA__09926__S0 _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10991_ _05219_ _05666_ _05673_ VGND VGND VPWR VPWR alu_out\[21\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13026__S _07032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12730_ _06336_ cpuregs.regs\[12\]\[30\] _06824_ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16041__A2 _02711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12661_ _06336_ cpuregs.regs\[30\]\[30\] _06787_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_723 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16337__S _02896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11612_ _06085_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__clkbuf_8
X_14400_ _03368_ _03378_ VGND VGND VPWR VPWR _08070_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08806__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15380_ cpuregs.regs\[12\]\[17\] cpuregs.regs\[13\]\[17\] cpuregs.regs\[14\]\[17\]
+ cpuregs.regs\[15\]\[17\] _02221_ _02222_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__mux4_1
X_12592_ _06784_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11543_ _06113_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__buf_2
X_14331_ decoded_imm_j\[2\] _07900_ _07907_ VGND VGND VPWR VPWR _08007_ sky130_fd_sc_hd__and3_1
XANTENNA__09459__B decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14262_ _05857_ _06254_ VGND VGND VPWR VPWR _07951_ sky130_fd_sc_hd__or2_1
X_17050_ clknet_leaf_190_clk _00224_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11474_ _06054_ irq_pending\[24\] _06056_ net17 VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__a31o_1
XFILLER_0_162_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11169__A2 _04710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13563__A0 _04602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12366__A1 _06575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13213_ _06968_ cpuregs.regs\[8\]\[12\] _07129_ VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__mux2_1
X_16001_ cpuregs.raddr1\[1\] _06006_ _06014_ _06015_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10425_ _05130_ _05131_ _04430_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14193_ _07900_ VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10377__B1 _04156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14381__A decoded_imm_j\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13144_ _07095_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09475__A _04072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10356_ cpuregs.regs\[8\]\[27\] cpuregs.regs\[9\]\[27\] cpuregs.regs\[10\]\[27\]
+ cpuregs.regs\[11\]\[27\] _04057_ _04060_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08990__A0 mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17952_ clknet_leaf_191_clk _01089_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dfxtp_1
X_13075_ _06966_ cpuregs.regs\[7\]\[11\] _07057_ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__mux2_1
XANTENNA__10129__B1 _04105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10287_ cpuregs.regs\[24\]\[25\] cpuregs.regs\[25\]\[25\] cpuregs.regs\[26\]\[25\]
+ cpuregs.regs\[27\]\[25\] _04291_ _04292_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_72_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12026_ _06466_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16903_ clknet_leaf_33_clk _00048_ VGND VGND VPWR VPWR mem_rdata_q\[22\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__11229__B _05864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09534__A2 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17883_ clknet_leaf_89_clk _01052_ VGND VGND VPWR VPWR count_cycle\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10614__B_N _05205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10775__S1 _05414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13725__A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16834_ _03160_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13618__A1 _07304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14815__B1 _01717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11629__B1 _06066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16765_ _06548_ cpuregs.regs\[13\]\[7\] _03116_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__mux2_1
X_13977_ _07737_ _07750_ VGND VGND VPWR VPWR _07751_ sky130_fd_sc_hd__and2_1
XANTENNA__14291__B2 _07960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18504_ clknet_leaf_151_clk _01569_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15716_ _02476_ _02523_ _02524_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__or3b_1
XFILLER_0_88_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12928_ _06972_ cpuregs.regs\[31\]\[14\] _06964_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__mux2_1
X_16696_ _03086_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16032__A2 _02634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18435_ clknet_leaf_145_clk _01500_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15466__S1 _02004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15647_ _03309_ _03411_ _03630_ _07905_ _02473_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__a41o_1
XFILLER_0_69_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12859_ _06929_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13460__A _03387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14594__A2 _07994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18366_ clknet_leaf_185_clk _01431_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15791__A1 is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15578_ _03687_ _02409_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10604__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17317_ clknet_leaf_148_clk _00491_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14529_ _08187_ _08188_ VGND VGND VPWR VPWR _08189_ sky130_fd_sc_hd__or2b_1
XANTENNA__09470__A1 _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18297_ clknet_leaf_5_clk _01365_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dfxtp_1
XANTENNA__09470__B2 _03226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17248_ clknet_leaf_175_clk _00422_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17179_ clknet_leaf_12_clk _00353_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09222__B2 _03888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16710__S _03087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08952_ _03657_ _03714_ _03692_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__a21o_1
XANTENNA__12015__S _06460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10215__S0 _04472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08959__S1 _03662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08883_ cpuregs.regs\[0\]\[2\] cpuregs.regs\[1\]\[2\] cpuregs.regs\[2\]\[2\] cpuregs.regs\[3\]\[2\]
+ _03645_ _03647_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__mux4_1
XFILLER_0_138_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16011__A instr_jalr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08729__A net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14806__B1 _01717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14282__A1 reg_pc\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14282__B2 _07960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09504_ _04234_ _04235_ _04121_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09435_ instr_retirq VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_140_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10994__A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09366_ _04067_ _04083_ _04097_ _04100_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__a211o_4
XFILLER_0_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08464__A net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15209__S1 _01971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09297_ net67 VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__inv_2
XANTENNA_40 _05923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08895__S0 _03658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_51 decoded_imm\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_84 net200 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_95 _02349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10210_ _04105_ count_cycle\[55\] _04013_ count_cycle\[23\] _04922_ VGND VGND VPWR
+ VPWR _04923_ sky130_fd_sc_hd__a221o_1
XANTENNA__11020__A1 _05244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11190_ _04198_ _05829_ _05833_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__o21a_4
XTAP_TAPCELL_ROW_37_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10141_ cpuregs.regs\[12\]\[21\] cpuregs.regs\[13\]\[21\] cpuregs.regs\[14\]\[21\]
+ cpuregs.regs\[15\]\[21\] _04282_ _04285_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput180 net180 VGND VGND VPWR VPWR mem_addr[27] sky130_fd_sc_hd__clkbuf_1
Xoutput191 net191 VGND VGND VPWR VPWR mem_addr[8] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10072_ cpuregs.regs\[20\]\[19\] cpuregs.regs\[21\]\[19\] cpuregs.regs\[22\]\[19\]
+ cpuregs.regs\[23\]\[19\] _04512_ _04513_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__mux4_1
X_13900_ _07697_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__clkbuf_1
X_14880_ count_cycle\[61\] count_cycle\[62\] _01804_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_50_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13831_ cpuregs.regs\[0\]\[12\] VGND VGND VPWR VPWR _07655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15470__B1 _03692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11087__A1 _05414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16550_ _03009_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13762_ _05076_ _07271_ _07597_ _07601_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__o22a_1
X_10974_ _04848_ _04810_ _05236_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15501_ cpuregs.regs\[28\]\[24\] cpuregs.regs\[29\]\[24\] cpuregs.regs\[30\]\[24\]
+ cpuregs.regs\[31\]\[24\] _01990_ _01992_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__mux4_1
XANTENNA__10834__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12713_ _06849_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15448__S1 _01977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16481_ cpuregs.regs\[17\]\[4\] _06542_ _02968_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__mux2_1
XANTENNA__12595__S _06751_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13693_ _04913_ _05261_ _07495_ _07279_ VGND VGND VPWR VPWR _07537_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18220_ clknet_leaf_92_clk _01291_ VGND VGND VPWR VPWR instr_rdinstrh sky130_fd_sc_hd__dfxtp_2
XFILLER_0_167_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15432_ cpuregs.regs\[4\]\[20\] cpuregs.regs\[5\]\[20\] cpuregs.regs\[6\]\[20\] cpuregs.regs\[7\]\[20\]
+ _01976_ _01977_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__mux4_1
X_12644_ _06812_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12587__A1 _06590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18151_ clknet_leaf_51_clk alu_out\[25\] VGND VGND VPWR VPWR alu_out_q\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15363_ cpuregs.regs\[8\]\[16\] cpuregs.regs\[9\]\[16\] cpuregs.regs\[10\]\[16\]
+ cpuregs.regs\[11\]\[16\] _01990_ _01992_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12575_ cpuregs.regs\[2\]\[21\] _06578_ _06774_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08886__S0 _03649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17102_ clknet_leaf_122_clk _00276_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_14314_ decoded_imm_j\[1\] _07972_ _07990_ VGND VGND VPWR VPWR _07991_ sky130_fd_sc_hd__a21oi_1
X_11526_ _06065_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__clkbuf_4
X_18082_ clknet_leaf_39_clk _01187_ VGND VGND VPWR VPWR mem_do_rdata sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15294_ cpuregs.regs\[24\]\[12\] cpuregs.regs\[25\]\[12\] cpuregs.regs\[26\]\[12\]
+ cpuregs.regs\[27\]\[12\] _02069_ _02070_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17033_ clknet_leaf_141_clk _00207_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10843__S _05390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11457_ irq_mask\[17\] _06042_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__or2_1
X_14245_ reg_next_pc\[15\] _05858_ _07922_ _07938_ VGND VGND VPWR VPWR _07939_ sky130_fd_sc_hd__o211a_2
XANTENNA__09204__A1 _03885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09204__B2 _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10408_ _05113_ _05114_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__and2_1
XANTENNA__15000__A _04227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14176_ count_instr\[59\] _07887_ _07826_ VGND VGND VPWR VPWR _07889_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output89_A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11388_ _03800_ _03804_ _05997_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__or3_1
XFILLER_0_110_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10339_ _05018_ _05019_ _05016_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__o21ai_1
X_13127_ _07086_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15384__S0 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17935_ clknet_leaf_68_clk _08375_ VGND VGND VPWR VPWR reg_out\[15\] sky130_fd_sc_hd__dfxtp_1
X_13058_ _06949_ cpuregs.regs\[7\]\[3\] _07046_ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__mux2_1
XANTENNA__13455__A _04466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12009_ _06336_ cpuregs.regs\[21\]\[30\] _06423_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__mux2_1
X_17866_ clknet_leaf_94_clk _01035_ VGND VGND VPWR VPWR count_cycle\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16817_ _06080_ _06823_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__nand2_4
X_17797_ clknet_leaf_57_clk _00966_ VGND VGND VPWR VPWR reg_pc\[5\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__15461__B1 _02298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11078__A1 _05323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16748_ _03114_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_105_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11406__C _06003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16679_ _06945_ cpuregs.regs\[19\]\[1\] _03076_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09220_ _03957_ _03962_ _03932_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18418_ clknet_leaf_127_clk _01483_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11703__A _06256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09151_ mem_rdata_q\[15\] _03781_ _03846_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__mux2_1
XANTENNA__11422__B _03308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18349_ clknet_leaf_33_clk _01417_ VGND VGND VPWR VPWR mem_rdata_q\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09443__A1 _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_923 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09082_ _03743_ _03781_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11849__S _06370_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_978 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput60 mem_rdata[5] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_1
XFILLER_0_82_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08731__B net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11538__C1 _06101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_55_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15819__A2 _06016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16440__S _02943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09984_ irq_mask\[16\] _04022_ timer\[16\] _04024_ _04027_ VGND VGND VPWR VPWR _04704_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__15375__S0 _01908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08935_ cpuregs.regs\[16\]\[3\] cpuregs.regs\[17\]\[3\] cpuregs.regs\[18\]\[3\] cpuregs.regs\[19\]\[3\]
+ _03658_ _03659_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__mux4_1
XANTENNA__11584__S _06086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15056__S _03664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08866_ _03309_ _03384_ _03305_ _03631_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_142_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08797_ net105 net73 VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__and2b_1
XFILLER_0_165_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16676__A _03075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14255__B2 reg_next_pc\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11069__A1 _05044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09357__S1 _04091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10816__A1 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15204__B1 _03675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10911__S1 _05413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13304__S _07176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09418_ reg_pc\[2\] decoded_imm\[2\] VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10690_ _05323_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__buf_4
XANTENNA__15755__A1 _05009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09434__A1 _04018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09349_ _00069_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__buf_8
XFILLER_0_124_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16615__S _03040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15839__A_N _03878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12360_ _06660_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09985__A2 _04145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13518__A0 _04466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11311_ reg_next_pc\[26\] reg_out\[26\] _05928_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__mux2_2
XFILLER_0_133_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15602__S1 _03684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10663__S _05363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12291_ _06623_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_91_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14030_ count_instr\[14\] _07784_ _07759_ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_73_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11242_ _05858_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10427__S0 _04487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11173_ net119 _04710_ _05821_ VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__a21o_2
XFILLER_0_38_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10124_ _04215_ _04839_ _04225_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15981_ _03783_ _02696_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14494__A1 _07986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17720_ clknet_leaf_77_clk _00889_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dfxtp_1
X_10055_ cpuregs.regs\[8\]\[18\] cpuregs.regs\[9\]\[18\] cpuregs.regs\[10\]\[18\]
+ cpuregs.regs\[11\]\[18\] _04477_ _04478_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__mux4_1
X_14932_ net201 net170 _01835_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__mux2_1
XANTENNA__09596__S1 _04277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17651_ clknet_leaf_49_clk _00820_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dfxtp_2
X_14863_ count_cycle\[55\] _01792_ count_cycle\[56\] VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__a21o_1
XANTENNA__10411__B decoded_imm\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output127_A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16602_ _03036_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_82_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13814_ _07646_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17582_ clknet_leaf_138_clk _00751_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15994__A1 _03867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14794_ _01748_ _08350_ _01749_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__and3b_1
X_16533_ cpuregs.regs\[17\]\[29\] _06594_ _02990_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13745_ _07254_ _07584_ _07585_ _07216_ VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_67_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10957_ _05640_ _05641_ _05517_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11523__A _06095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12009__A0 _06336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11480__A1 _06054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16464_ _02963_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__clkbuf_1
X_13676_ _07191_ _07516_ _07518_ _07520_ _07521_ VGND VGND VPWR VPWR _07522_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_14_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10888_ _05399_ _05574_ _05577_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_73_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18203_ clknet_leaf_29_clk _01274_ VGND VGND VPWR VPWR instr_sw sky130_fd_sc_hd__dfxtp_1
X_15415_ _03719_ _02255_ _00067_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12627_ _06803_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__clkbuf_1
X_16395_ _07001_ cpuregs.regs\[16\]\[28\] _02918_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16525__S _02990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10035__A2 _04710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18134_ clknet_leaf_42_clk alu_out\[8\] VGND VGND VPWR VPWR alu_out_q\[8\] sky130_fd_sc_hd__dfxtp_1
X_15346_ _02012_ _02190_ _02005_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12558_ cpuregs.regs\[2\]\[13\] _06561_ _06763_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13509__B1 _03311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10586__A3 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18065_ clknet_leaf_72_clk _01170_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfxtp_4
XANTENNA__16471__D _06081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11509_ latched_branch latched_store _03195_ _03293_ VGND VGND VPWR VPWR _06083_
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15277_ _02066_ _02125_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__or2_1
XANTENNA__16171__A1 net241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08551__B irq_pending\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12489_ _06201_ cpuregs.regs\[28\]\[13\] _06726_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10991__B1 _05673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17016_ clknet_leaf_169_clk _00190_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_14228_ _05856_ _06168_ VGND VGND VPWR VPWR _07927_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14159_ count_instr\[53\] _07874_ _07877_ VGND VGND VPWR VPWR _07878_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10743__A0 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09663__A _03385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08720_ net107 net75 VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__nor2_1
X_17918_ clknet_leaf_81_clk _01087_ VGND VGND VPWR VPWR count_cycle\[63\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_107_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09361__B1 _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08651_ timer\[21\] timer\[20\] timer\[23\] timer\[22\] VGND VGND VPWR VPWR _03418_
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_124_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17849_ clknet_leaf_108_clk _01018_ VGND VGND VPWR VPWR reg_next_pc\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08582_ _03345_ _03350_ _03355_ _03360_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__or4_2
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09602__S _04222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12799__A1 _06586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09113__B1 _03810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08726__B net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13124__S _07082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09203_ _03748_ _03879_ _03878_ _03844_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09134_ _03743_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09838__A _04561_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14463__B _07934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09065_ _03762_ _03774_ _03822_ _03826_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__or4_1
XFILLER_0_130_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08461__B _03244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15370__C1 _02020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13794__S _07224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15348__S0 _02074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09967_ cpuregs.regs\[24\]\[16\] cpuregs.regs\[25\]\[16\] cpuregs.regs\[26\]\[16\]
+ cpuregs.regs\[27\]\[16\] _04281_ _04470_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__mux4_1
XANTENNA__12487__A0 _06193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08918_ reg_sh\[2\] _03638_ _03682_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__a21oi_1
X_09898_ _04618_ _04619_ _04222_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__mux2_1
X_08849_ _03613_ _03614_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__nor2_1
XANTENNA__15425__B1 _03675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11860_ _06376_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15520__S0 _02111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10811_ _03507_ _05504_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_0_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _06116_ reg_next_pc\[30\] _06332_ _06334_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__a211o_4
XTAP_TAPCELL_ROW_0_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09655__B2 _04023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13034__S _07032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13530_ _03276_ _07380_ _07384_ _07385_ VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__a22o_1
X_10742_ _05398_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10673_ _04360_ _04456_ _04419_ _04466_ _05235_ _05237_ VGND VGND VPWR VPWR _05374_
+ sky130_fd_sc_hd__mux4_1
X_13461_ reg_pc\[6\] _07211_ _07321_ _07221_ VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__a211o_1
XANTENNA__16345__S _02896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09407__B2 _04052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_173_Right_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15200_ _02051_ _02052_ _03719_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12412_ _06688_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_62_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10648__S0 _05239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16180_ _02808_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09502__S1 _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13392_ _03276_ _07248_ _07249_ _07256_ VGND VGND VPWR VPWR _07257_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15131_ _03647_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__buf_6
XFILLER_0_90_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12343_ _06651_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15587__S0 _03641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12274_ _06614_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__clkbuf_1
X_15062_ _03666_ _01921_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10406__B decoded_imm\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11225_ _04456_ _05838_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__nand2_1
X_14013_ count_instr\[9\] _07773_ _07775_ VGND VGND VPWR VPWR _07776_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15339__S0 _02030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12902__A _06140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09483__A _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11156_ _05254_ net111 _04668_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__mux2_1
XANTENNA__13717__B _05227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output244_A net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10107_ _04821_ _04822_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__nand2_1
XANTENNA__13209__S _07129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11518__A latched_compr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11087_ _05414_ _05404_ _05545_ _05602_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__a211o_1
X_15964_ net224 VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__inv_2
XANTENNA__09569__S1 _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13675__C1 _07283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17703_ clknet_leaf_75_clk _00872_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dfxtp_1
XANTENNA__16208__A2 _06862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10038_ count_instr\[50\] _04104_ _04105_ count_cycle\[50\] VGND VGND VPWR VPWR _04756_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14915_ net223 net192 _01824_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__mux2_1
XANTENNA__11150__A0 _05286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11237__B _05864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15895_ is_alu_reg_imm _02611_ _02615_ _02616_ instr_addi VGND VGND VPWR VPWR _01268_
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_69_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15424__S _03713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17634_ clknet_leaf_52_clk _00803_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dfxtp_4
X_14846_ _01783_ _01753_ _01784_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__and3b_1
XFILLER_0_59_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17565_ clknet_leaf_113_clk _00734_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14777_ count_cycle\[28\] _01736_ _01717_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_170_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11989_ _06257_ cpuregs.regs\[21\]\[20\] _06446_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16516_ _02991_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__clkbuf_1
X_13728_ _07555_ _07558_ _07569_ VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__nand3_1
XFILLER_0_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17496_ clknet_leaf_165_clk _00665_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16447_ _06984_ cpuregs.regs\[29\]\[20\] _02954_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__mux2_1
X_13659_ _07488_ _07502_ _07504_ _07505_ VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__and4_1
XFILLER_0_155_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_185_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16378_ _02895_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__buf_6
XFILLER_0_60_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18117_ clknet_leaf_63_clk _01221_ VGND VGND VPWR VPWR irq_state\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15329_ cpuregs.regs\[12\]\[14\] cpuregs.regs\[13\]\[14\] cpuregs.regs\[14\]\[14\]
+ cpuregs.regs\[15\]\[14\] _02069_ _02070_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16144__A1 net227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14155__B1 _07834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18048_ clknet_leaf_51_clk _01153_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_112_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09821_ cpuregs.regs\[8\]\[12\] cpuregs.regs\[9\]\[12\] cpuregs.regs\[10\]\[12\]
+ cpuregs.regs\[11\]\[12\] _04085_ _04087_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_129_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14458__A1 _08071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10192__B2 _04052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12023__S _06460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09752_ _04086_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_123_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08703_ _03467_ _03468_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__and2_1
X_09683_ _04409_ _04410_ _04064_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__mux2_1
XANTENNA__11141__B1 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08634_ instr_slt instr_slti instr_blt VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15502__S0 _02022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08737__A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_138_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13362__B decoded_imm\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08565_ irq_mask\[3\] irq_pending\[3\] VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__and2b_2
XFILLER_0_162_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12641__A0 _06257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08496_ _03218_ _03278_ cpu_state\[6\] VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13789__S _05227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12693__S _06836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15186__A2 _02009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_170_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_170_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_137_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09496__S0 _04207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09117_ _03855_ _03873_ _03875_ _03861_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16135__A1 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10507__A _05209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15569__S0 _01973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11102__S _05413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09048_ _03728_ _03806_ _03808_ _03809_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__a31oi_4
XPHY_EDGE_ROW_147_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11010_ _03467_ _05213_ _05215_ _03469_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10722__A3 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11338__A _03229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _06296_ VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__buf_2
XANTENNA__12868__S _06928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13553__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14700_ count_cycle\[4\] _08340_ _07826_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__a21oi_1
X_11912_ _06405_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15680_ _04335_ _02479_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__nand2_1
XANTENNA__09971__S1 _04478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12892_ _06948_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_47_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14631_ _08281_ _08282_ _08278_ _08263_ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_157_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11843_ _06367_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10388__S _04320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_156_Left_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ clknet_leaf_185_clk _00519_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_14562_ _08212_ _07954_ VGND VGND VPWR VPWR _08219_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11774_ _06319_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__buf_2
XFILLER_0_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16301_ _06976_ cpuregs.regs\[15\]\[16\] _02870_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13513_ _07274_ _07368_ _07369_ _07190_ VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__a211o_1
X_10725_ _05243_ _05319_ _05423_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__o21a_1
X_17281_ clknet_leaf_186_clk _00455_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_161_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_161_clk sky130_fd_sc_hd__clkbuf_2
X_14493_ _07934_ _07937_ _07939_ _08119_ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__nand4_2
XFILLER_0_165_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16232_ _02840_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__clkbuf_1
X_13444_ _07304_ _04307_ _07305_ reg_pc\[5\] _07283_ VGND VGND VPWR VPWR _07306_ sky130_fd_sc_hd__a221o_1
X_10656_ _03534_ _05357_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output194_A net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16163_ net275 net237 _02797_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__mux2_1
X_10587_ net71 net72 net73 _04708_ _05229_ _05239_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__mux4_1
X_13375_ _03276_ _07230_ _07231_ _07240_ VGND VGND VPWR VPWR _07241_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12108__S _06507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09800__A1 _04272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16803__S _03138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15114_ _01968_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__buf_8
X_12326_ cpuregs.regs\[26\]\[1\] _06536_ _06641_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__mux2_1
XANTENNA__15334__C1 _02006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16094_ _02608_ _02755_ _05973_ _03845_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__a211o_1
XANTENNA__11947__S _06424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15045_ _03272_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__buf_4
XANTENNA__12699__A0 _06216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10851__S _05264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12257_ cpuregs.regs\[25\]\[1\] _06536_ _06604_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output71_A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11208_ reg_next_pc\[7\] reg_out\[7\] _05834_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_112_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12188_ _06558_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__clkbuf_1
X_11139_ _04040_ _04037_ _05808_ _04811_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__a211o_2
X_16996_ clknet_leaf_158_clk _00170_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_15947_ _04016_ _02650_ _02667_ _02669_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__a22o_1
XANTENNA__12778__S _06880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09867__B2 _04053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10477__A2 _04104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15878_ _02631_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14278__B _07944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14829_ _01773_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__clkbuf_1
X_17617_ clknet_leaf_136_clk _00786_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_18597_ clknet_leaf_146_clk _01662_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10229__A2 _04308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17548_ clknet_leaf_158_clk _00717_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17479_ clknet_leaf_178_clk _00648_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_152_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_152_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_982 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09478__S0 _04207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_667 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16117__A1 _03218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10937__B1 _05215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10401__A2 _05107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15837__B _03916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14741__B _08350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14679__A1 _03294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11857__S _06370_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_895 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16014__A mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13351__A1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09804_ count_instr\[43\] instr_rdinstrh instr_rdcycleh count_cycle\[43\] VGND VGND
+ VPWR VPWR _04529_ sky130_fd_sc_hd__a22o_1
XANTENNA__10260__S1 _04218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09735_ reg_pc\[10\] decoded_imm\[10\] VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09402__S0 _04071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11592__S _06086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11665__A1 _06186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09666_ _04392_ _04393_ _04356_ _04359_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__a211o_1
XFILLER_0_96_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08467__A _03240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08617_ irq_mask\[2\] irq_active _03241_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__o21a_1
X_09597_ _04324_ _04326_ _04223_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08548_ irq_mask\[4\] irq_pending\[4\] VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__and2b_4
XFILLER_0_9_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08479_ instr_bltu instr_bge instr_blt instr_bne VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__or4_1
XFILLER_0_119_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_143_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_143_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_42_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14521__B1_N _08012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11621__A _06183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13312__S _07176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10510_ instr_xor instr_xori VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11490_ _06064_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15564__C1 _02027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10441_ reg_pc\[30\] decoded_imm\[30\] VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08572__A_N irq_mask\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16623__S _03040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08597__A1 _03303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10372_ reg_pc\[27\] decoded_imm\[27\] VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13160_ _07103_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14651__B _07967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12111_ _06511_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__clkbuf_1
X_13091_ _06982_ cpuregs.regs\[7\]\[19\] _07057_ VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__mux2_1
X_12042_ _06201_ cpuregs.regs\[22\]\[13\] _06471_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__mux2_1
XANTENNA__09237__S _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16850_ _06565_ cpuregs.regs\[14\]\[15\] _03163_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10251__S1 _04219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15801_ _02584_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09761__A _04055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16781_ _03132_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09849__A1 _04018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13993_ _07761_ _07762_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__nor2_1
X_18520_ clknet_leaf_8_clk _01585_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_15732_ _04806_ _02506_ _02536_ _02481_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__o211a_1
XANTENNA__11656__A1 _06186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12853__A0 _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10003__S1 _04060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12944_ _06983_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10700__A _05244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16044__B1 mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18451_ clknet_leaf_155_clk _01516_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15663_ _04101_ _02477_ _02483_ _02485_ _07775_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__a221oi_1
X_12875_ _06937_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_130 net230 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output207_A net207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17402_ clknet_leaf_111_clk _00571_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12605__A0 _06114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14614_ _08225_ _08265_ _08266_ _08242_ VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__o211a_1
X_11826_ _06358_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__clkbuf_1
X_18382_ clknet_leaf_111_clk _01447_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08659__C_N _03425_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15594_ _02423_ _02424_ _02110_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17333_ clknet_leaf_115_clk _00507_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14545_ _07943_ _07946_ _08162_ _07998_ VGND VGND VPWR VPWR _08204_ sky130_fd_sc_hd__a31o_1
XFILLER_0_139_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_134_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_134_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11757_ _06304_ cpuregs.regs\[10\]\[26\] _06258_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15003__A _04561_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10708_ _05255_ _05261_ _05394_ _05407_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__a31o_1
X_17264_ clknet_leaf_110_clk _00438_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14476_ decoded_imm_j\[14\] _07937_ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__nor2_1
X_11688_ reg_pc\[19\] _06234_ _06101_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09001__A _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16215_ net40 mem_16bit_buffer\[0\] _02831_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13427_ _07287_ _07288_ _07289_ VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_114_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10639_ _03534_ _05340_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17195_ clknet_leaf_150_clk _00369_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16533__S _02990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16146_ net266 net228 _02786_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__mux2_1
X_13358_ _07224_ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15858__B1 _02617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12309_ cpuregs.regs\[25\]\[26\] _06588_ _06626_ VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__mux2_1
X_16077_ decoded_imm\[27\] _02750_ _02746_ mem_rdata_q\[27\] _02749_ VGND VGND VPWR
+ VPWR _01340_ sky130_fd_sc_hd__a221o_1
X_13289_ _06976_ cpuregs.regs\[5\]\[16\] _07165_ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__mux2_1
XANTENNA__10490__S1 _04218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15028_ irq_mask\[23\] _01865_ _01896_ _01891_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_110_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10147__A1 _04215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15181__S1 _01986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 irq[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
X_16979_ clknet_leaf_166_clk _00153_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09520_ net36 net53 _04039_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__mux2_1
XANTENNA__11647__A1 _06186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12301__S _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09451_ _04069_ _04179_ _04183_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__a21oi_1
X_18649_ clknet_leaf_117_clk _01709_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16708__S _03087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08402_ latched_branch latched_store VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10870__A2 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09382_ _04113_ _04114_ _04045_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__a21bo_1
XANTENNA__15794__C1 _06026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09068__A2 _03730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13640__B decoded_imm\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_125_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_125_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__08815__A2 _03460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13132__S _07082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12971__S _06985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16510__A1 _06571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16274__A0 _06949_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09718_ _04214_ _04444_ _04081_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__a21o_1
XANTENNA__12211__S _06555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09926__S1 _04478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10990_ _05425_ _05597_ _05672_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09700__B1 _04427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09649_ cpuregs.regs\[16\]\[7\] cpuregs.regs\[17\]\[7\] cpuregs.regs\[18\]\[7\] cpuregs.regs\[19\]\[7\]
+ _04216_ _04376_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12660_ _06820_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09520__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11611_ _06174_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__buf_2
XFILLER_0_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13260__A0 _06947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08806__A2 _03475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_116_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_116_clk sky130_fd_sc_hd__clkbuf_2
X_12591_ cpuregs.regs\[2\]\[29\] _06594_ _06774_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__mux2_1
XANTENNA__13042__S _07032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14330_ _08004_ _08005_ _07988_ VGND VGND VPWR VPWR _08006_ sky130_fd_sc_hd__o21ai_1
X_11542_ _06108_ _06109_ _06112_ _06093_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__o22a_2
XFILLER_0_151_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15758__A _05037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14261_ reg_pc\[19\] _07926_ _07950_ _07935_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11473_ irq_mask\[24\] _03428_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__or2_1
XANTENNA__16353__S _02896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16000_ cpuregs.raddr1\[0\] _03636_ _06005_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__o21a_1
XFILLER_0_162_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09767__B1 _04100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13212_ _07131_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10424_ cpuregs.regs\[12\]\[29\] cpuregs.regs\[13\]\[29\] cpuregs.regs\[14\]\[29\]
+ cpuregs.regs\[15\]\[29\] _04057_ _04060_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_59_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14192_ latched_branch irq_state\[0\] VGND VGND VPWR VPWR _07900_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09231__A2 _03864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09862__S0 _04273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13143_ _06966_ cpuregs.regs\[4\]\[11\] _07093_ VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__mux2_1
XANTENNA__12182__A _06174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10355_ cpuregs.regs\[12\]\[27\] cpuregs.regs\[13\]\[27\] cpuregs.regs\[14\]\[27\]
+ cpuregs.regs\[15\]\[27\] _04057_ _04060_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08990__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17951_ clknet_leaf_70_clk _08393_ VGND VGND VPWR VPWR reg_out\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11326__A0 _05086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13074_ _07058_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__clkbuf_1
X_10286_ cpuregs.regs\[28\]\[25\] cpuregs.regs\[29\]\[25\] cpuregs.regs\[30\]\[25\]
+ cpuregs.regs\[31\]\[25\] _04291_ _04292_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_72_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12025_ _06132_ cpuregs.regs\[22\]\[5\] _06460_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__mux2_1
X_16902_ clknet_leaf_33_clk _00047_ VGND VGND VPWR VPWR mem_rdata_q\[21\] sky130_fd_sc_hd__dfxtp_2
X_17882_ clknet_leaf_89_clk _01051_ VGND VGND VPWR VPWR count_cycle\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09491__A _04222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13725__B decoded_imm\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16833_ _06548_ cpuregs.regs\[14\]\[7\] _03152_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08819__B net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13217__S _07129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11526__A _06065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16764_ _03123_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12826__A0 _06132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13976_ _03328_ _07677_ _07681_ net154 VGND VGND VPWR VPWR _07750_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15715_ timer\[15\] _02521_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__or2_1
X_18503_ clknet_leaf_154_clk _01568_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11245__B _05877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12927_ _06207_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__buf_2
XANTENNA__10301__A1 _04010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16695_ _06961_ cpuregs.regs\[19\]\[9\] _03076_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15646_ _03199_ _02465_ _02471_ _02472_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__o211a_1
X_18434_ clknet_leaf_137_clk _01499_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__14579__B1 _07904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12858_ _06257_ cpuregs.regs\[6\]\[20\] _06928_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11491__B_N latched_store VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13460__B _04335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18365_ clknet_leaf_185_clk _01430_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11809_ _06096_ cpuregs.regs\[11\]\[1\] _06348_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15577_ cpuregs.regs\[24\]\[28\] cpuregs.regs\[25\]\[28\] cpuregs.regs\[26\]\[28\]
+ cpuregs.regs\[27\]\[28\] _01996_ _01997_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_107_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_107_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_113_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15791__A2 instr_jalr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12789_ cpuregs.regs\[9\]\[20\] _06575_ _06891_ VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__mux2_1
XANTENNA__08554__B irq_pending\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11261__A _04708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17316_ clknet_leaf_159_clk _00490_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15528__C1 _02006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14528_ decoded_imm_j\[18\] _07942_ _07946_ VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__nand3_1
X_18296_ clknet_leaf_5_clk _01364_ VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09470__A2 _04198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17247_ clknet_leaf_181_clk _00421_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14459_ _08106_ _08113_ _08114_ VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__or3_1
XFILLER_0_98_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12791__S _06891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14572__A _07954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17178_ clknet_leaf_188_clk _00352_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10368__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16129_ net289 _05255_ _02771_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08951_ _03711_ _03712_ _03713_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11317__A0 reg_next_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10215__S1 _04473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08882_ _03646_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__buf_8
XANTENNA__15834__C _03920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_4_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16011__B is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08729__B net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12031__S _06460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10340__A reg_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09503_ cpuregs.regs\[8\]\[4\] cpuregs.regs\[9\]\[4\] cpuregs.regs\[10\]\[4\] cpuregs.regs\[11\]\[4\]
+ _04232_ _04233_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__mux4_1
XANTENNA__11096__A2 _05086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13490__B1 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16438__S _02943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14747__A _03239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09434_ _04018_ count_cycle\[35\] _04165_ count_cycle\[3\] _04166_ VGND VGND VPWR
+ VPWR _04167_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15767__C1 _02488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08745__A net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10994__B _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09365_ net300 VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_111_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09296_ _04032_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__buf_4
XANTENNA_30 _04637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 _05923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10151__S0 _04579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08895__S1 _03659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 decoded_imm\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_63 net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15578__A _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_85 net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_96 _02349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_985 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09576__A _04227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10359__A1 _04215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16607__C_N cpuregs.waddr\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10515__A _05218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10140_ cpuregs.regs\[8\]\[21\] cpuregs.regs\[9\]\[21\] cpuregs.regs\[10\]\[21\]
+ cpuregs.regs\[11\]\[21\] _04282_ _04285_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_120_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput170 net170 VGND VGND VPWR VPWR mem_addr[17] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput181 net181 VGND VGND VPWR VPWR mem_addr[28] sky130_fd_sc_hd__clkbuf_1
Xoutput192 net192 VGND VGND VPWR VPWR mem_addr[9] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_54_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10071_ _04018_ count_cycle\[51\] _04013_ count_cycle\[19\] _04787_ VGND VGND VPWR
+ VPWR _04788_ sky130_fd_sc_hd__a221o_1
X_13830_ _07654_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15470__A1 _02066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11087__A2 _05404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13761_ _03631_ _07599_ _07600_ _07225_ VGND VGND VPWR VPWR _07601_ sky130_fd_sc_hd__o31ai_1
X_10973_ _03464_ _05367_ _05656_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12876__S _06928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11780__S _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15500_ _01982_ _02333_ _02335_ _02018_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__o211a_1
X_12712_ _06266_ cpuregs.regs\[12\]\[21\] _06847_ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__mux2_1
XANTENNA__10834__A2 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16480_ _02972_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__clkbuf_1
X_13692_ _07536_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10390__S0 _04290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15431_ cpuregs.regs\[8\]\[20\] cpuregs.regs\[9\]\[20\] cpuregs.regs\[10\]\[20\]
+ cpuregs.regs\[11\]\[20\] _02030_ _02031_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__mux4_1
X_12643_ _06266_ cpuregs.regs\[30\]\[21\] _06810_ VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__mux2_1
XANTENNA__14430__C1 _08097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18150_ clknet_leaf_46_clk alu_out\[24\] VGND VGND VPWR VPWR alu_out_q\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15362_ _03683_ _02205_ _02018_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ _06775_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11795__B1 _06101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08886__S1 _03643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17101_ clknet_leaf_120_clk _00275_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14313_ compressed_instr _07988_ _07989_ _06860_ VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__a211o_1
X_18081_ clknet_leaf_40_clk _01186_ VGND VGND VPWR VPWR mem_do_rinst sky130_fd_sc_hd__dfxtp_1
X_11525_ _06097_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__clkbuf_1
X_15293_ _01984_ _02140_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__or2_1
XANTENNA__12905__A _06149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17032_ clknet_leaf_142_clk _00206_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_14244_ _05857_ _06213_ VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__or2_1
XANTENNA__09486__A _04124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11456_ _06041_ irq_pending\[16\] _06046_ net8 VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10407_ reg_pc\[29\] decoded_imm\[29\] VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11011__A2 _05440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14175_ _07887_ _07888_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__nor2_1
XANTENNA__12116__S _06507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16811__S _03138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11387_ _03228_ _03979_ _03814_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13126_ _06949_ cpuregs.regs\[4\]\[3\] _07082_ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__mux2_1
X_10338_ _04391_ _05020_ _05047_ VGND VGND VPWR VPWR _08387_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15384__S1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11955__S _06424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17934_ clknet_leaf_69_clk _08374_ VGND VGND VPWR VPWR reg_out\[14\] sky130_fd_sc_hd__dfxtp_1
X_13057_ _07049_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__clkbuf_1
X_10269_ instr_retirq _04979_ _04980_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__a21o_1
XANTENNA__09912__B1 instr_rdinstr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12008_ _06456_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13455__B _05209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17865_ clknet_leaf_93_clk _01034_ VGND VGND VPWR VPWR count_cycle\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16816_ _03150_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__clkbuf_1
X_17796_ clknet_leaf_57_clk _00965_ VGND VGND VPWR VPWR reg_pc\[4\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__15461__A1 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13959_ _07737_ _07738_ VGND VGND VPWR VPWR _07739_ sky130_fd_sc_hd__and2_1
X_16747_ _03316_ _03112_ _03113_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__or3_1
XANTENNA__12786__S _06880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09140__A1 _03891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13471__A _04342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16678_ _03077_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18417_ clknet_leaf_117_clk _01482_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15629_ _01959_ _02449_ _02457_ _01932_ decoded_imm\[31\] VGND VGND VPWR VPWR _02458_
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_29_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10038__B1 _04105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13775__A1 _05227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09150_ _03861_ _03901_ _03905_ _03888_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18348_ clknet_leaf_30_clk _01416_ VGND VGND VPWR VPWR mem_rdata_q\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11250__A2 _05877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09081_ _03841_ _03237_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18279_ clknet_leaf_31_clk _01349_ VGND VGND VPWR VPWR is_sb_sh_sw sky130_fd_sc_hd__dfxtp_4
XFILLER_0_140_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13527__A1 _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput50 mem_rdata[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_2
XFILLER_0_13_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput61 mem_rdata[6] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_1
XANTENNA__11538__B1 _03344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09826__S0 _04216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16721__S _03098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10210__B1 _04013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09983_ _04051_ _04702_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_164_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15375__S1 _01909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11865__S _06370_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08934_ cpuregs.regs\[20\]\[3\] cpuregs.regs\[21\]\[3\] cpuregs.regs\[22\]\[3\] cpuregs.regs\[23\]\[3\]
+ _03658_ _03659_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__mux4_1
XANTENNA__16229__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16022__A _02611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08865_ _03311_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08459__B net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15861__A _03940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08796_ _03493_ _03560_ _03561_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_142_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11069__A2 _05013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13463__A0 _04342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09131__B2 _03888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15204__A1 _03654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16401__A0 _07007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09417_ _04143_ _04144_ _04148_ _04150_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15755__A2 _02486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10029__B1 _04747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09348_ _04070_ _04079_ _04082_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10944__S _05390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09279_ _04015_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__buf_4
XANTENNA__10675__S1 _05239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13320__S _07153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11310_ _05931_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_132_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12290_ cpuregs.regs\[25\]\[17\] _06569_ _06615_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09198__A1 _03730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11241_ _05875_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_4
XFILLER_0_121_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10427__S1 _04469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10201__B1 _04673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12741__A2 _06863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11172_ _04038_ _05254_ net102 _03297_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__a22o_1
XANTENNA__11775__S _06258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10123_ _04837_ _04838_ _04287_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__mux2_1
X_15980_ _03891_ _03767_ _02600_ _03862_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__a31o_1
X_10054_ cpuregs.regs\[12\]\[18\] cpuregs.regs\[13\]\[18\] cpuregs.regs\[14\]\[18\]
+ cpuregs.regs\[15\]\[18\] _04232_ _04233_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__mux4_1
X_14931_ _01840_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__clkbuf_1
X_17650_ clknet_leaf_47_clk _00819_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dfxtp_2
X_14862_ count_cycle\[55\] count_cycle\[56\] _01792_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15443__A1 _02020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16601_ _07003_ cpuregs.regs\[18\]\[29\] _03026_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__mux2_1
X_13813_ cpuregs.regs\[0\]\[3\] VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12257__A1 _06536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17581_ clknet_leaf_149_clk _00750_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14793_ count_cycle\[33\] _01745_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16532_ _02999_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13744_ _05174_ _04913_ _07276_ VGND VGND VPWR VPWR _07585_ sky130_fd_sc_hd__mux2_1
X_10956_ _03482_ _05627_ _03569_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_161_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16463_ _07001_ cpuregs.regs\[29\]\[28\] _02954_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__mux2_1
X_13675_ _07304_ _04871_ _07305_ reg_pc\[21\] _07283_ VGND VGND VPWR VPWR _07521_
+ sky130_fd_sc_hd__a221o_1
X_10887_ _03493_ _05357_ _05478_ _05575_ _05576_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_14_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18202_ clknet_leaf_43_clk _01273_ VGND VGND VPWR VPWR instr_andi sky130_fd_sc_hd__dfxtp_1
X_15414_ cpuregs.regs\[12\]\[19\] cpuregs.regs\[13\]\[19\] cpuregs.regs\[14\]\[19\]
+ cpuregs.regs\[15\]\[19\] _01936_ _03647_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_100_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12626_ _06201_ cpuregs.regs\[30\]\[13\] _06799_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16394_ _02926_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10115__S0 _04275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18133_ clknet_leaf_40_clk alu_out\[7\] VGND VGND VPWR VPWR alu_out_q\[7\] sky130_fd_sc_hd__dfxtp_1
X_15345_ cpuregs.regs\[20\]\[15\] cpuregs.regs\[21\]\[15\] cpuregs.regs\[22\]\[15\]
+ cpuregs.regs\[23\]\[15\] _02069_ _02070_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12557_ _06766_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15649__C _04006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15054__S0 _03658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13230__S _07140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18064_ clknet_leaf_73_clk _01169_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dfxtp_4
X_11508_ cpuregs.waddr\[3\] VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15276_ cpuregs.regs\[16\]\[11\] cpuregs.regs\[17\]\[11\] cpuregs.regs\[18\]\[11\]
+ cpuregs.regs\[19\]\[11\] _01985_ _01986_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__mux4_1
X_12488_ _06729_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10991__A1 _05219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17015_ clknet_leaf_177_clk _00189_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14227_ _07905_ VGND VGND VPWR VPWR _07926_ sky130_fd_sc_hd__clkbuf_4
X_11439_ irq_mask\[9\] _06030_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16541__S _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14158_ _06053_ VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10743__A1 _03524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11940__A0 _06336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11685__S _06176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13466__A _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13109_ _07076_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__clkbuf_1
X_14089_ count_instr\[33\] count_instr\[32\] _07824_ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17917_ clknet_leaf_82_clk _01086_ VGND VGND VPWR VPWR count_cycle\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09361__A1 _04053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08650_ timer\[25\] timer\[24\] timer\[27\] timer\[26\] VGND VGND VPWR VPWR _03417_
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_124_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17848_ clknet_leaf_64_clk _01017_ VGND VGND VPWR VPWR reg_next_pc\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12248__A1 _06598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08581_ _03356_ _03357_ _03358_ _03359_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__or4_1
X_17779_ clknet_leaf_86_clk _00948_ VGND VGND VPWR VPWR count_instr\[50\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__14297__A irq_pending\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16716__S _03087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09202_ _03767_ _03947_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__nor2_1
XANTENNA__14945__A0 net207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09133_ mem_rdata_q\[23\] _03889_ _03846_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10431__B1 _04100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09064_ mem_16bit_buffer\[9\] _03825_ _03727_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__mux2_4
XANTENNA__10982__A1 _05517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15856__A _03239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16451__S _02954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09854__A _04483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15348__S1 _02075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09966_ cpuregs.regs\[28\]\[16\] cpuregs.regs\[29\]\[16\] cpuregs.regs\[30\]\[16\]
+ cpuregs.regs\[31\]\[16\] _04579_ _04470_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__mux4_1
X_08917_ _03638_ _03313_ _03315_ _03681_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__a31o_1
X_09897_ cpuregs.regs\[8\]\[14\] cpuregs.regs\[9\]\[14\] cpuregs.regs\[10\]\[14\]
+ cpuregs.regs\[11\]\[14\] _04216_ _04376_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_96_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_2
X_08848_ net128 _03518_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__and2_1
XANTENNA__10004__S _04065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15425__A1 _03654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08779_ net126 _03524_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__or2b_1
XANTENNA__15520__S1 _03639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10810_ _05499_ _05503_ _05363_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _06072_ _03328_ _06098_ _06333_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09655__A2 _04308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10345__S0 _04758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10741_ _05436_ _05438_ _05278_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10670__A0 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14936__A0 net203 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13460_ _03387_ _04335_ VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10672_ _04198_ _04262_ _04251_ _04342_ _05235_ _05324_ VGND VGND VPWR VPWR _05373_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12411_ cpuregs.regs\[27\]\[9\] _06552_ _06678_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11214__A2 _05848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10648__S1 _05237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13391_ _07232_ _07251_ _07253_ _07255_ VGND VGND VPWR VPWR _07256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_23_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15130_ _01936_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__buf_8
XANTENNA__10422__B1 _04082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12342_ cpuregs.regs\[26\]\[9\] _06552_ _06641_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__mux2_1
XANTENNA__15587__S1 _03684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15061_ cpuregs.regs\[24\]\[0\] cpuregs.regs\[25\]\[0\] cpuregs.regs\[26\]\[0\] cpuregs.regs\[27\]\[0\]
+ _03670_ _03671_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__mux4_1
X_12273_ cpuregs.regs\[25\]\[9\] _06552_ _06604_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14012_ _03239_ VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_12_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11224_ _05852_ _05860_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__and2_2
XANTENNA__09040__A0 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15339__S1 _02031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11922__A0 _06266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11155_ _05812_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__buf_2
XFILLER_0_156_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16861__A0 _06575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10106_ reg_pc\[20\] decoded_imm\[20\] VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__or2_1
X_11086_ _03442_ _05761_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__xnor2_1
X_15963_ net65 _02673_ _02683_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__o21ai_1
XANTENNA_output237_A net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13675__B1 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_87_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_171_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17702_ clknet_leaf_75_clk _00871_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dfxtp_1
X_10037_ _04046_ _04754_ _04202_ irq_pending\[18\] VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__a22o_1
X_14914_ _01831_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11237__C _05868_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15894_ instr_sh _02635_ _02637_ is_sb_sh_sw VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11150__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15932__C mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ clknet_leaf_50_clk _00802_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_19_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14845_ count_cycle\[49\] _01780_ count_cycle\[50\] VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08827__B net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13225__S _07129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14776_ _01736_ _01737_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__nor2_1
X_17564_ clknet_leaf_105_clk _00733_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11988_ _06423_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__buf_6
XANTENNA__11989__A0 _06257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13727_ _07567_ _07568_ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_82_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16515_ cpuregs.regs\[17\]\[20\] _06575_ _02990_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__mux2_1
X_10939_ _05281_ _05618_ _05619_ _05625_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__a211o_1
XFILLER_0_156_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17495_ clknet_leaf_119_clk _00664_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15275__S0 _01982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13658_ _07472_ _07489_ VGND VGND VPWR VPWR _07505_ sky130_fd_sc_hd__or2b_1
XANTENNA__09939__A _04051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16446_ _02931_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__buf_6
XANTENNA__08843__A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12609_ _06132_ cpuregs.regs\[30\]\[5\] _06788_ VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__mux2_1
X_16377_ _02917_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13589_ _04659_ VGND VGND VPWR VPWR _07441_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12365__A _06640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_81_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18116_ clknet_leaf_82_clk _01220_ VGND VGND VPWR VPWR timer\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10413__B1 _04145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15328_ _02066_ _02173_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10964__B2 _05251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18047_ clknet_leaf_77_clk _00025_ VGND VGND VPWR VPWR irq_pending\[31\] sky130_fd_sc_hd__dfxtp_1
X_15259_ _02066_ _02108_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__or2_1
XANTENNA__14580__A _07954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09820_ count_instr\[44\] _04016_ count_cycle\[12\] _04013_ _04543_ VGND VGND VPWR
+ VPWR _04544_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09751_ _04084_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_78_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_2
X_08702_ net114 net82 VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__nand2_1
XANTENNA__13924__A _06053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09682_ cpuregs.regs\[16\]\[8\] cpuregs.regs\[17\]\[8\] cpuregs.regs\[18\]\[8\] cpuregs.regs\[19\]\[8\]
+ _04056_ _04091_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__mux4_1
XANTENNA__11141__A1 _03407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11141__B2 _04422_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10575__S0 _05277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15407__A1 _02004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09613__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08633_ _03404_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15502__S1 _02023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08737__B net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16080__A1 decoded_imm\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16080__B2 mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08564_ irq_mask\[23\] irq_pending\[23\] VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__and2b_1
XFILLER_0_119_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08495_ mem_do_prefetch _03237_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__and2_1
XANTENNA__12974__S _06985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14755__A _06053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08753__A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12275__A _06603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08472__B instr_jalr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09496__S1 _04208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09116_ mem_rdata_q\[21\] _03874_ _03846_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15569__S1 _01974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09047_ mem_16bit_buffer\[3\] _03728_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__nor2_1
XANTENNA__16181__S _02770_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_746 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15894__B2 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10523__A _05209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15646__A1 _03199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09949_ net39 _04034_ _04669_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_69_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _06994_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11132__A1 _05413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08928__A _00068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11911_ _06224_ cpuregs.regs\[20\]\[16\] _06398_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__mux2_1
XANTENNA__13553__B decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11683__A2 reg_next_pc\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12891_ _06947_ cpuregs.regs\[31\]\[2\] _06943_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11354__A _03215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14630_ _08269_ _08272_ _08280_ _08097_ VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__a31o_1
X_11842_ _06232_ cpuregs.regs\[11\]\[17\] _06359_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _03294_ _07954_ _07997_ _08217_ VGND VGND VPWR VPWR _08218_ sky130_fd_sc_hd__a22o_1
X_11773_ _06116_ reg_next_pc\[28\] _06316_ _06318_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__a211o_2
XFILLER_0_68_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13512_ _04456_ _05259_ _07332_ _07254_ VGND VGND VPWR VPWR _07369_ sky130_fd_sc_hd__o211a_1
XANTENNA__14909__A0 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16300_ _02876_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__clkbuf_1
X_10724_ _05242_ _05316_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__nand2_1
X_17280_ clknet_leaf_13_clk _00454_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08931__S0 _03641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14492_ _07934_ _07937_ _08119_ _07939_ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16231_ net49 mem_16bit_buffer\[8\] _02831_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13443_ _07211_ VGND VGND VPWR VPWR _07305_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15582__B1 _02412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10655_ _05356_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_152_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16162_ _02799_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__clkbuf_1
X_13374_ _07232_ _07233_ _07235_ _07239_ VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__a22o_1
X_10586_ net98 net68 net69 net70 _05229_ _05239_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15113_ _03654_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__buf_8
XFILLER_0_51_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12325_ _06642_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__clkbuf_1
X_16093_ is_sb_sh_sw _03636_ _02757_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14688__A2 _07948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15044_ irq_mask\[31\] _01865_ _01904_ _01891_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__a211o_1
X_12256_ _06605_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10159__C1 _04150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11207_ _05847_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__buf_4
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12187_ cpuregs.regs\[24\]\[11\] _06557_ _06555_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__mux2_1
XANTENNA__15098__C1 _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15637__A1 _03298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11138_ _04040_ _04033_ _05808_ _04811_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__a211o_2
X_16995_ clknet_leaf_131_clk _00169_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11963__S _06424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11069_ _05076_ _05044_ _05013_ _04959_ _05237_ _05266_ VGND VGND VPWR VPWR _05746_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__15865__C_N _03940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15946_ _04012_ _02650_ _02659_ _02669_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_0_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_2
X_15877_ instr_jalr _02630_ _03635_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__mux2_1
XANTENNA__08557__B irq_pending\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17616_ clknet_leaf_130_clk _00785_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_14828_ _01771_ _01753_ _01772_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__and3b_1
XFILLER_0_59_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18596_ clknet_leaf_138_clk _01661_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17547_ clknet_leaf_127_clk _00716_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14759_ count_cycle\[22\] _01722_ _01725_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08922__S0 _03641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17478_ clknet_leaf_17_clk _00647_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16429_ _02945_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09478__S1 _04208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16117__A2 _03199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12139__A0 _06312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14679__A2 _07971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15420__S0 _03645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15628__A1 _02017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16825__A0 _06540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09803_ instr_retirq _04526_ _04527_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09307__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09307__B2 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09734_ irq_pending\[9\] _04008_ _04451_ _04460_ VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_2_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08748__A net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09402__S1 _04073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09665_ reg_pc\[8\] decoded_imm\[8\] VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__or2_1
XANTENNA__11665__A2 reg_next_pc\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10489__S _04223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15487__S0 _03645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16053__A1 decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08616_ _03386_ _03390_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__or2_1
X_09596_ cpuregs.regs\[0\]\[6\] cpuregs.regs\[1\]\[6\] cpuregs.regs\[2\]\[6\] cpuregs.regs\[3\]\[6\]
+ _04325_ _04277_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__mux4_1
XFILLER_0_139_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08547_ irq_mask\[2\] irq_pending\[2\] VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__and2b_2
XFILLER_0_49_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14485__A decoded_imm_j\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15239__S0 _01985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08478_ instr_or instr_sra instr_srl instr_xor VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10440_ reg_pc\[30\] decoded_imm\[30\] VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09243__B1 _03867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10928__A1 _05517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08597__A2 _03254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10371_ _04391_ _05052_ _05079_ VGND VGND VPWR VPWR _08388_ sky130_fd_sc_hd__a21o_1
XANTENNA__13590__A2 _07441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15411__S0 _03670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12110_ _06201_ cpuregs.regs\[23\]\[13\] _06507_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__mux2_1
X_13090_ _07066_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12041_ _06474_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10253__A _04369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15800_ _08033_ _07994_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__and2_1
X_16780_ _06563_ cpuregs.regs\[13\]\[14\] _03127_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__mux2_1
X_13992_ count_instr\[2\] _07758_ _07759_ VGND VGND VPWR VPWR _07762_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_184_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15731_ timer\[19\] _02533_ _02535_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__o21ai_1
X_12943_ _06982_ cpuregs.regs\[31\]\[19\] _06964_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__mux2_1
XANTENNA__11656__A2 reg_next_pc\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16044__A1 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15478__S0 _01995_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18450_ clknet_leaf_125_clk _01515_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_15662_ _02482_ _02478_ _02484_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__o21a_1
XANTENNA_120 net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12874_ _06320_ cpuregs.regs\[6\]\[28\] _06928_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__mux2_1
XANTENNA_131 _01753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17401_ clknet_leaf_161_clk _00570_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_153 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11825_ _06166_ cpuregs.regs\[11\]\[9\] _06348_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__mux2_1
X_14613_ _07958_ _07959_ _08221_ VGND VGND VPWR VPWR _08266_ sky130_fd_sc_hd__o21ai_1
XANTENNA_output102_A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15593_ cpuregs.regs\[24\]\[29\] cpuregs.regs\[25\]\[29\] cpuregs.regs\[26\]\[29\]
+ cpuregs.regs\[27\]\[29\] _02221_ _02222_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__mux4_1
X_18381_ clknet_leaf_164_clk _01446_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12908__A _06156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17332_ clknet_leaf_112_clk _00506_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_14544_ _08201_ _08202_ _07972_ VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_138_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11756_ _06303_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__buf_2
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10092__A1 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10707_ _05298_ _05396_ _05406_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__a21bo_1
XANTENNA__14358__A1 _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17263_ clknet_leaf_122_clk _00437_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_14475_ decoded_imm_j\[14\] _07937_ VGND VGND VPWR VPWR _08139_ sky130_fd_sc_hd__and2_1
X_11687_ reg_pc\[19\] _06234_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13426_ _07260_ _07261_ _07259_ VGND VGND VPWR VPWR _07289_ sky130_fd_sc_hd__a21bo_1
X_16214_ _02830_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__clkbuf_4
X_10638_ _03538_ _05339_ _05323_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__mux2_1
X_17194_ clknet_leaf_147_clk _00368_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13030__A1 _06580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10919__A1 _05281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16145_ _02790_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__clkbuf_1
X_13357_ _07223_ VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10569_ _05271_ _05272_ _05240_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08840__B net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15858__A1 _03309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15858__B2 instr_beq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12308_ _06632_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16076_ decoded_imm\[26\] _02750_ _02746_ mem_rdata_q\[26\] _02749_ VGND VGND VPWR
+ VPWR _01339_ sky130_fd_sc_hd__a221o_1
X_13288_ _07171_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_137_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15027_ _04940_ _01885_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__nor2_1
XANTENNA__15954__A _03196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12239_ cpuregs.regs\[24\]\[28\] _06592_ _06576_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16807__A0 _06590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09952__A cpu_state\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12789__S _06891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14294__B1 _07971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16978_ clknet_leaf_111_clk _00152_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 irq[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
X_15929_ instr_and _02617_ _02627_ _02653_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__a22o_1
XANTENNA__11647__A2 reg_next_pc\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10304__C1 _04202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16035__A1 decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15469__S0 _02069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09450_ _04052_ _04182_ _00073_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__a21o_1
X_18648_ clknet_leaf_113_clk _01708_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08401_ mem_la_secondword VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09381_ _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__inv_2
XANTENNA__14597__B2 _03378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18579_ clknet_leaf_155_clk _01644_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10870__A3 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11722__A _06273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09473__B1 _04165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15546__B1 _03657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_0_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12029__S _06460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13021__A1 _06571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14752__B _08350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10138__A2 _04016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12699__S _06836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14285__B1 _07966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09717_ _04442_ _04443_ _04078_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__mux2_1
XANTENNA__11638__A2 _03352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09700__A1 _04391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10012__S _04121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09648_ cpuregs.regs\[20\]\[7\] cpuregs.regs\[21\]\[7\] cpuregs.regs\[22\]\[7\] cpuregs.regs\[23\]\[7\]
+ _04216_ _04376_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__mux4_1
XANTENNA__14037__B1 _07790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10947__S _05230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09579_ _04271_ _04307_ _04309_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_26_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12599__A0 _06078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11610_ _06170_ _06173_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__nor2_4
XFILLER_0_155_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12590_ _06783_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11541_ _06110_ _06111_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16634__S _03051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14260_ reg_next_pc\[19\] _05876_ _07922_ _07949_ VGND VGND VPWR VPWR _07950_ sky130_fd_sc_hd__o211a_2
XFILLER_0_34_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11472_ _06054_ irq_pending\[23\] _06055_ net16 VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15758__B _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13211_ _06966_ cpuregs.regs\[8\]\[11\] _07129_ VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10423_ cpuregs.regs\[8\]\[29\] cpuregs.regs\[9\]\[29\] cpuregs.regs\[10\]\[29\]
+ cpuregs.regs\[11\]\[29\] _04057_ _04060_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14191_ _07898_ VGND VGND VPWR VPWR _07899_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09862__S1 _04283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13142_ _07094_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09248__S _03757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10354_ _05061_ _05062_ _04211_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17950_ clknet_leaf_70_clk _08392_ VGND VGND VPWR VPWR reg_out\[30\] sky130_fd_sc_hd__dfxtp_1
X_13073_ _06963_ cpuregs.regs\[7\]\[10\] _07057_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10285_ _04287_ _04993_ _04995_ _04289_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__o211a_1
XANTENNA__10129__A2 _04104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13720__C1 _07221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12024_ _06465_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__clkbuf_1
X_16901_ clknet_leaf_33_clk _00046_ VGND VGND VPWR VPWR mem_rdata_q\[20\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_72_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Right_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17881_ clknet_leaf_89_clk _01050_ VGND VGND VPWR VPWR count_cycle\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16832_ _03159_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14276__B1 _07959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11629__A2 _03357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16763_ _06546_ cpuregs.regs\[13\]\[6\] _03116_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__mux2_1
X_13975_ _07749_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16809__S _03138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18502_ clknet_leaf_146_clk _01567_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_15714_ timer\[15\] _02521_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__and2_1
X_12926_ _06971_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__clkbuf_1
X_16694_ _03085_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14837__B _01753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18433_ clknet_leaf_147_clk _01498_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__14579__A1 _07898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15645_ _03239_ _03310_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__nor2_1
XANTENNA__14579__B2 reg_next_pc\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12857_ _06905_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15014__A _04737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18364_ clknet_leaf_174_clk _01429_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11808_ _06349_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__clkbuf_1
X_12788_ _06868_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__clkbuf_8
X_15576_ _02111_ _02407_ _01968_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__o21a_1
X_17315_ clknet_leaf_131_clk _00489_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11739_ _06288_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__buf_2
X_14527_ _07942_ _07946_ decoded_imm_j\[18\] VGND VGND VPWR VPWR _08187_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18295_ clknet_leaf_5_clk _01363_ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09207__A0 mem_rdata_q\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17246_ clknet_leaf_166_clk _00420_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__14200__A0 reg_next_pc\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08851__A net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14458_ _08071_ _08117_ _08118_ _08123_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__a211o_1
XFILLER_0_154_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14572__B _07988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13409_ _04419_ VGND VGND VPWR VPWR _07272_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17177_ clknet_leaf_14_clk _00351_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_14389_ decoded_imm_j\[7\] _07921_ VGND VGND VPWR VPWR _08060_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16128_ _02781_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08950_ _03652_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16059_ decoded_imm\[17\] _02720_ _02736_ _02742_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08881_ _00065_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10621__A _05230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14267__B1 _07954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16011__C is_alu_reg_imm VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10340__B decoded_imm\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16719__S _03098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09502_ cpuregs.regs\[12\]\[4\] cpuregs.regs\[13\]\[4\] cpuregs.regs\[14\]\[4\] cpuregs.regs\[15\]\[4\]
+ _04232_ _04233_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__mux4_1
XFILLER_0_154_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15623__S _03709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08497__A1 mem_do_wdata VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09433_ count_instr\[35\] _04104_ _04145_ count_instr\[3\] VGND VGND VPWR VPWR _04166_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08745__B _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13143__S _07093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13778__C1 _07221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09364_ cpuregs.raddr1\[3\] cpuregs.raddr1\[2\] cpuregs.raddr1\[4\] _04098_ VGND
+ VGND VPWR VPWR _04099_ sky130_fd_sc_hd__nor4_4
XFILLER_0_136_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11253__A0 reg_next_pc\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09295_ _04030_ _04031_ _03243_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_7_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_20 _03979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _04743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10151__S1 _04284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_42 _06141_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_53 decoded_imm_j\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_64 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08761__A net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_86 net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13379__A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 _03304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08421__A1 net262 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput160 net160 VGND VGND VPWR VPWR eoi[7] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_37_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput171 net171 VGND VGND VPWR VPWR mem_addr[18] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput182 net182 VGND VGND VPWR VPWR mem_addr[29] sky130_fd_sc_hd__buf_1
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10070_ count_instr\[51\] _04104_ _04011_ count_instr\[19\] VGND VGND VPWR VPWR _04787_
+ sky130_fd_sc_hd__a22o_1
Xoutput193 net193 VGND VGND VPWR VPWR mem_instr sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16247__A1 _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13318__S _07153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14258__B1 _07948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13760_ _07578_ _07581_ _07598_ VGND VGND VPWR VPWR _07600_ sky130_fd_sc_hd__a21oi_1
X_10972_ _05220_ _03466_ _03465_ _05440_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13481__A1 _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12711_ _06848_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__clkbuf_1
X_13691_ _04913_ _07535_ _07224_ VGND VGND VPWR VPWR _07536_ sky130_fd_sc_hd__mux2_1
XANTENNA__10834__A3 _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10390__S1 _04283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11362__A _03228_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12642_ _06811_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__clkbuf_1
X_15430_ cpuregs.regs\[12\]\[20\] cpuregs.regs\[13\]\[20\] cpuregs.regs\[14\]\[20\]
+ cpuregs.regs\[15\]\[20\] _01979_ _01980_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15361_ _02203_ _02204_ _01984_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__mux2_1
X_12573_ cpuregs.regs\[2\]\[20\] _06575_ _06774_ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__mux2_1
XANTENNA__16364__S _02907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17100_ clknet_leaf_180_clk _00274_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15605__S0 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11524_ _06096_ cpuregs.regs\[10\]\[1\] _06086_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__mux2_1
X_14312_ _05856_ _06088_ _07901_ _03190_ VGND VGND VPWR VPWR _07989_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_124_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18080_ clknet_leaf_26_clk _01185_ VGND VGND VPWR VPWR mem_do_prefetch sky130_fd_sc_hd__dfxtp_2
X_15292_ cpuregs.regs\[28\]\[12\] cpuregs.regs\[29\]\[12\] cpuregs.regs\[30\]\[12\]
+ cpuregs.regs\[31\]\[12\] _01985_ _01986_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14243_ reg_pc\[14\] _07926_ _07937_ _07935_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__a22o_1
X_17031_ clknet_leaf_147_clk _00205_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_11455_ irq_mask\[16\] _06042_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10406_ reg_pc\[29\] decoded_imm\[29\] VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14174_ count_instr\[58\] _07884_ _07877_ VGND VGND VPWR VPWR _07888_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11386_ _03845_ _03971_ _05991_ _05995_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13125_ _07085_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__clkbuf_1
X_10337_ irq_pending\[26\] _04007_ _05043_ _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12921__A _06192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17933_ clknet_leaf_66_clk _08373_ VGND VGND VPWR VPWR reg_out\[13\] sky130_fd_sc_hd__dfxtp_1
X_13056_ _06947_ cpuregs.regs\[7\]\[2\] _07046_ VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__mux2_1
X_10268_ irq_mask\[24\] _04308_ timer\[24\] instr_timer _04025_ VGND VGND VPWR VPWR
+ _04980_ sky130_fd_sc_hd__a221o_1
X_12007_ _06328_ cpuregs.regs\[21\]\[29\] _06446_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__mux2_1
XANTENNA__11537__A _06098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17864_ clknet_leaf_96_clk _01033_ VGND VGND VPWR VPWR count_cycle\[9\] sky130_fd_sc_hd__dfxtp_1
X_10199_ net81 VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_109_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16815_ _06598_ cpuregs.regs\[13\]\[31\] _03115_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__mux2_1
XANTENNA__09007__A _03767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10160__B decoded_imm\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17795_ clknet_leaf_57_clk _00964_ VGND VGND VPWR VPWR reg_pc\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15944__D_N mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16746_ reg_sh\[0\] _03399_ _04046_ reg_sh\[1\] VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__o211a_1
X_13958_ _03342_ _07727_ _07728_ net147 VGND VGND VPWR VPWR _07738_ sky130_fd_sc_hd__a22o_1
XANTENNA__09676__B1 _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09140__A2 _03892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15749__B1 _02488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13471__B _05259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12909_ _06959_ cpuregs.regs\[31\]\[8\] _06943_ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16677_ _06941_ cpuregs.regs\[19\]\[0\] _03076_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13889_ _07675_ _07689_ VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_122_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18416_ clknet_leaf_108_clk _01481_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15628_ _02017_ _02452_ _02456_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_17_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13775__A2 _05334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18347_ clknet_leaf_35_clk _01415_ VGND VGND VPWR VPWR mem_rdata_q\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16274__S _02859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15559_ _02066_ _02391_ _03692_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__o21a_1
X_09080_ _03229_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__buf_2
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08581__A _03356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18278_ clknet_leaf_29_clk _01348_ VGND VGND VPWR VPWR is_jalr_addi_slti_sltiu_xori_ori_andi
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput40 mem_rdata[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17229_ clknet_leaf_121_clk _00403_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12307__S _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput51 mem_rdata[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
XANTENNA__11538__A1 irq_state\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput62 mem_rdata[7] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_1
XFILLER_0_71_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11538__B2 _06072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09826__S1 _04376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10210__A1 _04105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09982_ _04689_ _04693_ _04100_ _04701_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__a211o_4
XFILLER_0_40_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08933_ _03695_ _03696_ _03687_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13138__S _07082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11447__A _03305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08864_ _03601_ _03603_ _03629_ _03626_ _03623_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__o32a_2
XANTENNA__12042__S _06471_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11710__A1 alu_out_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08795_ net104 net72 VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_142_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16449__S _02954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13662__A _03276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11069__A3 _04959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11474__B1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09762__S0 _04487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09416_ _04149_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11182__A _03219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14412__B1 _07997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10029__A1 _04150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09347_ _04081_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14963__A1 irq_active VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14493__A _07934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09587__A _04283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09278_ instr_rdinstrh VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08491__A cpu_state\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12726__A0 _06320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11240_ _04566_ _05874_ _05827_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09198__A2 _03867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11171_ net118 _04710_ _05820_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__a21o_2
XANTENNA__10201__B2 _04914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10122_ cpuregs.regs\[16\]\[20\] cpuregs.regs\[17\]\[20\] cpuregs.regs\[18\]\[20\]
+ cpuregs.regs\[19\]\[20\] _04282_ _04285_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13151__A0 _06974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13048__S _07009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10053_ _04321_ _04770_ _04069_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__o21a_1
X_14930_ net200 net169 _01835_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__mux2_1
XANTENNA__11701__A1 _06252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14861_ count_cycle\[55\] _01792_ _01794_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__o21a_1
XANTENNA__15979__B1 _02695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14668__A _08232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13572__A _04754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16640__A1 _06215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16600_ _03035_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__clkbuf_1
X_13812_ _07645_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__clkbuf_1
X_17580_ clknet_leaf_115_clk _00749_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08666__A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14792_ count_cycle\[32\] count_cycle\[33\] count_cycle\[31\] _01741_ VGND VGND VPWR
+ VPWR _01748_ sky130_fd_sc_hd__and4_2
XANTENNA__10268__B2 instr_timer VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16531_ cpuregs.regs\[17\]\[28\] _06592_ _02990_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10955_ _03480_ _05629_ _03481_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__a21boi_1
X_13743_ _03583_ _07315_ _07583_ VGND VGND VPWR VPWR _07584_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09753__S0 _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16462_ _02962_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__clkbuf_1
X_10886_ _03492_ _05398_ _05367_ _03491_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__o22a_1
X_13674_ _04913_ _07277_ _07519_ _07238_ VGND VGND VPWR VPWR _07520_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18201_ clknet_leaf_43_clk _01272_ VGND VGND VPWR VPWR instr_ori sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15413_ _02252_ _02253_ _03664_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12625_ _06802_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15499__A _01989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16393_ _06999_ cpuregs.regs\[16\]\[27\] _02918_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10115__S1 _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18132_ clknet_leaf_28_clk alu_out\[6\] VGND VGND VPWR VPWR alu_out_q\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12556_ cpuregs.regs\[2\]\[12\] _06559_ _06763_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__mux2_1
X_15344_ _02066_ _02188_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15054__S1 _03659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11507_ cpuregs.waddr\[4\] VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__clkbuf_4
X_18063_ clknet_leaf_73_clk _01168_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dfxtp_4
XANTENNA__10436__A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12487_ _06193_ cpuregs.regs\[28\]\[12\] _06726_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__mux2_1
X_15275_ _02120_ _02121_ _02122_ _02123_ _01982_ _02088_ VGND VGND VPWR VPWR _02124_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12127__S _06518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17014_ clknet_leaf_126_clk _00188_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_output94_A net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14226_ reg_pc\[9\] _07906_ _07925_ _07912_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__a22o_1
X_11438_ _06029_ irq_pending\[8\] _06036_ net31 VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14157_ count_instr\[53\] _07874_ VGND VGND VPWR VPWR _07876_ sky130_fd_sc_hd__and2_1
X_11369_ _03885_ _05981_ _05979_ _03634_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_146_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13108_ _06999_ cpuregs.regs\[7\]\[27\] _07068_ VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__mux2_1
XANTENNA__13466__B decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14088_ count_instr\[32\] _07824_ _07827_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11267__A _04744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17916_ clknet_leaf_82_clk _01085_ VGND VGND VPWR VPWR count_cycle\[61\] sky130_fd_sc_hd__dfxtp_1
X_13039_ _07039_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13693__A1 _04913_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17847_ clknet_leaf_60_clk _01016_ VGND VGND VPWR VPWR reg_next_pc\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12797__S _06891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08580_ irq_mask\[8\] irq_pending\[8\] VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__and2b_2
X_17778_ clknet_leaf_86_clk _00947_ VGND VGND VPWR VPWR count_instr\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08576__A _03351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11456__B1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16729_ _06995_ cpuregs.regs\[19\]\[25\] _03098_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09201_ _03779_ _03789_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14945__A1 net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12956__A0 _06991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11730__A _06280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09132_ _03850_ _03819_ _03820_ _03849_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__a22o_1
XANTENNA__08624__A1 _03309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09063_ _03823_ _03824_ _03203_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_7_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15856__B _02610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15370__B2 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10065__B decoded_imm\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12184__A1 _06554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10290__S0 _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09965_ _04683_ _04684_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_51_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15872__A _02612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08916_ _03677_ _03679_ _03680_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__a21oi_1
X_09896_ cpuregs.regs\[12\]\[14\] cpuregs.regs\[13\]\[14\] cpuregs.regs\[14\]\[14\]
+ cpuregs.regs\[15\]\[14\] _04216_ _04376_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__mux4_1
XANTENNA__10512__C _05213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10498__A1 _04271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09870__A _04592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10042__S0 _04758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08847_ net128 net96 VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16179__S _02770_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08778_ _03529_ _03542_ _03543_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11116__S _05324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10345__S1 _04759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10740_ _05437_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10670__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10671_ _05371_ _05304_ _05309_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12947__A0 _06984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12410_ _06687_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11640__A _06200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13331__S _04211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13390_ _03312_ _04342_ _05259_ _07254_ VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_62_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_973 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12341_ _06650_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10422__A1 _04070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09110__A _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16642__S _03051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10973__A2 _05367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15060_ cpuregs.regs\[28\]\[0\] cpuregs.regs\[29\]\[0\] cpuregs.regs\[30\]\[0\] cpuregs.regs\[31\]\[0\]
+ _01918_ _01919_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12272_ _06613_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__clkbuf_1
X_14011_ _07773_ _07774_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__nor2_1
XANTENNA__08918__A2 _03638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11223_ _05852_ _05860_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09040__A1 mem_rdata_q\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09256__S _03757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11154_ _05292_ net109 _04745_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__mux2_1
XANTENNA__16310__A0 _06984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13124__A0 _06947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10105_ reg_pc\[20\] decoded_imm\[20\] VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11085_ _03591_ _05760_ _05363_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__mux2_1
X_15962_ _02674_ _02676_ _02681_ _02682_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__o211a_1
XANTENNA__13675__A1 _07304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17701_ clknet_leaf_75_clk _00870_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dfxtp_1
X_10036_ net76 VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__clkbuf_4
X_14913_ net222 net191 _01824_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__mux2_1
XANTENNA__09974__S0 _04057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15893_ instr_sb _02635_ _02636_ is_sb_sh_sw VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__a22o_1
XANTENNA__11237__D _05871_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15932__D mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16613__A1 _06104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ clknet_leaf_172_clk _00801_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_14844_ count_cycle\[49\] count_cycle\[50\] _01780_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_86_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11438__B1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17563_ clknet_leaf_165_clk _00732_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14775_ count_cycle\[27\] _01732_ _01723_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_102_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11987_ _06445_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__clkbuf_1
X_16514_ _02967_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__clkbuf_8
X_13726_ _05013_ decoded_imm\[25\] VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10938_ _05620_ _05301_ _05484_ _05601_ _05624_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_82_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17494_ clknet_leaf_98_clk _00663_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15275__S1 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15900__A_N _03940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16445_ _02953_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__clkbuf_1
X_13657_ _07459_ _07503_ _07490_ _07474_ VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__a211o_1
XANTENNA__08773__A_N net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10869_ _05278_ _05559_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__nor2_1
XANTENNA__09939__B _04659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12608_ _06793_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16376_ _06982_ cpuregs.regs\[16\]\[19\] _02907_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__mux2_1
X_13588_ _07217_ _07438_ _07439_ _07190_ VGND VGND VPWR VPWR _07440_ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18115_ clknet_leaf_82_clk _01219_ VGND VGND VPWR VPWR timer\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09020__A _03747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15327_ cpuregs.regs\[8\]\[14\] cpuregs.regs\[9\]\[14\] cpuregs.regs\[10\]\[14\]
+ cpuregs.regs\[11\]\[14\] _01996_ _01997_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12539_ cpuregs.regs\[2\]\[4\] _06542_ _06752_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18046_ clknet_leaf_77_clk _00024_ VGND VGND VPWR VPWR irq_pending\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15258_ cpuregs.regs\[0\]\[10\] cpuregs.regs\[1\]\[10\] cpuregs.regs\[2\]\[10\] cpuregs.regs\[3\]\[10\]
+ _01990_ _01992_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14580__B _07956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14209_ irq_state\[0\] _07913_ VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15189_ cpuregs.regs\[0\]\[7\] cpuregs.regs\[1\]\[7\] cpuregs.regs\[2\]\[7\] cpuregs.regs\[3\]\[7\]
+ _03670_ _03671_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__mux4_1
XANTENNA__15104__A1 _03677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11709__B _06118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09582__A2 _04008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09750_ _04054_ _04475_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__nand2_1
X_08701_ net114 net82 VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__or2_1
X_09681_ cpuregs.regs\[20\]\[8\] cpuregs.regs\[21\]\[8\] cpuregs.regs\[22\]\[8\] cpuregs.regs\[23\]\[8\]
+ _04056_ _04091_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__mux4_1
XFILLER_0_146_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11141__A2 _05286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08632_ _03402_ _03403_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08563_ irq_mask\[24\] irq_pending\[24\] VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__and2b_1
XANTENNA__16727__S _03098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16368__A0 _06974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08494_ net66 VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10791__A2_N _05440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10652__A1 _05281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08753__B net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13151__S _07093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08472__C instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09115_ _03850_ _03791_ _03792_ _03849_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12990__S _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09046_ _03231_ _03807_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_758 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15894__A2 _02635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10804__A _05498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10263__S0 _04071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09948_ _03297_ _04361_ _04668_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__a21o_1
XANTENNA__10015__S _04064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ net71 VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__clkbuf_4
X_11910_ _06404_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12230__S _06576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12890_ _06104_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__buf_2
XFILLER_0_99_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10891__A1 _05414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09708__S0 _04274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11841_ _06366_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12093__A0 _06132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _06252_ _03354_ _06253_ _06317_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14560_ _07998_ _08209_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10723_ _05310_ _05314_ _05295_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__mux2_1
X_13511_ _04342_ _04611_ _07315_ VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08931__S1 _03684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14491_ _08140_ _08152_ _08150_ VGND VGND VPWR VPWR _08154_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15031__B1 _03240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16230_ _02839_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15582__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13442_ _07209_ VGND VGND VPWR VPWR _07304_ sky130_fd_sc_hd__clkbuf_4
X_10654_ instr_xor instr_xori VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__nor2_2
XFILLER_0_125_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13373_ _03312_ _04262_ _07236_ _07238_ VGND VGND VPWR VPWR _07239_ sky130_fd_sc_hd__a31o_1
X_16161_ net273 net235 _02797_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__mux2_1
X_10585_ _05287_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__16372__S _02907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09261__B2 _03888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15112_ _05255_ _01906_ _01967_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12324_ cpuregs.regs\[26\]\[0\] _06531_ _06641_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15334__B2 _02037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16092_ _03781_ _03935_ _02756_ _05987_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__a211o_1
XFILLER_0_161_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13345__B1 _07211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13297__A _07153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15043_ _05200_ _01863_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__nor2_1
X_12255_ cpuregs.regs\[25\]\[0\] _06531_ _06604_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__mux2_1
XANTENNA__12405__S _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11206_ _04342_ _05846_ _05827_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__mux2_1
X_12186_ _06183_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15098__B1 decoded_imm\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_79_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11137_ _04030_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__inv_2
X_16994_ clknet_leaf_181_clk _00168_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09714__S _04223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18733_ net128 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10006__S0 _04072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11068_ _05530_ _05700_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__nor2_1
X_15945_ _02664_ _02668_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__nor2_2
XANTENNA__13236__S _07140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15017__A _03240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10019_ _04737_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__inv_2
XANTENNA__10331__B1 _04009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15876_ _03790_ _03816_ _02628_ _02629_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17615_ clknet_leaf_145_clk _00784_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16062__A2 decoded_imm_j\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14827_ count_cycle\[43\] _01768_ count_cycle\[44\] VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__a21o_1
X_18595_ clknet_leaf_149_clk _01660_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16547__S _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15270__B1 _02118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17546_ clknet_leaf_182_clk _00715_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_14758_ count_cycle\[22\] _01722_ _01717_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_931 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14575__B _07956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13709_ _07524_ _07549_ VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17477_ clknet_leaf_2_clk _00646_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08922__S1 _03684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14689_ _03240_ VGND VGND VPWR VPWR _08335_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16428_ _06966_ cpuregs.regs\[29\]\[11\] _02943_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13584__B1 _03311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16359_ _02908_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16282__S _02859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_1010 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10398__B1 net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14591__A _07958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11595__C1 _06118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10937__A2 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18029_ clknet_leaf_65_clk _00005_ VGND VGND VPWR VPWR irq_pending\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15420__S1 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12315__S _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_97_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09802_ irq_mask\[11\] _04308_ timer\[11\] instr_timer _04025_ VGND VGND VPWR VPWR
+ _04527_ sky130_fd_sc_hd__a221o_1
XANTENNA__15626__S _03666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10570__A0 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09307__A2 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09733_ _03385_ _04454_ _04455_ _04459_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08748__B net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12311__A1 _06590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16038__C1 _02634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12050__S _06471_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16589__A0 _06991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09664_ reg_pc\[8\] decoded_imm\[8\] VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__nand2_1
XANTENNA__10873__A1 _05287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08615_ is_lb_lh_lw_lbu_lhu _03269_ _03388_ _03389_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__or4_1
XANTENNA__15487__S1 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09595_ _04273_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16457__S _02954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15361__S _01984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12075__A0 _06328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ irq_mask\[26\] irq_pending\[26\] VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__and2b_1
XANTENNA__08764__A net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10625__A1 _05255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15239__S1 _01986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10625__B2 _05225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08477_ instr_sll instr_sub instr_add instr_andi VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__or4_1
XFILLER_0_119_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15564__A1 _01969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12378__A1 _06588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10389__B1 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09243__A1 _03891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09595__A _04273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10370_ irq_pending\[27\] _04007_ _05075_ _05078_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__o22a_1
XANTENNA__10484__S0 _04274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09029_ net46 mem_rdata_q\[21\] _03729_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__mux2_1
XANTENNA__15411__S1 _03671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12040_ _06193_ cpuregs.regs\[22\]\[12\] _06471_ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10561__A0 _04754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08939__A _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13991_ count_instr\[2\] count_instr\[1\] count_instr\[0\] _07755_ VGND VGND VPWR
+ VPWR _07761_ sky130_fd_sc_hd__and4_1
XANTENNA__13056__S _07046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15730_ timer\[19\] _02533_ _02488_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12942_ _06247_ VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__buf_2
XFILLER_0_99_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15478__S1 _01937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15661_ _03301_ _04024_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__nand2_2
X_12873_ _06936_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_110 reg_next_pc\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13580__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17400_ clknet_leaf_164_clk _00569_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14612_ _08219_ _08231_ _08241_ _08254_ VGND VGND VPWR VPWR _08265_ sky130_fd_sc_hd__or4_1
X_11824_ _06357_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__clkbuf_1
X_18380_ clknet_leaf_163_clk _01445_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13802__A1 _05044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15592_ cpuregs.regs\[28\]\[29\] cpuregs.regs\[29\]\[29\] cpuregs.regs\[30\]\[29\]
+ cpuregs.regs\[31\]\[29\] _01908_ _01909_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__mux4_1
XANTENNA__08674__A net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11813__A0 _06114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17331_ clknet_leaf_165_clk _00505_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_14543_ _08198_ _08200_ VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__nand2_1
X_11755_ _06226_ reg_next_pc\[26\] _06300_ _06302_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__a211o_2
XFILLER_0_83_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10706_ _03528_ _05398_ _05400_ _05404_ _05405_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__o221a_1
XANTENNA__10092__A2 _04788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17262_ clknet_leaf_97_clk _00436_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14474_ _08133_ _08135_ _08138_ _07905_ reg_next_pc\[13\] VGND VGND VPWR VPWR _01005_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_153_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11686_ _06241_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16213_ _03218_ _02685_ _02827_ _02829_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__a211o_2
X_13425_ net93 decoded_imm\[4\] VGND VGND VPWR VPWR _07288_ sky130_fd_sc_hd__nor2_1
X_10637_ _05300_ _05338_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17193_ clknet_leaf_135_clk _00367_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12924__A _06200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09234__B2 _03888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11577__C1 _06118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16144_ net265 net227 _02786_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__mux2_1
X_10568_ _05044_ _05076_ _05263_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__mux2_1
X_13356_ _03316_ _07222_ _03281_ VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08993__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15858__A2 _02611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12307_ cpuregs.regs\[25\]\[25\] _06586_ _06626_ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__mux2_1
XANTENNA__12135__S _06518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16075_ decoded_imm\[25\] _02750_ _02746_ mem_rdata_q\[25\] _02749_ VGND VGND VPWR
+ VPWR _01338_ sky130_fd_sc_hd__a221o_1
X_10499_ _04010_ _05183_ _05203_ _03302_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__o211a_1
X_13287_ _06974_ cpuregs.regs\[5\]\[15\] _07165_ VGND VGND VPWR VPWR _07171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15026_ irq_mask\[22\] _01880_ _01895_ _01891_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__a211o_1
XANTENNA__11259__B _05889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15954__B net299 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12238_ _06319_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11974__S _06435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13755__A _05069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12169_ _06545_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__clkbuf_1
X_16977_ clknet_leaf_161_clk _00151_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14294__B2 _07960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 irq[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
XANTENNA__15970__A mem_rdata_q\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15928_ instr_or _02617_ _02626_ _02653_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__a22o_1
XANTENNA__16035__A2 _02711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15469__S1 _02070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18647_ clknet_leaf_112_clk _01707_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_15859_ _02616_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12057__A0 _06257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09380_ _04045_ _04113_ _04114_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__and3b_1
XFILLER_0_143_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15794__A1 latched_branch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18578_ clknet_leaf_128_clk _01643_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17529_ clknet_leaf_114_clk _00698_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10619__A instr_sub VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09473__A1 _04018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15546__A1 _03675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16743__B1 _01929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13557__A0 _04611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11884__S _06387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13665__A _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15157__S0 _01970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08759__A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14285__A1 reg_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14285__B2 _07960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11185__A _03219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09716_ cpuregs.regs\[16\]\[9\] cpuregs.regs\[17\]\[9\] cpuregs.regs\[18\]\[9\] cpuregs.regs\[19\]\[9\]
+ _04072_ _04074_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09647_ _04124_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_26_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08494__A net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09578_ irq_mask\[5\] _04308_ timer\[5\] _04023_ _04026_ VGND VGND VPWR VPWR _04309_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_26_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08529_ is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__buf_4
XFILLER_0_154_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08898__S0 _03661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11540_ reg_pc\[2\] _06090_ reg_pc\[3\] VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11471_ irq_mask\[23\] _03428_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13210_ _07130_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__clkbuf_1
X_10422_ _04070_ _05128_ _04082_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14190_ _03293_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_59_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10231__C1 _04149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13141_ _06963_ cpuregs.regs\[4\]\[10\] _07093_ VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__mux2_1
X_10353_ cpuregs.regs\[0\]\[27\] cpuregs.regs\[1\]\[27\] cpuregs.regs\[2\]\[27\] cpuregs.regs\[3\]\[27\]
+ _04207_ _04208_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__mux4_1
XFILLER_0_104_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15396__S0 _02046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13072_ _07045_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__clkbuf_8
X_10284_ _04430_ _04994_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__or2_1
X_12023_ _06125_ cpuregs.regs\[22\]\[4\] _06460_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__mux2_1
XANTENNA__15266__S _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16900_ clknet_leaf_31_clk _00045_ VGND VGND VPWR VPWR mem_rdata_q\[19\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13720__B1 _07211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13575__A _03387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17880_ clknet_leaf_88_clk _01049_ VGND VGND VPWR VPWR count_cycle\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10534__A0 _04036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08669__A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16831_ _06546_ cpuregs.regs\[14\]\[6\] _03152_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__mux2_1
XANTENNA__14276__A1 reg_pc\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14276__B2 _07960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16762_ _03122_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__clkbuf_1
X_13974_ _07737_ _07748_ VGND VGND VPWR VPWR _07749_ sky130_fd_sc_hd__and2_1
X_18501_ clknet_leaf_138_clk _01566_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_15713_ _04631_ _02477_ _02522_ _07775_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__a211oi_1
X_12925_ _06970_ cpuregs.regs\[31\]\[13\] _06964_ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__mux2_1
XANTENNA_output212_A net212 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16693_ _06959_ cpuregs.regs\[19\]\[8\] _03076_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18432_ clknet_leaf_143_clk _01497_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_15644_ _02468_ _02470_ _02465_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__or3b_1
X_12856_ _06927_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14579__A2 _07956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08835__C _03600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18363_ clknet_leaf_179_clk _01428_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11807_ _06078_ cpuregs.regs\[11\]\[0\] _06348_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__mux2_1
XANTENNA__15014__B _01885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15575_ cpuregs.regs\[28\]\[28\] cpuregs.regs\[29\]\[28\] cpuregs.regs\[30\]\[28\]
+ cpuregs.regs\[31\]\[28\] _02030_ _02031_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__mux4_1
XANTENNA__14984__C1 _08335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12787_ _06890_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16825__S _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17314_ clknet_leaf_183_clk _00488_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16725__A0 _06991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14526_ _08182_ _08184_ _08186_ _07905_ reg_next_pc\[17\] VGND VGND VPWR VPWR _01009_
+ sky130_fd_sc_hd__a32o_1
X_11738_ _06226_ reg_next_pc\[24\] _06285_ _06287_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__a211o_2
XANTENNA__08663__C1 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15528__B2 _02037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18294_ clknet_leaf_5_clk _01362_ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17245_ clknet_leaf_187_clk _00419_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09207__A1 _03892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14457_ _08119_ _08122_ VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__nor2_1
X_11669_ _06071_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08851__B net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11014__A1 instr_sub VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13408_ _07224_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10448__S0 _04472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17176_ clknet_leaf_176_clk _00350_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_14388_ reg_next_pc\[6\] _07905_ _08051_ _07899_ _08059_ VGND VGND VPWR VPWR _00998_
+ sky130_fd_sc_hd__a221o_1
X_16127_ net288 _05414_ _02771_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__mux2_1
X_13339_ _04054_ _07205_ _04296_ VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15387__S0 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16058_ _03402_ decoded_imm_j\[17\] _03403_ mem_rdata_q\[17\] VGND VGND VPWR VPWR
+ _02742_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_149_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13485__A net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09915__C1 _04149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15009_ irq_mask\[14\] _01880_ _01886_ _01876_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_166_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08880_ _03640_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_127_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09902__S _04078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09501_ _04091_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11733__A reg_pc\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_1006 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09432_ _03253_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15311__S0 _01990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08857__A_N _03604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13778__B1 _07211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14975__C1 _08335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09363_ cpuregs.raddr1\[1\] cpuregs.raddr1\[0\] VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__or2_1
XANTENNA__16735__S _03098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09294_ mem_wordsize\[2\] mem_wordsize\[1\] VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_10 _02298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_21 _04065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_32 _04923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_43 _06149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_54 is_alu_reg_reg VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16192__A1 net257 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08761__B net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_76 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_87 net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_98 _03346_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_183_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13379__B decoded_imm\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12753__A1 _06540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08421__A2 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15152__C1 _02006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput150 net150 VGND VGND VPWR VPWR eoi[27] sky130_fd_sc_hd__clkbuf_1
Xoutput161 net161 VGND VGND VPWR VPWR eoi[8] sky130_fd_sc_hd__clkbuf_1
XANTENNA__13395__A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput172 net172 VGND VGND VPWR VPWR mem_addr[19] sky130_fd_sc_hd__buf_1
Xoutput183 net183 VGND VGND VPWR VPWR mem_addr[2] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput194 net194 VGND VGND VPWR VPWR mem_la_addr[10] sky130_fd_sc_hd__buf_1
XANTENNA__08489__A is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11627__B _06118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14258__A1 _07899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14258__B2 reg_pc\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10971_ _05255_ _05394_ _05597_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__o21a_1
XANTENNA__09685__A1 _04231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15207__A0 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13481__A2 _05260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15115__A _01918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12710_ _06257_ cpuregs.regs\[12\]\[20\] _06847_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13690_ _07232_ _07529_ _07531_ _07533_ _07534_ VGND VGND VPWR VPWR _07535_ sky130_fd_sc_hd__o41a_1
XFILLER_0_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_136_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12641_ _06257_ cpuregs.regs\[30\]\[20\] _06810_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15360_ cpuregs.regs\[24\]\[16\] cpuregs.regs\[25\]\[16\] cpuregs.regs\[26\]\[16\]
+ cpuregs.regs\[27\]\[16\] _02022_ _02023_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08645__C1 _03304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12572_ _06751_ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__buf_6
XFILLER_0_65_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11789__S _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14311_ _07987_ VGND VGND VPWR VPWR _07988_ sky130_fd_sc_hd__buf_2
X_11523_ _06095_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__buf_2
XANTENNA__15605__S1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15291_ _02135_ _02136_ _02137_ _02138_ _01982_ _03683_ VGND VGND VPWR VPWR _02139_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__16183__A1 net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17030_ clknet_leaf_139_clk _00204_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14242_ reg_next_pc\[14\] _05876_ _07922_ _07936_ VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__o211a_2
XANTENNA__14194__B1 _07901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11454_ _06041_ irq_pending\[15\] _06045_ net7 VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12744__A1 cpuregs.waddr\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10405_ _05084_ _05085_ _05112_ VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12744__B2 _06861_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14173_ count_instr\[58\] count_instr\[57\] count_instr\[56\] _07881_ VGND VGND VPWR
+ VPWR _07887_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_74_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11385_ _03739_ _03923_ _05994_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13124_ _06947_ cpuregs.regs\[4\]\[2\] _07082_ VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__mux2_1
X_10336_ _04046_ _05044_ _04752_ _05045_ _04202_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14497__A1 _07899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15694__B1 _03240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_17932_ clknet_leaf_50_clk _08372_ VGND VGND VPWR VPWR reg_out\[12\] sky130_fd_sc_hd__dfxtp_1
X_13055_ _07048_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__clkbuf_1
X_10267_ _04966_ _04970_ _04978_ _04133_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__o211a_4
X_12006_ _06455_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__clkbuf_1
X_17863_ clknet_leaf_96_clk _01032_ VGND VGND VPWR VPWR count_cycle\[8\] sky130_fd_sc_hd__dfxtp_1
X_10198_ _04268_ _04890_ _04911_ _04149_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__o211a_1
XANTENNA__11180__A0 reg_next_pc\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10441__B decoded_imm\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16814_ _03149_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15541__S0 _03645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17794_ clknet_leaf_22_clk _00963_ VGND VGND VPWR VPWR reg_pc\[2\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_161_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16745_ _03680_ _01955_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_89_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13957_ _03304_ VGND VGND VPWR VPWR _07737_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09676__A1 _04053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13244__S _07140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15025__A _04908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12908_ _06156_ VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__buf_2
X_16676_ _03075_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09140__A3 _03880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13888_ _03344_ _07678_ _07682_ net156 VGND VGND VPWR VPWR _07689_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_122_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15627_ _00068_ _02455_ _03657_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__a21o_1
X_18415_ clknet_leaf_109_clk _01480_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12839_ _06184_ cpuregs.regs\[6\]\[11\] _06917_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16555__S _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10038__A2 _04104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18346_ clknet_leaf_30_clk _01414_ VGND VGND VPWR VPWR mem_rdata_q\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10669__S0 _05230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15558_ cpuregs.regs\[24\]\[27\] cpuregs.regs\[25\]\[27\] cpuregs.regs\[26\]\[27\]
+ cpuregs.regs\[27\]\[27\] _02069_ _02070_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14509_ _08161_ _08163_ _08170_ VGND VGND VPWR VPWR _08171_ sky130_fd_sc_hd__a21o_1
X_18277_ clknet_leaf_28_clk _01347_ VGND VGND VPWR VPWR is_slli_srli_srai sky130_fd_sc_hd__dfxtp_2
XFILLER_0_4_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15489_ cpuregs.regs\[12\]\[23\] cpuregs.regs\[13\]\[23\] cpuregs.regs\[14\]\[23\]
+ cpuregs.regs\[15\]\[23\] _03661_ _03662_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__mux4_1
XFILLER_0_83_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08581__B _03357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14185__B1 _07826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17228_ clknet_leaf_151_clk _00402_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 irq[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_2
XFILLER_0_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput41 mem_rdata[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
XANTENNA__15921__A1 is_alu_reg_reg VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput52 mem_rdata[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
XANTENNA__15921__B2 _05517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput63 mem_rdata[8] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11538__A2 reg_next_pc\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17159_ clknet_leaf_144_clk _00333_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09981_ _04231_ _04696_ _04700_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12499__A0 _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08932_ cpuregs.regs\[28\]\[3\] cpuregs.regs\[29\]\[3\] cpuregs.regs\[30\]\[3\] cpuregs.regs\[31\]\[3\]
+ _03641_ _03684_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08863_ instr_bne _03624_ _03627_ _03628_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13943__A _07677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08794_ _03496_ _03499_ _03556_ _03559_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__a31o_1
XANTENNA__15532__S0 _01995_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09116__A0 mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11474__A1 _06054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09762__S1 _04469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09415_ _03301_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__16465__S _02954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14412__A1 _03294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09868__A _04133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09346_ _04080_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_33_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16165__A1 net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09277_ _04013_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__buf_4
XFILLER_0_117_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15599__S0 _01908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14176__B1 _07826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11170_ _04038_ _05292_ net101 _03297_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__a22o_1
XANTENNA__10201__A2 _04913_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10121_ cpuregs.regs\[20\]\[20\] cpuregs.regs\[21\]\[20\] cpuregs.regs\[22\]\[20\]
+ cpuregs.regs\[23\]\[20\] _04282_ _04285_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__18131__D alu_out\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12233__S _06576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_42_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10052_ cpuregs.regs\[4\]\[18\] cpuregs.regs\[5\]\[18\] cpuregs.regs\[6\]\[18\] cpuregs.regs\[7\]\[18\]
+ _04472_ _04473_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__mux4_1
XANTENNA__11162__A0 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15428__A0 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14860_ count_cycle\[55\] _01792_ _01714_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15979__A1 _04024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15523__S0 _02069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14668__B _07969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13811_ cpuregs.regs\[0\]\[2\] VGND VGND VPWR VPWR _07645_ sky130_fd_sc_hd__clkbuf_1
X_14791_ _01747_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08666__B net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13064__S _07046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16530_ _02998_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13742_ _05013_ _05258_ VGND VGND VPWR VPWR _07583_ sky130_fd_sc_hd__nor2_1
XANTENNA__10268__A2 _04308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10954_ _05361_ _05631_ _05632_ _05639_ VGND VGND VPWR VPWR alu_out\[18\] sky130_fd_sc_hd__a31o_1
XANTENNA__09753__S1 _04478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16461_ _06999_ cpuregs.regs\[29\]\[27\] _02954_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__mux2_1
X_13673_ _04848_ _05258_ VGND VGND VPWR VPWR _07519_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10885_ _05278_ _05437_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_191_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_191_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_84_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14684__A _08232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18200_ clknet_leaf_42_clk _01271_ VGND VGND VPWR VPWR instr_xori sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_51_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15412_ cpuregs.regs\[0\]\[19\] cpuregs.regs\[1\]\[19\] cpuregs.regs\[2\]\[19\] cpuregs.regs\[3\]\[19\]
+ _03670_ _03671_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_14_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12624_ _06193_ cpuregs.regs\[30\]\[12\] _06799_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16392_ _02925_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_100_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08682__A net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18131_ clknet_leaf_40_clk alu_out\[5\] VGND VGND VPWR VPWR alu_out_q\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15343_ cpuregs.regs\[16\]\[15\] cpuregs.regs\[17\]\[15\] cpuregs.regs\[18\]\[15\]
+ cpuregs.regs\[19\]\[15\] _01996_ _01997_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12555_ _06765_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16156__A1 net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09291__C1 _04027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18062_ clknet_leaf_73_clk _01167_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dfxtp_4
XANTENNA__14167__B1 _07826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11506_ _06079_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__buf_4
XFILLER_0_81_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15274_ cpuregs.regs\[0\]\[11\] cpuregs.regs\[1\]\[11\] cpuregs.regs\[2\]\[11\] cpuregs.regs\[3\]\[11\]
+ _02085_ _02086_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__mux4_1
X_12486_ _06728_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17013_ clknet_leaf_117_clk _00187_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_14225_ _05857_ _06159_ _07922_ _05859_ VGND VGND VPWR VPWR _07925_ sky130_fd_sc_hd__o211a_2
X_11437_ irq_mask\[8\] _06030_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16404__A _02931_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09717__S _04078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output87_A net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14156_ _07874_ _07875_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11368_ _03215_ _05970_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_60_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15667__B1 _02488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _07075_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12143__S _06518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10319_ cpuregs.regs\[8\]\[26\] cpuregs.regs\[9\]\[26\] cpuregs.regs\[10\]\[26\]
+ cpuregs.regs\[11\]\[26\] _04071_ _04073_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__mux4_1
X_14087_ count_instr\[32\] _07824_ _07826_ VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__a21oi_1
X_11299_ reg_next_pc\[24\] _05898_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_163_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17915_ clknet_leaf_82_clk _01084_ VGND VGND VPWR VPWR count_cycle\[60\] sky130_fd_sc_hd__dfxtp_1
X_13038_ cpuregs.regs\[3\]\[26\] _06588_ _07032_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__mux2_1
XANTENNA__10171__B decoded_imm\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09441__S0 _04071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13693__A2 _05261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11982__S _06435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10900__A0 _04642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17846_ clknet_leaf_63_clk _01015_ VGND VGND VPWR VPWR reg_next_pc\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_124_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17777_ clknet_leaf_86_clk _00946_ VGND VGND VPWR VPWR count_instr\[48\] sky130_fd_sc_hd__dfxtp_1
X_14989_ irq_mask\[6\] _01864_ _01874_ _08335_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__a211o_1
XANTENNA__08576__B _03352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14297__C irq_pending\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16728_ _03103_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16659_ cpuregs.regs\[1\]\[24\] _06288_ _03062_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_182_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_182_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09200_ mem_rdata_q\[9\] _03826_ _03846_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08592__A _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09131_ _03861_ _03877_ _03887_ _03888_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__a22o_1
X_18329_ clknet_leaf_37_clk _01397_ VGND VGND VPWR VPWR mem_16bit_buffer\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08624__A2 _03385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09062_ net50 mem_rdata_q\[25\] _03729_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13381__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15107__C1 _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13149__S _07093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09964_ _04681_ _04682_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_984 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10290__S1 _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08915_ _03312_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__14330__B1 _07988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15872__B _02613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11144__B1 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09895_ _04214_ _04616_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__nand2_1
XANTENNA__12988__S _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11892__S _06387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13673__A _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10512__D _05215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08846_ _03610_ _03611_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__nor2_1
XANTENNA__10042__S1 _04759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15505__S0 _01990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08767__A net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08777_ net125 net93 VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__and2b_1
XANTENNA__14633__A1 _07899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_108_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_173_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_173_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09598__A _04052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10670_ net73 net74 _05229_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09329_ _04063_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__buf_8
XANTENNA__16138__A1 net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12340_ cpuregs.regs\[26\]\[8\] _06550_ _06641_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_985 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_117_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12271_ cpuregs.regs\[25\]\[8\] _06550_ _06604_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14010_ count_instr\[8\] _07771_ _07759_ VGND VGND VPWR VPWR _07774_ sky130_fd_sc_hd__o21ai_1
X_11222_ reg_out\[9\] _05857_ _05859_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09671__S0 _04072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11368__A _03215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11153_ _05811_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__buf_2
X_10104_ _04683_ _04716_ _04815_ _04819_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__a31oi_1
X_11084_ _05759_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__inv_2
X_15961_ mem_state\[0\] _02677_ _03227_ _02676_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__or4_1
XANTENNA__13675__A2 _04871_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17700_ clknet_leaf_75_clk _00869_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dfxtp_1
X_10035_ net42 _04710_ _04667_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__a21o_1
X_14912_ _01830_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__clkbuf_1
X_15892_ instr_lhu _02635_ _02625_ _02640_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__a22o_1
XANTENNA__09974__S1 _04060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08677__A net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ count_cycle\[49\] _01780_ _01782_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__o21a_1
X_17631_ clknet_leaf_163_clk _00800_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output125_A net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17562_ clknet_leaf_106_clk _00731_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_14774_ _01735_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_102_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11986_ _06248_ cpuregs.regs\[21\]\[19\] _06435_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16513_ _02989_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__clkbuf_1
X_13725_ net84 decoded_imm\[25\] VGND VGND VPWR VPWR _07567_ sky130_fd_sc_hd__or2_1
X_10937_ _03487_ _05222_ _05215_ _03488_ _05623_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17493_ clknet_leaf_100_clk _00662_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_164_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_164_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__12927__A _06207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16444_ _06982_ cpuregs.regs\[29\]\[19\] _02943_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__mux2_1
X_13656_ _07445_ _07460_ VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__or2b_1
XFILLER_0_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10868_ _05290_ _05306_ _05331_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09301__A _04036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12607_ _06125_ cpuregs.regs\[30\]\[4\] _06788_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16375_ _02916_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16129__A1 _05255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13587_ _04611_ _05259_ _07389_ _07254_ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__o211a_1
XANTENNA__09803__A1 instr_retirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16833__S _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10799_ _03512_ _03549_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18114_ clknet_leaf_82_clk _01218_ VGND VGND VPWR VPWR timer\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11071__C1 _05251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15326_ _02168_ _02169_ _02170_ _02171_ _01982_ _03639_ VGND VGND VPWR VPWR _02172_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10413__A2 _04016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12538_ _06756_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09020__B _03781_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18045_ clknet_leaf_82_clk _00022_ VGND VGND VPWR VPWR irq_pending\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13758__A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10881__S _05264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15257_ _02020_ _02106_ _02006_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12469_ _06719_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14208_ reg_next_pc\[4\] _06117_ _03189_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15188_ cpuregs.regs\[4\]\[7\] cpuregs.regs\[5\]\[7\] cpuregs.regs\[6\]\[7\] cpuregs.regs\[7\]\[7\]
+ _03670_ _03671_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14139_ _07862_ _07863_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15104__A2 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14312__B1 _07901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08700_ _03464_ _03465_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__and2b_1
XANTENNA__13493__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12874__A0 _06320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12601__S _06788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09680_ _04406_ _04407_ _04078_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__mux2_1
XANTENNA__08587__A instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08631_ _03257_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__buf_2
X_17829_ clknet_leaf_57_clk _00998_ VGND VGND VPWR VPWR reg_next_pc\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15812__B1 _03965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08562_ irq_mask\[27\] irq_pending\[27\] VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__and2b_1
XFILLER_0_147_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08493_ _03275_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_155_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_155_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_162_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14379__B1 _08050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12048__S _06471_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09114_ _03870_ _03872_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__or2_1
XANTENNA__10404__A2 _04049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08472__D _03255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15867__B _03940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14771__B _08350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09045_ net58 mem_rdata_q\[3\] _03730_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12572__A _06751_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10168__A1 _03384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15883__A _02611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10263__S1 _04073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09947_ mem_wordsize\[2\] mem_wordsize\[1\] VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__nor2_4
XANTENNA__15500__C1 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09405__S0 _04123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13607__S _07374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10820__A _05292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09878_ _04535_ _04542_ _04599_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_5_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16210__C _03215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08829_ net122 net90 VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__and2b_1
XFILLER_0_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12617__A0 _06166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11840_ _06224_ cpuregs.regs\[11\]\[16\] _06359_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__mux2_1
XANTENNA__09708__S1 _04317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11771_ reg_out\[28\] alu_out_q\[28\] _06069_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_146_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_146_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_64_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13510_ _07365_ _07366_ VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10722_ net126 _04262_ _05222_ _05420_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__a31o_1
X_14490_ _08140_ _08150_ _08152_ VGND VGND VPWR VPWR _08153_ sky130_fd_sc_hd__or3_1
XFILLER_0_83_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09121__A _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13441_ _03275_ _07299_ _07300_ _07302_ VGND VGND VPWR VPWR _07303_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10653_ net121 net89 VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__and2_1
XANTENNA__15582__A2 _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16653__S _03062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_637 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16160_ _02798_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__clkbuf_1
X_13372_ _07237_ VGND VGND VPWR VPWR _07238_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_840 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10584_ _05244_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11797__S _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09892__S0 _04290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15111_ _03396_ _03726_ _01966_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12323_ _06640_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_161_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16091_ _03878_ _02607_ _02755_ _03783_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__and4b_1
XFILLER_0_106_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15042_ irq_mask\[30\] _01865_ _01903_ _01891_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__a211o_1
XANTENNA__13345__B2 reg_next_pc\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12254_ _06603_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10159__A1 _04010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09644__S0 _04325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15793__A _03302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11205_ _05844_ _05845_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__and2b_1
XFILLER_0_103_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12185_ _06556_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15098__B2 _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11136_ _04040_ _04033_ _04030_ _04422_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__a2bb2o_2
XANTENNA_output242_A net242 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16993_ clknet_leaf_183_clk _00167_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_18732_ net127 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10006__S1 _04074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11067_ _05529_ _05621_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__and2_1
X_15944_ mem_rdata_q\[20\] mem_rdata_q\[22\] mem_rdata_q\[23\] mem_rdata_q\[21\] VGND
+ VGND VPWR VPWR _02668_ sky130_fd_sc_hd__or4b_1
XANTENNA__14202__A _06860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10018_ _04724_ _04728_ net300 _04736_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__a211o_4
X_15875_ _03768_ _03916_ _02603_ _02608_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__and4b_1
XFILLER_0_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14826_ count_cycle\[43\] count_cycle\[44\] _01768_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__and3_1
X_17614_ clknet_leaf_136_clk _00783_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_18594_ clknet_leaf_159_clk _01659_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15270__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ _01722_ _01724_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__nor2_1
XANTENNA__13281__A0 _06968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17545_ clknet_leaf_185_clk _00714_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_137_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_137_clk sky130_fd_sc_hd__clkbuf_2
X_11969_ _06436_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13708_ _07499_ _07550_ _07511_ VGND VGND VPWR VPWR _07551_ sky130_fd_sc_hd__o21a_1
XANTENNA__15033__A _05037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17476_ clknet_leaf_7_clk _00645_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14688_ reg_next_pc\[31\] _07948_ _08326_ _08334_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__a22o_1
XANTENNA__15022__A1 _03303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10190__S0 _04084_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11280__B _05906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13639_ _07483_ _07485_ _07486_ _07284_ VGND VGND VPWR VPWR _07487_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_119_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16427_ _02944_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16358_ _06963_ cpuregs.regs\[16\]\[10\] _02907_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08870__A _03635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11595__B1 _06098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15309_ _02154_ _02155_ _01984_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12392__A _06677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16289_ _06963_ cpuregs.regs\[15\]\[10\] _02870_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18028_ clknet_leaf_65_clk _00004_ VGND VGND VPWR VPWR irq_pending\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09635__S0 _04274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10116__S _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09801_ _04227_ _04517_ _04525_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__nor3_4
XANTENNA__10570__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09732_ _03637_ _04456_ _04458_ _03225_ _04266_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__a221o_1
XANTENNA__12847__A0 _06216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09206__A _03730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09663_ _03385_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__clkbuf_4
X_08614_ _03271_ _03254_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__or2_1
X_09594_ cpuregs.regs\[4\]\[6\] cpuregs.regs\[5\]\[6\] cpuregs.regs\[6\]\[6\] cpuregs.regs\[7\]\[6\]
+ _04291_ _04292_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__mux4_1
XFILLER_0_173_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08545_ _03320_ _03321_ _03322_ _03323_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_46_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_128_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_128_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_119_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13162__S _07104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10086__B1 _04237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10625__A2 _05261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08476_ instr_fence instr_and _03257_ _03259_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__or4_1
XFILLER_0_147_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10181__S0 _04281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16473__S _02968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10389__A1 _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10484__S1 _04317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12506__S _06737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09028_ _03206_ _03213_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_130_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10561__A1 _04810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15118__A _01918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13990_ _07758_ _07760_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12941_ _06981_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16648__S _03051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15660_ _02482_ _02478_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__nand2_1
XANTENNA__15788__C1 _06026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_100 _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12872_ _06312_ cpuregs.regs\[6\]\[27\] _06928_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__mux2_1
XANTENNA_111 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_122 net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14611_ _07988_ _08263_ VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__nand2_1
XANTENNA__13580__B decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 _05517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _06157_ cpuregs.regs\[11\]\[8\] _06348_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _02420_ _02421_ _02110_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_119_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_119_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA_144 net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08674__B net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13802__A2 _05260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17330_ clknet_leaf_111_clk _00504_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14542_ _08198_ _08200_ VGND VGND VPWR VPWR _08201_ sky130_fd_sc_hd__or2_1
X_11754_ _06252_ _03325_ _06253_ _06301_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10705_ _03527_ _05221_ _05356_ _03529_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__o22a_1
X_17261_ clknet_leaf_97_clk _00435_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14473_ _06863_ _08137_ VGND VGND VPWR VPWR _08138_ sky130_fd_sc_hd__nand2_1
X_11685_ _06240_ cpuregs.regs\[10\]\[18\] _06176_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16383__S _02918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16212_ _03753_ _03223_ _02828_ _02821_ _01821_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__o311ai_1
X_13424_ net93 decoded_imm\[4\] VGND VGND VPWR VPWR _07287_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10636_ net67 net99 _05231_ _03242_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__a22o_1
X_17192_ clknet_leaf_133_clk _00366_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11577__B1 _06098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09865__S0 _04280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16143_ _02789_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__clkbuf_1
X_13355_ cpu_state\[2\] _07221_ _05211_ _03400_ VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10567_ _04959_ _05013_ _05236_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12416__S _06689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16504__A1 _06565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11320__S _03219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12306_ _06631_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16074_ decoded_imm\[24\] _02750_ _02746_ mem_rdata_q\[24\] _02749_ VGND VGND VPWR
+ VPWR _01337_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13286_ _07170_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__clkbuf_1
X_10498_ _04271_ _05201_ _05202_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15025_ _04908_ _01885_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__nor2_1
X_12237_ _06591_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16268__A0 _06941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12168_ cpuregs.regs\[24\]\[5\] _06544_ _06534_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__mux2_1
X_11119_ _03436_ _05222_ _05596_ _05254_ _05792_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__a221o_1
X_12099_ _06157_ cpuregs.regs\[23\]\[8\] _06496_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__mux2_1
X_16976_ clknet_leaf_164_clk _00150_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15927_ _02625_ _02651_ _02656_ _02616_ instr_sra VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__a32o_1
Xinput6 irq[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XANTENNA__15970__B mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10304__A1 _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10304__B2 _05014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09170__A1 _03920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13771__A net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18646_ clknet_leaf_168_clk _01706_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_15858_ _03309_ _02611_ _02615_ _02617_ instr_beq VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__a32o_1
XANTENNA__08865__A _03311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14809_ count_cycle\[37\] _01756_ count_cycle\[38\] VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__a21o_1
XANTENNA__09458__C1 _04150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18577_ clknet_leaf_119_clk _01642_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_15789_ _03385_ _03292_ _03318_ _06069_ _06026_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__o221a_1
XFILLER_0_148_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17528_ clknet_leaf_165_clk _00697_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_173_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17459_ clknet_leaf_151_clk _00628_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16293__S _02870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16743__B2 _03638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13557__A1 _04566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18224__D _01295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12326__S _06641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13665__B decoded_imm\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15157__S1 _01971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08759__B _03524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13157__S _07093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12061__S _06482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09715_ cpuregs.regs\[20\]\[9\] cpuregs.regs\[21\]\[9\] cpuregs.regs\[22\]\[9\] cpuregs.regs\[23\]\[9\]
+ _04072_ _04074_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__mux4_1
XANTENNA__12996__S _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09646_ _04373_ _04374_ _04321_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09577_ instr_maskirq VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_167_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ irq_mask\[1\] irq_active _03307_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__nor3_4
XFILLER_0_148_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08898__S1 _03662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08459_ _03242_ net67 VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13620__S _07374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11470_ _06053_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10421_ _05126_ _05127_ _04121_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12236__S _06576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13140_ _07081_ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10352_ cpuregs.regs\[4\]\[27\] cpuregs.regs\[5\]\[27\] cpuregs.regs\[6\]\[27\] cpuregs.regs\[7\]\[27\]
+ _04207_ _04208_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__mux4_1
XANTENNA__15396__S1 _02047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13071_ _07056_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__clkbuf_1
X_10283_ cpuregs.regs\[16\]\[25\] cpuregs.regs\[17\]\[25\] cpuregs.regs\[18\]\[25\]
+ cpuregs.regs\[19\]\[25\] _04291_ _04292_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13720__A1 _07209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12022_ _06464_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13720__B2 reg_pc\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13575__B _04631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10534__A1 _04160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08669__B net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16830_ _03158_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__clkbuf_1
X_13973_ _03337_ _07727_ _07728_ net152 VGND VGND VPWR VPWR _07748_ sky130_fd_sc_hd__a22o_1
X_16761_ _06544_ cpuregs.regs\[13\]\[5\] _03116_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__mux2_1
XANTENNA__09688__C1 _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18500_ clknet_leaf_143_clk _01565_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15282__S _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10298__B1 _04133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15712_ _02484_ _02520_ _02521_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__and3_1
X_12924_ _06200_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__buf_2
X_16692_ _03084_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08685__A net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10393__S0 _04123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18431_ clknet_leaf_133_clk _01496_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13236__A0 _06991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15643_ mem_do_prefetch _03410_ _02469_ _03301_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__a22o_1
X_12855_ _06248_ cpuregs.regs\[6\]\[19\] _06917_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__mux2_1
XANTENNA_output205_A net205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14579__A3 _08050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11806_ _06347_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__buf_6
XFILLER_0_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15574_ _02404_ _02405_ _03687_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__mux2_1
X_18362_ clknet_leaf_18_clk _01427_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12786_ cpuregs.regs\[9\]\[19\] _06573_ _06880_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10145__S0 _04758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11798__B1 _06098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17313_ clknet_leaf_184_clk _00487_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_14525_ _08120_ _08185_ VGND VGND VPWR VPWR _08186_ sky130_fd_sc_hd__or2_1
X_11737_ _06252_ _03342_ _06253_ _06286_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__a22o_1
XANTENNA__10696__S1 _05287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18293_ clknet_leaf_5_clk _01361_ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15084__S0 _03669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17244_ clknet_leaf_13_clk _00418_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_14456_ _07932_ _08102_ _08121_ VGND VGND VPWR VPWR _08122_ sky130_fd_sc_hd__o21ai_1
X_11668_ _06225_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13407_ _07270_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08415__A0 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11014__A2 _04913_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10619_ instr_sub VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17175_ clknet_leaf_156_clk _00349_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10448__S1 _04473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14387_ _08056_ _08057_ _08058_ VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__and3b_1
X_11599_ _06162_ _06163_ _06075_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_12_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16126_ _02780_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13338_ _07203_ _07204_ _04575_ VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15387__S1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11970__A0 _06184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15457__S _01907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16057_ decoded_imm\[16\] _02720_ _02736_ _02741_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__o22a_1
X_13269_ _07161_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_149_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15008_ _04631_ _01885_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__nor2_1
XANTENNA__13485__B decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15981__A _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16959_ clknet_leaf_180_clk _00133_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_127_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09500_ _04084_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_144_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10289__B1 _04225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09431_ _04151_ _04159_ _04164_ _04008_ irq_pending\[2\] VGND VGND VPWR VPWR _08391_
+ sky130_fd_sc_hd__o32a_2
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18629_ clknet_leaf_182_clk _01689_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15767__A2 _02560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15311__S1 _01992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13778__A1 _07304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13778__B2 reg_pc\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09362_ _04070_ _04090_ _04096_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_170_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09293_ _03242_ mem_wordsize\[2\] VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__nand2_4
XFILLER_0_170_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_11 _02397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_22 _04151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_33 _04982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10461__B1 _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_44 _06165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16192__A2 net259 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 mem_do_wdata VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09829__S0 _04329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_66 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_77 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_88 net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16751__S _03116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 _03880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15875__B _03916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11961__A0 _06150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput140 net140 VGND VGND VPWR VPWR eoi[18] sky130_fd_sc_hd__buf_1
Xoutput151 net151 VGND VGND VPWR VPWR eoi[28] sky130_fd_sc_hd__buf_1
XFILLER_0_100_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput162 net162 VGND VGND VPWR VPWR eoi[9] sky130_fd_sc_hd__buf_1
XANTENNA__13395__B decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput173 net173 VGND VGND VPWR VPWR mem_addr[20] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput184 net184 VGND VGND VPWR VPWR mem_addr[30] sky130_fd_sc_hd__clkbuf_1
Xoutput195 net195 VGND VGND VPWR VPWR mem_la_addr[11] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11196__A _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14258__A2 _07944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10970_ _03466_ _05653_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__xor2_1
XFILLER_0_168_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09629_ _04356_ _04357_ _04347_ _04351_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__o211a_1
XANTENNA__18129__D alu_out\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12640_ _06787_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12571_ _06773_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12441__A1 _06582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_50_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14310_ _03364_ _07986_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__and2_1
XANTENNA__15131__A _03647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11522_ _06066_ _06088_ _06089_ _06094_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__a211o_4
XFILLER_0_136_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15290_ cpuregs.regs\[8\]\[12\] cpuregs.regs\[9\]\[12\] cpuregs.regs\[10\]\[12\]
+ cpuregs.regs\[11\]\[12\] _02085_ _02086_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14241_ _05857_ _06205_ VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15391__B1 _02233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11453_ irq_mask\[15\] _06042_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__or2_1
XANTENNA__10275__A reg_pc\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14970__A _03301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16661__S _03062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10404_ irq_pending\[28\] _04049_ _05111_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12744__A2 _06862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14172_ _07886_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15785__B _03364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11384_ _03789_ _05992_ _05993_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_74_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13123_ _07084_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__clkbuf_1
X_10335_ net51 _04811_ _04667_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15694__A1 _02484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17931_ clknet_leaf_55_clk _08371_ VGND VGND VPWR VPWR reg_out\[11\] sky130_fd_sc_hd__dfxtp_1
X_13054_ _06945_ cpuregs.regs\[7\]\[1\] _07046_ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__mux2_1
X_10266_ _04328_ _04973_ _04977_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__a21o_1
XANTENNA_output155_A net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12005_ _06320_ cpuregs.regs\[21\]\[28\] _06446_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__mux2_1
X_17862_ clknet_leaf_93_clk _01031_ VGND VGND VPWR VPWR count_cycle\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10197_ _04271_ _04909_ _04910_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16813_ _06596_ cpuregs.regs\[13\]\[30\] _03115_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17793_ clknet_leaf_22_clk _00962_ VGND VGND VPWR VPWR reg_pc\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15541__S1 _03647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09125__B2 _03767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16744_ reg_sh\[0\] _07274_ _03111_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_89_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13956_ _07736_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_89_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09304__A _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15025__B _01885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12907_ _06958_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__clkbuf_1
X_13887_ _07688_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__clkbuf_1
X_16675_ _06346_ _02894_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_122_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14957__A0 net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18414_ clknet_leaf_107_clk _01479_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_15626_ _02453_ _02454_ _03666_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__mux2_1
X_12838_ _06918_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10118__S0 _04275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14864__B _01753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18345_ clknet_leaf_29_clk _01413_ VGND VGND VPWR VPWR mem_rdata_q\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10884__S _05288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12769_ _06881_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__clkbuf_1
X_15557_ _01984_ _02389_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16137__A _02770_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__13260__S _07154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15041__A _05169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14508_ _07972_ _08168_ _08169_ _08050_ _07941_ VGND VGND VPWR VPWR _08170_ sky130_fd_sc_hd__a32o_1
XANTENNA__14709__B1 _07826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15488_ _02323_ _02324_ _03653_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__mux2_1
X_18276_ clknet_leaf_29_clk _01346_ VGND VGND VPWR VPWR is_lb_lh_lw_lbu_lhu sky130_fd_sc_hd__dfxtp_2
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08581__C _03358_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput20 irq[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
XFILLER_0_141_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17227_ clknet_leaf_150_clk _00401_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput31 irq[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
X_14439_ _08104_ _08105_ VGND VGND VPWR VPWR _08106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 mem_rdata[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput53 mem_rdata[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
XFILLER_0_4_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput64 mem_rdata[9] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09061__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17158_ clknet_leaf_137_clk _00332_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_168_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16109_ mem_do_wdata _03220_ _01821_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__and3_1
X_09980_ _04069_ _04699_ _04095_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__a21o_1
X_17089_ clknet_leaf_183_clk _00263_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09185__S _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08931_ cpuregs.regs\[24\]\[3\] cpuregs.regs\[25\]\[3\] cpuregs.regs\[26\]\[3\] cpuregs.regs\[27\]\[3\]
+ _03641_ _03684_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08862_ instr_bgeu _03625_ _03599_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__mux2_1
XANTENNA__11171__A1 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08793_ _03496_ _03557_ _03558_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__a21o_1
XANTENNA__15532__S1 _01937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15988__A2 _03737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09116__A1 _03874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15216__A _02066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12120__A0 _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09414_ count_cycle\[2\] _04014_ _04147_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__a21o_1
XANTENNA__15296__S0 _01999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09345_ _00073_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__inv_2
XANTENNA__13620__A0 _04744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10029__A3 _04743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13170__S _07104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_2
X_09276_ _03253_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15599__S1 _01909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15373__B1 _02197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16481__S _02968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10198__C1 _04149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11934__A0 _06312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12514__S _06737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16873__A0 _06588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10120_ _04834_ _04835_ _04430_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_99_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10051_ _04430_ _04768_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__or2_1
XANTENNA__11162__A1 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15428__A1 _02268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09823__S _04369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10969__S _05363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15979__A2 _02635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15523__S1 _02070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13810_ _07644_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__clkbuf_1
X_14790_ _01745_ _08350_ _01746_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__and3b_1
XANTENNA__09658__A2 _04013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10348__S0 _04207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13741_ _07568_ _07571_ _07580_ VGND VGND VPWR VPWR _07582_ sky130_fd_sc_hd__nand3_1
X_10953_ _05337_ _05597_ _05635_ _05281_ _05638_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_1013 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10673__A0 _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15287__S0 _01970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13672_ _04744_ _07236_ _07517_ _07217_ VGND VGND VPWR VPWR _07518_ sky130_fd_sc_hd__o211a_1
X_16460_ _02961_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__clkbuf_1
X_10884_ _05570_ _05573_ _05288_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08963__A _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14684__B _07971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15411_ cpuregs.regs\[4\]\[19\] cpuregs.regs\[5\]\[19\] cpuregs.regs\[6\]\[19\] cpuregs.regs\[7\]\[19\]
+ _03670_ _03671_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__mux4_1
X_12623_ _06801_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_84_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08618__B1 _03244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12414__A1 _06554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16391_ _06997_ cpuregs.regs\[16\]\[26\] _02918_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08682__B net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_23_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_54_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18130_ clknet_leaf_27_clk alu_out\[4\] VGND VGND VPWR VPWR alu_out_q\[4\] sky130_fd_sc_hd__dfxtp_1
X_15342_ _02183_ _02184_ _02185_ _02186_ _02111_ _02088_ VGND VGND VPWR VPWR _02187_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_109_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12554_ cpuregs.regs\[2\]\[11\] _06557_ _06763_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10976__B2 _05251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11505_ cpuregs.waddr\[0\] cpuregs.waddr\[1\] VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__and2b_1
X_18061_ clknet_leaf_73_clk _01166_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dfxtp_4
X_15273_ cpuregs.regs\[4\]\[11\] cpuregs.regs\[5\]\[11\] cpuregs.regs\[6\]\[11\] cpuregs.regs\[7\]\[11\]
+ _01976_ _01977_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__mux4_1
X_12485_ _06184_ cpuregs.regs\[28\]\[11\] _06726_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__mux2_1
XANTENNA__16391__S _02918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17012_ clknet_leaf_112_clk _00186_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_14224_ reg_pc\[8\] _07906_ _07924_ _07912_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__a22o_1
X_11436_ _06029_ irq_pending\[7\] _06035_ net30 VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__a31o_1
XANTENNA__09043__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14155_ count_instr\[52\] _07872_ _07834_ VGND VGND VPWR VPWR _07875_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13390__A2 _04342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12424__S _06689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11367_ _05967_ _05979_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15211__S0 _01976_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13106_ _06997_ cpuregs.regs\[7\]\[26\] _07068_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__mux2_1
X_10318_ _04068_ _05027_ _04080_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_146_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14086_ _03239_ VGND VGND VPWR VPWR _07826_ sky130_fd_sc_hd__buf_4
X_11298_ _03460_ _05829_ _05921_ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__o21ai_4
XFILLER_0_119_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_163_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17914_ clknet_leaf_84_clk _01083_ VGND VGND VPWR VPWR count_cycle\[59\] sky130_fd_sc_hd__dfxtp_1
X_13037_ _07038_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__clkbuf_1
X_10249_ count_instr\[56\] _04015_ _04017_ count_cycle\[56\] VGND VGND VPWR VPWR _04961_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09441__S1 _04073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17845_ clknet_leaf_60_clk _01014_ VGND VGND VPWR VPWR reg_next_pc\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10900__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16092__A1 _03781_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17776_ clknet_leaf_87_clk _00945_ VGND VGND VPWR VPWR count_instr\[47\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_182_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14988_ _04335_ _01869_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__nor2_1
XANTENNA__08576__C _03353_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_9 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16727_ _06993_ cpuregs.regs\[19\]\[24\] _03098_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__mux2_1
X_13939_ _07724_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11456__A2 irq_pending\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16566__S _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15278__S0 _02069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09969__A _04054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16658_ _03066_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15609_ _02437_ _02438_ _02110_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16589_ _06991_ cpuregs.regs\[18\]\[23\] _03026_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_33_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09130_ _03835_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18328_ clknet_leaf_19_clk _01396_ VGND VGND VPWR VPWR cpuregs.waddr\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09282__B1 _04018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08624__A3 _03237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09061_ net64 mem_rdata_q\[9\] _03729_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__mux2_1
X_18259_ clknet_leaf_28_clk _01330_ VGND VGND VPWR VPWR decoded_imm\[17\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_72_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15450__S0 _02111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11739__A _06288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15107__B1 decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13381__A2 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12334__S _06641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15658__A1 _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15202__S0 _03640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09963_ _04681_ _04682_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_135_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08914_ cpuregs.raddr2\[3\] cpuregs.raddr2\[4\] _03678_ VGND VGND VPWR VPWR _03679_
+ sky130_fd_sc_hd__or3_4
X_09894_ _04614_ _04615_ _04222_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__mux2_1
XANTENNA__11144__A1 _03407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15872__C _03940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11144__B2 _04422_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08845_ net67 _03609_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__and2_1
XANTENNA__14968__A1_N irq_active VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11875__A_N _06082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_1002 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15505__S1 _01992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08767__B net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08776_ _03531_ net92 _03541_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__a21o_1
XANTENNA__14094__B1 _07790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14633__A2 _07964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09879__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09328_ _00071_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_75_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15346__B1 _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09259_ _03996_ _03997_ _03737_ _03932_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__o211a_1
XFILLER_0_173_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12270_ _06612_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11221_ reg_next_pc\[9\] _05858_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09671__S1 _04074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11152_ _05277_ net108 _04745_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__mux2_1
X_10103_ reg_pc\[19\] decoded_imm\[19\] _04815_ _04817_ _04818_ VGND VGND VPWR VPWR
+ _04819_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11083_ _03448_ _03451_ _05752_ _03447_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__a31o_1
X_15960_ _01821_ _02680_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__nand2_1
XANTENNA__11135__A1 _05219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10034_ _04673_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__buf_2
X_14911_ net221 net190 _01824_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__mux2_1
X_15891_ instr_lbu _02635_ _02623_ _02640_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__a22o_1
XANTENNA__16074__A1 decoded_imm\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08677__B net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13075__S _07057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17630_ clknet_leaf_124_clk _00799_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16074__B2 mem_rdata_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14842_ count_cycle\[49\] _01780_ _01714_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_19_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14624__A2 _07948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17561_ clknet_leaf_114_clk _00730_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_14773_ count_cycle\[25\] count_cycle\[26\] count_cycle\[27\] _01729_ VGND VGND VPWR
+ VPWR _01735_ sky130_fd_sc_hd__and4_1
X_11985_ _06444_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output118_A net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16512_ cpuregs.regs\[17\]\[19\] _06573_ _02979_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__mux2_1
XANTENNA__08934__S0 _03658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13724_ _07566_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__clkbuf_1
X_10936_ _05284_ _05622_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__nor2_1
X_17492_ clknet_leaf_152_clk _00661_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16443_ _02952_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13655_ _07450_ _07461_ _07474_ _07490_ VGND VGND VPWR VPWR _07502_ sky130_fd_sc_hd__or4_1
X_10867_ _05288_ _05422_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__nor2_1
XANTENNA__14388__B2 _07899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12606_ _06792_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13586_ _04532_ _04810_ _07315_ VGND VGND VPWR VPWR _07438_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16374_ _06980_ cpuregs.regs\[16\]\[18\] _02907_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10798_ _03550_ _04419_ _05322_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_156_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09803__A2 _04526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18113_ clknet_leaf_81_clk _01217_ VGND VGND VPWR VPWR timer\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15337__B1 _02181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15325_ cpuregs.regs\[16\]\[14\] cpuregs.regs\[17\]\[14\] cpuregs.regs\[18\]\[14\]
+ cpuregs.regs\[19\]\[14\] _02085_ _02086_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__mux4_1
X_12537_ cpuregs.regs\[2\]\[3\] _06540_ _06752_ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15432__S0 _01976_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18044_ clknet_leaf_76_clk _00021_ VGND VGND VPWR VPWR irq_pending\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13758__B decoded_imm\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15256_ _02104_ _02105_ _03687_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__mux2_1
X_12468_ _06114_ cpuregs.regs\[28\]\[3\] _06715_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09567__A1 _04272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11419_ _05969_ _03920_ _06024_ _05973_ cpuregs.raddr1\[4\] VGND VGND VPWR VPWR _06025_
+ sky130_fd_sc_hd__a32o_1
X_14207_ reg_pc\[3\] _07906_ _07911_ _07912_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__a22o_1
X_15187_ net127 _01906_ _02039_ _02040_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__o22a_1
X_12399_ cpuregs.regs\[27\]\[3\] _06540_ _06678_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14138_ count_instr\[47\] _07860_ _07834_ VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11993__S _06446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08790__A2 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14069_ count_instr\[27\] count_instr\[26\] _07811_ VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__and3_1
XANTENNA__11126__A1 _05517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__13493__B decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08630_ instr_jal VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__buf_2
X_17828_ clknet_leaf_57_clk _00997_ VGND VGND VPWR VPWR reg_next_pc\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15812__A1 decoded_imm_j\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08561_ _03324_ _03329_ _03334_ _03339_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__or4_4
X_17759_ clknet_leaf_90_clk _00928_ VGND VGND VPWR VPWR count_instr\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08925__S0 _03658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08492_ _03274_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10101__A2 decoded_imm\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14379__A1 _07986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15576__B1 _01968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15040__A2 _01865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09113_ _03862_ _03863_ _03810_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15867__C _02612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15423__S0 _03640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09044_ _03203_ _03805_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11038__B1_N _05254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11469__A _03277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09946_ _04666_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__buf_2
XANTENNA__09405__S1 _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _04535_ _04542_ _04599_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_5_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09730__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08828_ _03592_ net87 _03445_ _03593_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__a31o_1
XANTENNA__09730__B2 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14067__B1 _07775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08759_ net126 _03524_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11770_ _06314_ _06315_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__nor2_1
XANTENNA__09494__B1 _04225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _03523_ _05301_ _05215_ _03526_ _05419_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__a221o_1
XANTENNA__18137__D alu_out\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12239__S _06576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15031__A2 _01863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13440_ _04040_ _05259_ _07301_ _07216_ VGND VGND VPWR VPWR _07302_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10652_ _05281_ _05345_ _05353_ _05298_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09121__B _03213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09341__S0 _04072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13371_ cpu_state\[4\] _03313_ VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__and2_1
XANTENNA__15319__B1 _02027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10583_ _05266_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09892__S1 _04276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15414__S0 _01936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12322_ _06639_ _06532_ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15110_ is_slli_srli_srai cpuregs.raddr2\[4\] decoded_imm\[4\] _01932_ _01934_ VGND
+ VGND VPWR VPWR _01966_ sky130_fd_sc_hd__a221o_1
X_16090_ _03228_ _03815_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15041_ _05169_ _01863_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11379__A _03916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12253_ _06602_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_79_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11204_ _05831_ _05835_ _05840_ _05843_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__a31o_1
XANTENNA__09644__S1 _04277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12184_ cpuregs.regs\[24\]\[10\] _06554_ _06555_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11135_ _05219_ _05800_ _05807_ VGND VGND VPWR VPWR alu_out\[31\] sky130_fd_sc_hd__o21ai_2
XANTENNA__13594__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11108__A1 _05219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16992_ clknet_leaf_186_clk _00166_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08688__A net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13502__C1 _07283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18731_ net126 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_1
X_11066_ _05743_ VGND VGND VPWR VPWR alu_out\[26\] sky130_fd_sc_hd__clkbuf_1
X_15943_ _04018_ _02650_ _02665_ _02667_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__a22o_1
XANTENNA_output235_A net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16047__A1 mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10017_ _04070_ _04731_ _04735_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14058__B1 _07775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15874_ _03833_ _03770_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__nor2_1
XANTENNA__10331__A2 _04145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17613_ clknet_leaf_145_clk _00782_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13805__A0 _05174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14825_ count_cycle\[43\] _01768_ _01770_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__o21a_1
X_18593_ clknet_leaf_129_clk _01658_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08907__S0 _03670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ clknet_leaf_173_clk _00713_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ count_cycle\[21\] _01719_ _01723_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11968_ _06175_ cpuregs.regs\[21\]\[10\] _06435_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10095__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11292__A0 _04913_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13707_ _04880_ decoded_imm\[21\] VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__nor2_1
XANTENNA__15033__B _01885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10919_ _05281_ _05599_ _05601_ _05480_ _05606_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__a221o_1
X_17475_ clknet_leaf_16_clk _00644_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16844__S _03163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11899_ _06175_ cpuregs.regs\[20\]\[10\] _06398_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14687_ _08327_ _08328_ _08329_ _08333_ VGND VGND VPWR VPWR _08334_ sky130_fd_sc_hd__a211o_1
XANTENNA__15022__A2 _04022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10190__S1 _04086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16426_ _06963_ cpuregs.regs\[29\]\[10\] _02943_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__mux2_1
XANTENNA__09237__A0 mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13638_ _07281_ _04806_ _07282_ reg_pc\[19\] VGND VGND VPWR VPWR _07486_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16357_ _02895_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13569_ _07420_ _07421_ VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15308_ cpuregs.regs\[24\]\[13\] cpuregs.regs\[25\]\[13\] cpuregs.regs\[26\]\[13\]
+ cpuregs.regs\[27\]\[13\] _02022_ _02023_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08460__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16288_ _02858_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_132_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18027_ clknet_leaf_65_clk _00003_ VGND VGND VPWR VPWR irq_pending\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__14533__A1 _07986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15730__B1 _02488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15239_ cpuregs.regs\[28\]\[9\] cpuregs.regs\[29\]\[9\] cpuregs.regs\[30\]\[9\] cpuregs.regs\[31\]\[9\]
+ _01985_ _01986_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__mux4_1
XANTENNA__10193__A _04133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09635__S1 _04317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09800_ _04272_ _04520_ _04524_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09193__S _03757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_163_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09731_ _04420_ _04457_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16038__B2 mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09662_ _04156_ _04358_ _04359_ _04390_ VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_2_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15246__C1 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08613_ is_slli_srli_srai _03387_ is_jalr_addi_slti_sltiu_xori_ori_andi VGND VGND
+ VPWR VPWR _03388_ sky130_fd_sc_hd__or3_1
X_09593_ _04206_ _04322_ _04225_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08544_ irq_mask\[9\] irq_pending\[9\] VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__and2b_2
XFILLER_0_77_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10086__A1 _04328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15549__A0 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11471__B _03428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09571__S0 _04217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08475_ instr_sw instr_sh _03258_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12059__S _06482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10181__S1 _04470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13679__A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11130__S0 _05324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09243__A3 _03810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08451__A1 _03199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09027_ _03206_ _03213_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12522__S _06737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14288__B1 _07944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15485__C1 _01968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09929_ _04231_ _04649_ _04082_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10849__B1 _05367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12940_ _06980_ cpuregs.regs\[31\]\[18\] _06964_ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__mux2_1
XANTENNA__09831__S _04369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08911__C1 _03675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12871_ _06935_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_101 _04532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_123 net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15134__A _03666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14610_ _07961_ _08258_ VGND VGND VPWR VPWR _08263_ sky130_fd_sc_hd__and2_1
XANTENNA_134 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _06356_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15860__B_N _02612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15590_ cpuregs.regs\[16\]\[29\] cpuregs.regs\[17\]\[29\] cpuregs.regs\[18\]\[29\]
+ cpuregs.regs\[19\]\[29\] _02221_ _02222_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__mux4_1
XANTENNA_145 _04342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11753_ reg_out\[26\] alu_out_q\[26\] _06069_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09562__S0 _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14541_ _08180_ _08199_ _08187_ VGND VGND VPWR VPWR _08200_ sky130_fd_sc_hd__a21o_1
X_10704_ _05403_ _05247_ _05246_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__mux2_2
X_17260_ clknet_leaf_151_clk _00434_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13015__A1 _06565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11684_ _06239_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__buf_2
X_14472_ _08035_ _08136_ VGND VGND VPWR VPWR _08137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16211_ net33 net44 VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10635_ _05332_ _05336_ _05278_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__mux2_1
X_13423_ _07191_ _07275_ _07280_ _07285_ VGND VGND VPWR VPWR _07286_ sky130_fd_sc_hd__o31a_1
XANTENNA__13589__A _04659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17191_ clknet_leaf_144_clk _00365_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11577__A1 _06072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09865__S1 _04091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13354_ _07220_ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16142_ net264 net226 _02786_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10566_ _05268_ _05269_ _05266_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output185_A net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12305_ cpuregs.regs\[25\]\[24\] _06584_ _06626_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13285_ _06972_ cpuregs.regs\[5\]\[14\] _07165_ VGND VGND VPWR VPWR _07170_ sky130_fd_sc_hd__mux2_1
XANTENNA__10217__S _04065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16073_ decoded_imm\[23\] _02750_ _02746_ mem_rdata_q\[23\] _02749_ VGND VGND VPWR
+ VPWR _01336_ sky130_fd_sc_hd__a221o_1
X_10497_ irq_mask\[31\] _04021_ timer\[31\] _04023_ _04188_ VGND VGND VPWR VPWR _05202_
+ sky130_fd_sc_hd__a221o_1
X_15024_ _03303_ _04022_ _04871_ _01894_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__a31o_1
X_12236_ cpuregs.regs\[24\]\[27\] _06590_ _06576_ VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09942__B2 _03253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12432__S _06689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12167_ _06131_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__buf_2
X_11118_ _03435_ _05221_ _05356_ _03438_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__o22ai_1
X_12098_ _06504_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__clkbuf_1
X_16975_ clknet_leaf_120_clk _00149_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_11049_ _05513_ _05621_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__and2_1
X_15926_ _02625_ _02649_ _02651_ _02616_ instr_srl VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10304__A2 _05013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput7 irq[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_127_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13771__B decoded_imm\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18645_ clknet_leaf_111_clk _01705_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_15857_ _02616_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15779__B1 _07905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14808_ count_cycle\[37\] count_cycle\[38\] _01756_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18576_ clknet_leaf_108_clk _01641_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_135_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15788_ latched_store _02573_ _02577_ _06026_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__o211a_1
XANTENNA__10068__A1 reg_pc\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11291__B _05915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17527_ clknet_leaf_117_clk _00696_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_173_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14739_ count_cycle\[16\] count_cycle\[17\] _08365_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__and3_1
XANTENNA__16574__S _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17458_ clknet_leaf_147_clk _00627_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08881__A _00065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16409_ _06947_ cpuregs.regs\[29\]\[2\] _02932_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17389_ clknet_leaf_153_clk _00558_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12607__S _06788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11568__A1 _06116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_144_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16259__A1 _03878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12342__S _06641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13962__A _07737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09714_ _04439_ _04440_ _04223_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__mux2_1
X_09645_ cpuregs.regs\[24\]\[7\] cpuregs.regs\[25\]\[7\] cpuregs.regs\[26\]\[7\] cpuregs.regs\[27\]\[7\]
+ _04325_ _04317_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_153_Left_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09576_ _04227_ _04298_ _04306_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__nor3_4
XFILLER_0_96_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14442__B1 _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08527_ cpu_state\[2\] _03269_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_26_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15617__S0 _02046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08458_ net78 VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11008__A0 _04945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13548__A2 _07392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11559__A1 alu_out_q\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10420_ cpuregs.regs\[16\]\[29\] cpuregs.regs\[17\]\[29\] cpuregs.regs\[18\]\[29\]
+ cpuregs.regs\[19\]\[29\] _04477_ _04478_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__mux4_1
XANTENNA__08424__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_162_Left_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10231__A1 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10351_ _04215_ _05059_ _04225_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13070_ _06961_ cpuregs.regs\[7\]\[9\] _07046_ VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__mux2_1
X_10282_ cpuregs.regs\[20\]\[25\] cpuregs.regs\[21\]\[25\] cpuregs.regs\[22\]\[25\]
+ cpuregs.regs\[23\]\[25\] _04275_ _04278_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__mux4_1
XANTENNA__09385__C1 _04049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12021_ _06114_ cpuregs.regs\[22\]\[3\] _06460_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__mux2_1
XANTENNA__11657__A _06215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15129__A _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13720__A2 _04979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14033__A _06053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10534__A2 _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15458__C1 _02004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16659__S _03062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13872__A _06072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16760_ _03121_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__clkbuf_1
X_13972_ _07747_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14681__B1 _07986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_171_Left_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15711_ timer\[13\] timer\[14\] _02516_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__or3_1
X_12923_ _06969_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09783__S0 _04282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16691_ _06957_ cpuregs.regs\[19\]\[7\] _03076_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08685__B net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13083__S _07057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18430_ clknet_leaf_183_clk _01495_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10393__S1 _04124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15642_ is_lb_lh_lw_lbu_lhu _03270_ _03396_ is_sb_sh_sw VGND VGND VPWR VPWR _02469_
+ sky130_fd_sc_hd__a22o_1
X_12854_ _06926_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18361_ clknet_leaf_187_clk _01426_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11805_ _06084_ _06346_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__nand2_2
XANTENNA_output100_A net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15573_ cpuregs.regs\[20\]\[28\] cpuregs.regs\[21\]\[28\] cpuregs.regs\[22\]\[28\]
+ cpuregs.regs\[23\]\[28\] _01918_ _01919_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__mux4_1
X_12785_ _06889_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11798__A1 _06072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10145__S1 _04759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17312_ clknet_leaf_175_clk _00486_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15608__S0 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14524_ _07943_ _08162_ VGND VGND VPWR VPWR _08185_ sky130_fd_sc_hd__nand2_1
X_11736_ reg_out\[24\] alu_out_q\[24\] _06068_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__mux2_2
X_18292_ clknet_leaf_38_clk _01360_ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10470__A1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15084__S1 _03646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17243_ clknet_leaf_13_clk _00417_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10470__B2 _05175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14455_ _06860_ _08120_ VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__nor2_2
XFILLER_0_142_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11667_ _06224_ cpuregs.regs\[10\]\[16\] _06176_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13406_ _04198_ _07269_ _07225_ VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__mux2_1
X_10618_ _05311_ _05320_ _05292_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__mux2_1
XANTENNA__11489__A_N net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17174_ clknet_leaf_126_clk _00348_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14386_ _08038_ _08054_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__or2_1
X_11598_ reg_pc\[8\] _06146_ reg_pc\[9\] VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_12_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16125_ net285 _05413_ _02771_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__mux2_1
X_10549_ _05224_ _05225_ _05252_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__or3_1
X_13337_ cpuregs.regs\[8\]\[0\] cpuregs.regs\[9\]\[0\] cpuregs.regs\[10\]\[0\] cpuregs.regs\[11\]\[0\]
+ _04579_ _04284_ VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16056_ _03402_ decoded_imm_j\[16\] _03403_ mem_rdata_q\[16\] VGND VGND VPWR VPWR
+ _02741_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13268_ _06955_ cpuregs.regs\[5\]\[6\] _07154_ VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15007_ _01862_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13258__S _07154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15039__A _05138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12162__S _06534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12219_ _06579_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13199_ _07124_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_166_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10081__S0 _04512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13782__A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15473__S _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16661__A1 _06296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16958_ clknet_leaf_18_clk _00132_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_127_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08876__A _03640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14672__B1 _08055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10289__A1 _04206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11486__B1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15909_ is_alu_reg_imm _02611_ _02620_ _02647_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_144_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16889_ clknet_leaf_33_clk _00059_ VGND VGND VPWR VPWR mem_rdata_q\[8\] sky130_fd_sc_hd__dfxtp_1
X_09430_ _03680_ _04160_ _04163_ _03226_ _04049_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18628_ clknet_leaf_184_clk _01688_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11238__B1 _05871_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09361_ _04053_ _04094_ _04095_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__a21o_1
XANTENNA__13778__A2 _05107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18559_ clknet_leaf_131_clk _01624_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09203__C _03878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11789__A1 alu_out_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09292_ _04010_ _04020_ _04028_ _03303_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_12 _02397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_23 _04271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09500__A _04084_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10461__A1 _04053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 _05110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_45 _06165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09829__S1 _04218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 mem_rdata_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_78 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09603__B1 _04237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_89 net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13957__A _03304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09646__S _04321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15152__B2 _02004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput130 net130 VGND VGND VPWR VPWR cpi_rs2[9] sky130_fd_sc_hd__buf_1
Xoutput141 net141 VGND VGND VPWR VPWR eoi[19] sky130_fd_sc_hd__buf_1
XFILLER_0_101_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput152 net152 VGND VGND VPWR VPWR eoi[29] sky130_fd_sc_hd__buf_1
XANTENNA__13168__S _07104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput163 net163 VGND VGND VPWR VPWR mem_addr[10] sky130_fd_sc_hd__clkbuf_1
Xoutput174 net174 VGND VGND VPWR VPWR mem_addr[21] sky130_fd_sc_hd__buf_1
XFILLER_0_100_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput185 net185 VGND VGND VPWR VPWR mem_addr[31] sky130_fd_sc_hd__buf_1
Xoutput196 net196 VGND VGND VPWR VPWR mem_la_addr[12] sky130_fd_sc_hd__buf_1
XANTENNA__08489__C _03272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10072__S0 _04512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16479__S _02968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08590__B1 instr_waitirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09628_ reg_pc\[7\] decoded_imm\[7\] VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09559_ _04055_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__buf_6
XFILLER_0_66_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12570_ cpuregs.regs\[2\]\[19\] _06573_ _06763_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__mux2_1
XANTENNA__08645__A1 irq_mask\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09264__B1_N _03763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11521_ _06090_ _06091_ _06093_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08771__B_N net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10556__A _05259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11452_ _06041_ irq_pending\[14\] _06044_ net6 VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__a31o_1
X_14240_ reg_pc\[13\] _07926_ _07934_ _07935_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__a22o_1
XANTENNA__15391__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10275__B decoded_imm\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14970__B _04448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10403_ _03680_ _05086_ _04752_ _05087_ _05110_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14171_ _07884_ _07815_ _07885_ VGND VGND VPWR VPWR _07886_ sky130_fd_sc_hd__and3b_1
XFILLER_0_21_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11383_ _03781_ _03789_ _03768_ _03736_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__or4_1
XANTENNA__15785__C _07984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10334_ net85 VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__clkbuf_4
X_13122_ _06945_ cpuregs.regs\[4\]\[1\] _07082_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17930_ clknet_leaf_62_clk _08370_ VGND VGND VPWR VPWR reg_out\[10\] sky130_fd_sc_hd__dfxtp_1
X_13053_ _07047_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11387__A _03228_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14497__A3 _07992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10265_ _04068_ _04976_ _04080_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__a21o_1
XANTENNA__10291__A _04223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12004_ _06454_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09373__A2 _04014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17861_ clknet_leaf_93_clk _01030_ VGND VGND VPWR VPWR count_cycle\[6\] sky130_fd_sc_hd__dfxtp_1
X_10196_ irq_mask\[22\] _04308_ timer\[22\] instr_timer _04026_ VGND VGND VPWR VPWR
+ _04910_ sky130_fd_sc_hd__a221o_1
XANTENNA__16389__S _02918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output148_A net148 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16812_ _03148_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17792_ clknet_leaf_82_clk _00961_ VGND VGND VPWR VPWR count_instr\[63\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12710__S _06847_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08696__A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11468__B1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16743_ reg_sh\[0\] _03314_ _01929_ _03638_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13955_ _07714_ _07735_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_89_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11326__S _03219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12906_ _06957_ cpuregs.regs\[31\]\[7\] _06943_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16674_ _03074_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__clkbuf_1
X_13886_ _07675_ _07687_ VGND VGND VPWR VPWR _07688_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18413_ clknet_leaf_161_clk _01478_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__14957__A1 net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ cpuregs.regs\[28\]\[31\] cpuregs.regs\[29\]\[31\] cpuregs.regs\[30\]\[31\]
+ cpuregs.regs\[31\]\[31\] _03640_ _03642_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_122_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12837_ _06175_ cpuregs.regs\[6\]\[10\] _06917_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12968__A0 _06999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10118__S1 _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18344_ clknet_leaf_36_clk _01412_ VGND VGND VPWR VPWR mem_16bit_buffer\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15556_ cpuregs.regs\[28\]\[27\] cpuregs.regs\[29\]\[27\] cpuregs.regs\[30\]\[27\]
+ cpuregs.regs\[31\]\[27\] _01996_ _01997_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12768_ cpuregs.regs\[9\]\[10\] _06554_ _06880_ VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12665__B _06082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14507_ _08166_ _08167_ VGND VGND VPWR VPWR _08169_ sky130_fd_sc_hd__or2_1
XANTENNA__15041__B _01863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11719_ reg_out\[22\] alu_out_q\[22\] _06068_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__mux2_1
X_18275_ clknet_leaf_23_clk _01345_ VGND VGND VPWR VPWR compressed_instr sky130_fd_sc_hd__dfxtp_1
XANTENNA__16852__S _03163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15487_ cpuregs.regs\[24\]\[23\] cpuregs.regs\[25\]\[23\] cpuregs.regs\[26\]\[23\]
+ cpuregs.regs\[27\]\[23\] _03645_ _01991_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__mux4_1
XANTENNA__11061__S _05322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12699_ _06216_ cpuregs.regs\[12\]\[15\] _06836_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__mux2_1
XANTENNA__08581__D _03359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17226_ clknet_leaf_147_clk _00400_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14438_ decoded_imm_j\[11\] _07930_ VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__or2_1
Xinput10 irq[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 irq[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
XFILLER_0_141_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput32 irq[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xinput43 mem_rdata[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
XANTENNA__13393__A0 _04160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput54 mem_rdata[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_2
X_17157_ clknet_leaf_148_clk _00331_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput65 mem_ready VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14369_ _03368_ _08041_ VGND VGND VPWR VPWR _08042_ sky130_fd_sc_hd__nand2_1
XANTENNA__09061__A1 mem_rdata_q\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09466__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16108_ _03286_ _03220_ _01821_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__and3_1
X_17088_ clknet_leaf_186_clk _00262_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13145__A0 _06968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11297__A _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08930_ _03683_ _03688_ _03693_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__a21o_1
X_16039_ decoded_imm\[8\] _02711_ _02731_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14893__B1 _05200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09990__A _04668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10054__S0 _04232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08861_ _03626_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__inv_2
XANTENNA__16299__S _02870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11171__A2 _04710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16634__A1 _06192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16095__C1 _06026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08792_ net103 net71 VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__and2b_1
XANTENNA__13448__A1 _03524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12620__S _06799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09413_ count_instr\[2\] _04145_ _04009_ _04146_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__a211o_1
XANTENNA__15296__S1 _02000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09344_ _04075_ _04076_ _04078_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10434__A1 _04168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09275_ _04011_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12067__S _06482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15373__A1 decoded_imm\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14790__B _08350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13687__A _03575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14884__B1 _01714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10050_ cpuregs.regs\[0\]\[18\] cpuregs.regs\[1\]\[18\] cpuregs.regs\[2\]\[18\] cpuregs.regs\[3\]\[18\]
+ _04057_ _04060_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__mux4_1
XANTENNA__16625__A1 _06156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10348__S1 _04208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09512__C1 _04150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13740_ _07568_ _07571_ _07580_ VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10952_ _05512_ _05600_ _05603_ _05345_ _05637_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10673__A1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15287__S1 _01971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13671_ _03584_ _05257_ VGND VGND VPWR VPWR _07517_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10883_ _05572_ _05511_ _05395_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__mux2_1
X_15410_ _02251_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15142__A _03647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12622_ _06184_ cpuregs.regs\[30\]\[11\] _06799_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08618__A1 mem_do_wdata VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16390_ _02924_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11622__A0 _06184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15341_ cpuregs.regs\[0\]\[15\] cpuregs.regs\[1\]\[15\] cpuregs.regs\[2\]\[15\] cpuregs.regs\[3\]\[15\]
+ _02085_ _02086_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12553_ _06764_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14981__A _04185_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09291__B2 _04024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18060_ clknet_leaf_73_clk _01165_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_124_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11504_ _06077_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__buf_2
X_15272_ cpuregs.regs\[8\]\[11\] cpuregs.regs\[9\]\[11\] cpuregs.regs\[10\]\[11\]
+ cpuregs.regs\[11\]\[11\] _01973_ _01974_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12484_ _06727_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17011_ clknet_leaf_20_clk _00185_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14223_ reg_next_pc\[8\] _05858_ _07922_ _07923_ VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__o211a_2
XFILLER_0_62_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11435_ irq_mask\[7\] _06030_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__or2_1
XANTENNA__12705__S _06836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14154_ count_instr\[52\] count_instr\[51\] _07865_ _07868_ VGND VGND VPWR VPWR _07874_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_132_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11366_ _03783_ _03213_ _03876_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__and3_1
XANTENNA__13390__A3 _05259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15211__S1 _01977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10317_ _05025_ _05026_ _04077_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__mux2_1
X_13105_ _07074_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _07824_ _07825_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__nor2_1
X_11297_ _03841_ _05919_ _05920_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_163_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913_ clknet_leaf_84_clk _01082_ VGND VGND VPWR VPWR count_cycle\[58\] sky130_fd_sc_hd__dfxtp_1
X_10248_ net49 _04811_ _04667_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__a21o_2
XANTENNA__09977__S0 _04487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13036_ cpuregs.regs\[3\]\[25\] _06586_ _07032_ VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10587__S1 _05239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17844_ clknet_leaf_108_clk _01013_ VGND VGND VPWR VPWR reg_next_pc\[21\] sky130_fd_sc_hd__dfxtp_1
X_10179_ _04891_ _04892_ _04065_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__mux2_1
XANTENNA__14221__A _07901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10900__A2 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16092__A2 _03935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08857__C _03605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17775_ clknet_leaf_87_clk _00944_ VGND VGND VPWR VPWR count_instr\[46\] sky130_fd_sc_hd__dfxtp_1
X_14987_ irq_mask\[5\] _01864_ _01873_ _08335_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_141_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16726_ _03102_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__clkbuf_1
X_13938_ _07714_ _07723_ VGND VGND VPWR VPWR _07724_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15278__S1 _02070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16657_ cpuregs.regs\[1\]\[23\] _06280_ _03062_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13869_ cpuregs.regs\[0\]\[31\] VGND VGND VPWR VPWR _07674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15608_ cpuregs.regs\[24\]\[30\] cpuregs.regs\[25\]\[30\] cpuregs.regs\[26\]\[30\]
+ cpuregs.regs\[27\]\[30\] _02221_ _02222_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__mux4_1
XANTENNA__15052__A _03666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16588_ _03029_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18327_ clknet_leaf_19_clk _01395_ VGND VGND VPWR VPWR cpuregs.waddr\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09901__S0 _04329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15539_ _02367_ _02369_ _02372_ _02017_ _01968_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__a221o_1
XANTENNA__14891__A _03631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09060_ mem_16bit_buffer\[7\] _03821_ _03727_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__mux2_2
XFILLER_0_114_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18258_ clknet_leaf_24_clk _01329_ VGND VGND VPWR VPWR decoded_imm\[16\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_72_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17209_ clknet_leaf_14_clk _00383_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15450__S1 _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09034__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12615__S _06788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18189_ clknet_leaf_31_clk _01260_ VGND VGND VPWR VPWR instr_jalr sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15107__B2 _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15202__S1 _03642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09962_ reg_pc\[16\] decoded_imm\[16\] VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09924__S _04065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08913_ cpuregs.raddr2\[1\] cpuregs.raddr2\[0\] cpuregs.raddr2\[2\] VGND VGND VPWR
+ VPWR _03678_ sky130_fd_sc_hd__or3_1
X_09893_ cpuregs.regs\[0\]\[14\] cpuregs.regs\[1\]\[14\] cpuregs.regs\[2\]\[14\] cpuregs.regs\[3\]\[14\]
+ _04290_ _04276_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__mux4_1
XANTENNA__11144__A2 _05254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13446__S _07225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08844_ net67 _03609_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1014 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08775_ _03531_ net92 _03540_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16757__S _03116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14397__A2 _07994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15897__A _03304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09327_ cpuregs.regs\[24\]\[1\] cpuregs.regs\[25\]\[1\] cpuregs.regs\[26\]\[1\] cpuregs.regs\[27\]\[1\]
+ _04057_ _04060_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09895__A _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15346__A1 _02012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09258_ _03775_ _03995_ _03763_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09189_ _03785_ _03934_ _03937_ _03932_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11220_ _05834_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__buf_2
XFILLER_0_31_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11151_ _05810_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__buf_2
XFILLER_0_101_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10591__A0 _03524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10102_ reg_pc\[18\] decoded_imm\[18\] _04783_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__and3_1
XANTENNA__09834__S _04077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11082_ _05758_ VGND VGND VPWR VPWR alu_out\[27\] sky130_fd_sc_hd__clkbuf_1
X_10033_ _04714_ _04718_ _04749_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__a21oi_1
X_14910_ _01829_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15137__A _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15890_ is_lb_lh_lw_lbu_lhu _02611_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ _01780_ _01781_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14976__A _04101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16667__S _03062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13880__A _07675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ clknet_leaf_109_clk _00729_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_14772_ _01734_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__clkbuf_1
X_11984_ _06240_ cpuregs.regs\[21\]\[18\] _06435_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14695__B _07815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16511_ _02988_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__clkbuf_1
X_13723_ _04959_ _07565_ _07224_ VGND VGND VPWR VPWR _07566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10935_ _05244_ _05621_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__nand2_1
X_17491_ clknet_leaf_156_clk _00660_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08934__S1 _03659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13091__S _07057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16442_ _06980_ cpuregs.regs\[29\]\[18\] _02943_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13654_ _07499_ _07500_ VGND VGND VPWR VPWR _07501_ sky130_fd_sc_hd__nand2_1
XANTENNA__16782__A0 _06565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14388__A2 _07905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10866_ _05226_ _05227_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12399__A1 _06540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12605_ _06114_ cpuregs.regs\[30\]\[3\] _06788_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16373_ _02915_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09264__A1 _03737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13585_ _07435_ _07436_ VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10797_ _03512_ _05468_ _03511_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_156_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18112_ clknet_leaf_81_clk _01216_ VGND VGND VPWR VPWR timer\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_639 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11071__A1 _05277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15324_ cpuregs.regs\[20\]\[14\] cpuregs.regs\[21\]\[14\] cpuregs.regs\[22\]\[14\]
+ cpuregs.regs\[23\]\[14\] _01976_ _01977_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__mux4_1
XFILLER_0_109_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15337__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12536_ _06755_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18043_ clknet_leaf_82_clk _00020_ VGND VGND VPWR VPWR irq_pending\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15432__S1 _01977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15255_ cpuregs.regs\[28\]\[10\] cpuregs.regs\[29\]\[10\] cpuregs.regs\[30\]\[10\]
+ cpuregs.regs\[31\]\[10\] _02022_ _02023_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__mux4_1
X_12467_ _06718_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12435__S _06700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output92_A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12813__B_N _06082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14206_ _03294_ VGND VGND VPWR VPWR _07912_ sky130_fd_sc_hd__clkbuf_4
X_11418_ _06003_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__inv_2
X_15186_ decoded_imm\[6\] _02009_ _01963_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_134_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12398_ _06681_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14137_ count_instr\[47\] count_instr\[46\] _07859_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__and3_1
X_11349_ _03891_ _03767_ _03770_ _03736_ _05963_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14068_ count_instr\[26\] _07811_ _07813_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__o21a_1
XANTENNA__09724__C1 _04150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13266__S _07154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13019_ cpuregs.regs\[3\]\[17\] _06569_ _07021_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__mux2_1
XANTENNA__15047__A _03664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17827_ clknet_leaf_57_clk _00996_ VGND VGND VPWR VPWR reg_next_pc\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12087__A0 _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08560_ _03335_ _03336_ _03337_ _03338_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__or4_1
X_17758_ clknet_leaf_89_clk _00927_ VGND VGND VPWR VPWR count_instr\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08884__A _03640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08491_ cpu_state\[6\] cpu_state\[5\] VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__or2_2
XFILLER_0_7_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16709_ _03093_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08925__S1 _03659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17689_ clknet_leaf_108_clk _00858_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15576__A1 _02111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15120__S0 _01973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09112_ _03852_ _03861_ _03871_ _03855_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10270__C1 _04149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13339__B1 _04296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09043_ net43 mem_rdata_q\[19\] _03730_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15423__S1 _03642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12345__S _06652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12562__A1 _06565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13965__A _07737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09945_ _04665_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__buf_2
XANTENNA__15500__A1 _01982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13511__A0 _04342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13176__S _07104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09876_ _04597_ _04598_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__nand2_1
XANTENNA__10325__B1 _00073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16056__A2 decoded_imm_j\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08827_ net120 net88 VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__and2b_1
XANTENNA__10876__A1 _05219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10420__S0 _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16487__S _02968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08758_ net94 VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11825__A0 _06166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ net116 net84 VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__nor2_1
XANTENNA__09494__A1 _04215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10720_ _05400_ _05418_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13578__A0 _04611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10651_ _05349_ _05352_ _05287_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__mux2_1
XANTENNA__09246__B2 _03888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10582_ _05284_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__inv_2
X_13370_ _05258_ VGND VGND VPWR VPWR _07236_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09341__S1 _04074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10487__S0 _04325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10800__A1 _05323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15414__S1 _03647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12321_ cpuregs.waddr\[0\] cpuregs.waddr\[1\] VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__or2b_2
XANTENNA__12255__S _06604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18731__A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15040_ irq_mask\[29\] _01865_ _01902_ _01891_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_181_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12252_ cpuregs.waddr\[2\] cpuregs.waddr\[4\] cpuregs.waddr\[3\] _06601_ VGND VGND
+ VPWR VPWR _06602_ sky130_fd_sc_hd__and4b_1
XFILLER_0_32_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13750__A0 _05044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09954__C1 _04674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13875__A _03292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11203_ _05831_ _05835_ _05840_ _05843_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__and4_1
X_12183_ _06533_ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10564__A0 _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15178__S0 _02030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09564__S _04223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13594__B decoded_imm\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11134_ _05456_ _05700_ _05802_ _05806_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_112_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16991_ clknet_leaf_181_clk _00165_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08688__B net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12305__A1 _06584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13502__B1 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18730_ net125 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_1
X_11065_ _05727_ _05735_ _05742_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__or3_1
X_15942_ _02666_ mem_rdata_q\[26\] mem_rdata_q\[27\] _02658_ VGND VGND VPWR VPWR _02667_
+ sky130_fd_sc_hd__and4bb_4
X_10016_ _04053_ _04734_ _04095_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output130_A net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15873_ instr_bgeu _02618_ _02622_ _02627_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__a22o_1
XANTENNA__16397__S _02918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output228_A net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14824_ count_cycle\[43\] _01768_ _01717_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__a21oi_1
X_17612_ clknet_leaf_160_clk _00781_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_18592_ clknet_leaf_182_clk _01657_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17543_ clknet_leaf_178_clk _00712_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14755_ _06053_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08907__S1 _03671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11967_ _06423_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_158_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13706_ net82 decoded_imm\[23\] VGND VGND VPWR VPWR _07549_ sky130_fd_sc_hd__nor2_1
X_10918_ _03485_ _05220_ _05249_ _05603_ _05605_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__a221o_1
XANTENNA__09312__B cpu_state\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17474_ clknet_leaf_1_clk _00643_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14686_ _08330_ _08331_ _08332_ VGND VGND VPWR VPWR _08333_ sky130_fd_sc_hd__o21a_1
X_11898_ _06386_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_168_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15022__A3 _04842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_134_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16425_ _02931_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__buf_6
X_13637_ _07274_ _07484_ _07191_ VGND VGND VPWR VPWR _07485_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09237__A1 _03977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10849_ _03498_ _05398_ _05367_ _03497_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__o22a_1
XFILLER_0_157_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_171_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16356_ _02906_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13568_ _07406_ _07409_ _07407_ VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_136_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08996__A0 mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11595__A2 _03323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15307_ cpuregs.regs\[28\]\[13\] cpuregs.regs\[29\]\[13\] cpuregs.regs\[30\]\[13\]
+ cpuregs.regs\[31\]\[13\] _01990_ _01992_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12519_ _06745_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16287_ _02869_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12165__S _06534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13499_ _04419_ _05260_ _07316_ _07279_ VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_149_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18026_ clknet_leaf_65_clk _00002_ VGND VGND VPWR VPWR irq_pending\[10\] sky130_fd_sc_hd__dfxtp_1
X_15238_ _02082_ _02083_ _02084_ _02087_ _01982_ _02088_ VGND VGND VPWR VPWR _02089_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_132_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15169_ _03647_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09960__A2 decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08598__B irq_state\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__15494__B1 _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09730_ net50 _04030_ _04034_ net64 _04423_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__o221a_1
XFILLER_0_66_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16038__A2 decoded_imm_j\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09661_ irq_pending\[7\] _04049_ _04389_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_2_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08612_ is_lui_auipc_jal VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__clkbuf_4
X_09592_ _04318_ _04319_ _04321_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__mux2_1
XANTENNA__15341__S0 _02085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11807__A0 _06078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08543_ irq_mask\[5\] irq_pending\[5\] VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__and2b_2
XFILLER_0_49_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13025__A _07009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15549__A1 _02382_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12480__A0 _06166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16746__B1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08474_ instr_lbu instr_lb VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__or2_1
XANTENNA__09571__S1 _04219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16336__A _02895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15240__A _01984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13679__B decoded_imm\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11130__S1 _05286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12075__S _06482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09026_ _03787_ _03749_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__nor2_1
XANTENNA__11199__B _05840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12803__S _06891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09928_ _04647_ _04648_ _04121_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__mux2_1
X_09859_ _04206_ _04581_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__nand2_1
XANTENNA__15788__A1 latched_store VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15332__S0 _02074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12870_ _06304_ cpuregs.regs\[6\]\[26\] _06928_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_102 _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_113 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11821_ _06150_ cpuregs.regs\[11\]\[7\] _06348_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__18148__D alu_out\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_124 net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_135 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18726__A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11154__S _04745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_146 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14540_ _08177_ _08188_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__and2_1
X_11752_ reg_pc\[26\] _06291_ _06299_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__o21a_1
XANTENNA__09562__S1 _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10703_ _05402_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09219__A1 _03864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14471_ _07934_ _08119_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11683_ _06226_ reg_next_pc\[18\] _06236_ _06238_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__a211o_2
X_16210_ _03187_ _03198_ _03215_ _03217_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_153_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _07281_ _04241_ _07282_ reg_pc\[4\] _07284_ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__a221o_1
XFILLER_0_165_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11026__B2 _05254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10634_ _05333_ _05335_ _05295_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__mux2_1
X_17190_ clknet_leaf_137_clk _00364_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11577__A2 _03349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16141_ _02788_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__clkbuf_1
X_13353_ cpu_state\[4\] _03274_ VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__or2_1
X_10565_ net81 _04945_ _05236_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12304_ _06630_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_114_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16072_ decoded_imm\[22\] _02750_ _02746_ mem_rdata_q\[22\] _02749_ VGND VGND VPWR
+ VPWR _01335_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13284_ _07169_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__clkbuf_1
X_10496_ _05200_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__inv_2
XANTENNA__13723__A0 _04959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output178_A net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15023_ irq_mask\[21\] _01863_ _01714_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12235_ _06311_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__buf_2
XANTENNA__10537__A0 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08699__A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09942__A2 _04145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12166_ _06543_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14279__A1 reg_pc\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15476__B1 _02197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11117_ _05790_ _05764_ _05729_ _05702_ _05286_ _05277_ VGND VGND VPWR VPWR _05791_
+ sky130_fd_sc_hd__mux4_1
X_12097_ _06150_ cpuregs.regs\[23\]\[7\] _06496_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__mux2_1
XANTENNA__15571__S0 _02111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16974_ clknet_leaf_101_clk _00148_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11048_ _05726_ VGND VGND VPWR VPWR alu_out\[25\] sky130_fd_sc_hd__clkbuf_1
X_15925_ instr_xor _02617_ _02623_ _02653_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__a22o_1
XANTENNA__15228__B1 _01963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 irq[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12949__A _06265_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13345__A2_N _07208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15856_ _03239_ _02610_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__nor2_2
XANTENNA__15323__S0 _01973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18644_ clknet_leaf_164_clk _01704_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15779__B2 _06186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14807_ count_cycle\[37\] _01756_ _01758_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__o21a_1
XANTENNA__14987__C1 _08335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15787_ _03384_ _02574_ _02576_ _03226_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__a211o_1
XANTENNA__09458__A1 _04010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18575_ clknet_leaf_20_clk _01640_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_12999_ _07018_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10068__A2 decoded_imm\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12462__A0 _06078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14738_ count_cycle\[16\] _08365_ _08367_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17526_ clknet_leaf_97_clk _00695_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_173_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11999__S _06446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17457_ clknet_leaf_132_clk _00626_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14669_ _08232_ _07969_ VGND VGND VPWR VPWR _08317_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16408_ _02934_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_41_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17388_ clknet_leaf_116_clk _00557_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10916__B _05398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08969__A0 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16339_ _06945_ cpuregs.regs\[16\]\[1\] _02896_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18009_ clknet_leaf_78_clk _01146_ VGND VGND VPWR VPWR irq_mask\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08402__A latched_branch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09713_ cpuregs.regs\[24\]\[9\] cpuregs.regs\[25\]\[9\] cpuregs.regs\[26\]\[9\] cpuregs.regs\[27\]\[9\]
+ _04217_ _04219_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__mux4_1
XANTENNA__09932__S _04121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15235__A _01919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09644_ cpuregs.regs\[28\]\[7\] cpuregs.regs\[29\]\[7\] cpuregs.regs\[30\]\[7\] cpuregs.regs\[31\]\[7\]
+ _04325_ _04277_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09575_ _04272_ _04301_ _04305_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_167_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16765__S _03116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _03305_ _03246_ _03247_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_26_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16719__A0 _06984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13650__C1 _07283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15617__S1 _02047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16195__A1 net257 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08457_ reg_next_pc\[0\] _03199_ net66 VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__and3_1
XANTENNA__08791__B net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11008__A1 _04913_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10231__A2 _04923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10350_ _05057_ _05058_ _04211_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09009_ net51 mem_rdata_q\[26\] _03729_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__mux2_1
X_10281_ count_instr\[25\] _04012_ count_cycle\[25\] _04165_ _04991_ VGND VGND VPWR
+ VPWR _04992_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10519__B1 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12533__S _06752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12020_ _06463_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10534__A3 _04198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15844__S _03635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15553__S0 _01973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13872__B _03298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13971_ _07737_ _07746_ VGND VGND VPWR VPWR _07747_ sky130_fd_sc_hd__and2_1
XANTENNA__09688__B2 _04023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14681__A1 _07971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15710_ timer\[13\] _02516_ timer\[14\] VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15145__A _03647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12922_ _06968_ cpuregs.regs\[31\]\[12\] _06964_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__mux2_1
X_16690_ _03083_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09783__S1 _04285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15641_ _07992_ _02466_ _02467_ _03410_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__a211oi_1
X_12853_ _06240_ cpuregs.regs\[6\]\[18\] _06917_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__mux2_1
XANTENNA__15630__A0 net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14433__B2 _08033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11247__A1 _05829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11804_ _06345_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__buf_4
X_18360_ clknet_leaf_10_clk _01425_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_15572_ cpuregs.regs\[16\]\[28\] cpuregs.regs\[17\]\[28\] cpuregs.regs\[18\]\[28\]
+ cpuregs.regs\[19\]\[28\] _01918_ _01919_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__mux4_1
X_12784_ cpuregs.regs\[9\]\[18\] _06571_ _06880_ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17311_ clknet_leaf_181_clk _00485_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15608__S1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14523_ _07898_ _07943_ _07997_ _08183_ VGND VGND VPWR VPWR _08184_ sky130_fd_sc_hd__a22o_1
X_11735_ _06283_ _06118_ _06284_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__and3b_1
X_18291_ clknet_leaf_5_clk _01359_ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17242_ clknet_leaf_186_clk _00416_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10470__A2 _05174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14454_ _03364_ _07986_ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__nand2_2
XFILLER_0_126_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11666_ _06223_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__buf_2
XFILLER_0_126_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10736__B _05259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13405_ _03276_ _07262_ _07263_ _07268_ VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10617_ _05314_ _05319_ _05295_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17173_ clknet_leaf_116_clk _00347_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_14385_ _08024_ _08028_ _08040_ _08054_ VGND VGND VPWR VPWR _08057_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11597_ reg_pc\[9\] reg_pc\[8\] _06146_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16124_ _02779_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__clkbuf_1
X_13336_ cpuregs.regs\[12\]\[0\] cpuregs.regs\[13\]\[0\] cpuregs.regs\[14\]\[0\] cpuregs.regs\[15\]\[0\]
+ _04579_ _04284_ VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__mux4_1
XFILLER_0_150_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10548_ _05228_ _05245_ _05249_ _05251_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16055_ decoded_imm\[15\] _02720_ _02736_ _02740_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__o22a_1
XANTENNA__12443__S _06700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13267_ _07160_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__clkbuf_1
X_10479_ cpuregs.regs\[20\]\[31\] cpuregs.regs\[21\]\[31\] cpuregs.regs\[22\]\[31\]
+ cpuregs.regs\[23\]\[31\] _04291_ _04292_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__mux4_1
XFILLER_0_122_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15006_ irq_mask\[13\] _01880_ _01884_ _01876_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__a211o_1
XANTENNA__09318__A _04052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12218_ cpuregs.regs\[24\]\[21\] _06578_ _06576_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__mux2_1
XANTENNA__15039__B _01863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11183__A0 _04160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13198_ _06953_ cpuregs.regs\[8\]\[5\] _07118_ VGND VGND VPWR VPWR _07124_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_166_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10081__S1 _04513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12149_ _06077_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__buf_2
XANTENNA__10930__A0 _04744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15544__S0 _03640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09128__B1 _03885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13782__B decoded_imm\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16957_ clknet_leaf_187_clk _00131_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_127_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13274__S _07154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11583__A _06149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11486__A1 _06054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15908_ _02645_ _02646_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_144_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16888_ clknet_leaf_33_clk _00058_ VGND VGND VPWR VPWR mem_rdata_q\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_144_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09053__A _03810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18627_ clknet_leaf_174_clk _01687_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10199__A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16585__S _03026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15839_ _03878_ _03885_ _03895_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__and3b_1
XFILLER_0_149_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09988__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09360_ _00073_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__clkbuf_8
X_18558_ clknet_leaf_182_clk _01623_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12986__A1 _06536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17509_ clknet_leaf_1_clk _00678_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09291_ irq_mask\[0\] _04022_ timer\[0\] _04024_ _04027_ VGND VGND VPWR VPWR _04028_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__16177__A1 net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18489_ clknet_leaf_1_clk _01554_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_13 _02412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14188__B1 _03240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_24 _04289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 _05313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_46 _06752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 reg_next_pc\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_68 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09603__A1 _04328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15688__B1 _02476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12353__S _06652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput120 net120 VGND VGND VPWR VPWR cpi_rs2[29] sky130_fd_sc_hd__buf_1
XANTENNA__10662__A _05323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput131 net131 VGND VGND VPWR VPWR eoi[0] sky130_fd_sc_hd__buf_1
Xoutput142 net142 VGND VGND VPWR VPWR eoi[1] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15850__B_N decoder_trigger VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput153 net153 VGND VGND VPWR VPWR eoi[2] sky130_fd_sc_hd__buf_1
XANTENNA__11477__B _03428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput164 net164 VGND VGND VPWR VPWR mem_addr[11] sky130_fd_sc_hd__clkbuf_1
XANTENNA__11174__B1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput175 net175 VGND VGND VPWR VPWR mem_addr[22] sky130_fd_sc_hd__clkbuf_1
Xoutput186 net186 VGND VGND VPWR VPWR mem_addr[3] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput197 net197 VGND VGND VPWR VPWR mem_la_addr[13] sky130_fd_sc_hd__buf_1
XANTENNA__16101__A1 _03635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10072__S1 _04513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09119__A0 mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08590__A1 decoder_trigger VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13184__S _07081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12674__A0 _06114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09627_ reg_pc\[7\] decoded_imm\[7\] VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15612__B1 _02441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09558_ _04214_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08509_ cpu_state\[1\] VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08645__A2 _03412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09489_ cpuregs.regs\[16\]\[4\] cpuregs.regs\[17\]\[4\] cpuregs.regs\[18\]\[4\] cpuregs.regs\[19\]\[4\]
+ _04217_ _04219_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11520_ _06092_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11451_ irq_mask\[14\] _06042_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15391__A2 _01906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10048__S _04065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10402_ _04009_ _05089_ _05109_ _03301_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14170_ count_instr\[56\] _07881_ count_instr\[57\] VGND VGND VPWR VPWR _07885_ sky130_fd_sc_hd__a21o_1
X_11382_ _03816_ _03736_ _03853_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_12_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13359__S _07225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13121_ _07083_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__clkbuf_1
X_10333_ _05038_ _05039_ _05042_ _03302_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12263__S _06604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13052_ _06941_ cpuregs.regs\[7\]\[0\] _07046_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__mux2_1
XANTENNA__11387__B _03979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10264_ _04974_ _04975_ _04077_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15574__S _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12003_ _06312_ cpuregs.regs\[21\]\[27\] _06446_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__mux2_1
XANTENNA__13883__A _07675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10195_ _04908_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__inv_2
XANTENNA__15526__S0 _02074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17860_ clknet_leaf_93_clk _01029_ VGND VGND VPWR VPWR count_cycle\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08977__A _03213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14103__B1 _07675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16811_ _06594_ cpuregs.regs\[13\]\[29\] _03138_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__mux2_1
XANTENNA__15300__C1 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17791_ clknet_leaf_82_clk _00960_ VGND VGND VPWR VPWR count_instr\[62\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13094__S _07068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13954_ _03343_ _07727_ _07728_ net146 VGND VGND VPWR VPWR _07735_ sky130_fd_sc_hd__a22o_1
X_16742_ _03110_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_161_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12905_ _06149_ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__buf_2
XANTENNA_output210_A net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16673_ cpuregs.regs\[1\]\[31\] _06342_ _03039_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__mux2_1
X_13885_ _03326_ _07678_ _07682_ net153 VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18412_ clknet_leaf_109_clk _01477_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ cpuregs.regs\[24\]\[31\] cpuregs.regs\[25\]\[31\] cpuregs.regs\[26\]\[31\]
+ cpuregs.regs\[27\]\[31\] _03640_ _03642_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__mux4_1
X_12836_ _06905_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _02384_ _02385_ _02386_ _02387_ _02111_ _02004_ VGND VGND VPWR VPWR _02388_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__16159__A1 net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18343_ clknet_leaf_37_clk _01411_ VGND VGND VPWR VPWR mem_16bit_buffer\[14\] sky130_fd_sc_hd__dfxtp_1
X_12767_ _06868_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11025__A2_N _05221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14506_ _08166_ _08167_ VGND VGND VPWR VPWR _08168_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11718_ _06268_ _06269_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18274_ clknet_leaf_25_clk _00033_ VGND VGND VPWR VPWR is_lui_auipc_jal sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15486_ cpuregs.regs\[28\]\[23\] cpuregs.regs\[29\]\[23\] cpuregs.regs\[30\]\[23\]
+ cpuregs.regs\[31\]\[23\] _03645_ _01991_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12698_ _06841_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17225_ clknet_leaf_135_clk _00399_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14437_ decoded_imm_j\[11\] _07930_ VGND VGND VPWR VPWR _08104_ sky130_fd_sc_hd__nand2_1
X_11649_ _06208_ cpuregs.regs\[10\]\[14\] _06176_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput11 irq[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput22 irq[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
XFILLER_0_142_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput33 mem_rdata[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11944__B_N cpuregs.waddr\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput44 mem_rdata[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17156_ clknet_leaf_143_clk _00330_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput55 mem_rdata[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_1
X_14368_ _08024_ _08028_ _08040_ VGND VGND VPWR VPWR _08041_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput66 resetn VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_168_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16107_ _03309_ _03255_ _02618_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13319_ _07187_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__clkbuf_1
X_17087_ clknet_leaf_181_clk _00261_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10482__A _04289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14299_ irq_pending\[24\] irq_pending\[25\] irq_pending\[26\] irq_pending\[27\] VGND
+ VGND VPWR VPWR _07976_ sky130_fd_sc_hd__or4_1
XFILLER_0_110_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16038_ _02715_ decoded_imm_j\[8\] _02726_ mem_rdata_q\[28\] _02634_ VGND VGND VPWR
+ VPWR _02731_ sky130_fd_sc_hd__a221o_1
XANTENNA__11156__A0 _05254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13696__A2 _04941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09444__S0 _04084_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15484__S _03653_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14893__B2 _03387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08860_ is_slti_blt_slt _03431_ _03625_ _03430_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__a211o_1
XANTENNA__10054__S1 _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15517__S0 _02030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08791_ net102 net70 VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__and2b_1
XANTENNA__13448__A2 decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17989_ clknet_leaf_105_clk _01126_ VGND VGND VPWR VPWR irq_mask\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15842__B1 _06016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10421__S _04121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_185_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_185_clk sky130_fd_sc_hd__clkbuf_2
X_09412_ count_instr\[34\] _04015_ _04017_ count_cycle\[34\] VGND VGND VPWR VPWR _04146_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09343_ _04077_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__buf_6
XFILLER_0_48_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10434__A2 _05139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09274_ instr_rdinstr VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15358__C1 _02006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13968__A _07737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15373__A2 _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14581__B1 _07956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10198__A1 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12083__S _06496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11147__B1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14799__A _03304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08989_ _03738_ _03750_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__nor2_1
XANTENNA__10370__B2 _05078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10951_ _03482_ _05215_ _05334_ _05254_ _05636_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_176_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_176_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13670_ _07514_ _07515_ VGND VGND VPWR VPWR _07516_ sky130_fd_sc_hd__and2b_1
XANTENNA__10673__A2 _04419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10882_ _05571_ _05543_ _05240_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12621_ _06800_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08618__A2 _03218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11162__S _04668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15340_ cpuregs.regs\[4\]\[15\] cpuregs.regs\[5\]\[15\] cpuregs.regs\[6\]\[15\] cpuregs.regs\[7\]\[15\]
+ _01976_ _01977_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__mux4_1
X_12552_ cpuregs.regs\[2\]\[10\] _06554_ _06763_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09291__A2 _04022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11503_ _06066_ _06070_ _06073_ _06076_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__a211o_2
XFILLER_0_47_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13878__A _07681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15271_ cpuregs.regs\[12\]\[11\] cpuregs.regs\[13\]\[11\] cpuregs.regs\[14\]\[11\]
+ cpuregs.regs\[15\]\[11\] _01970_ _01971_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__mux4_1
XFILLER_0_109_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12483_ _06175_ cpuregs.regs\[28\]\[10\] _06726_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__mux2_1
X_17010_ clknet_leaf_111_clk _00184_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13375__A1 _03276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14222_ _05856_ _06153_ VGND VGND VPWR VPWR _07923_ sky130_fd_sc_hd__or2_1
X_11434_ _06029_ irq_pending\[6\] _06034_ net29 VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09674__S0 _04056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13089__S _07057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14153_ _07872_ _07873_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__nor2_1
X_11365_ cpuregs.raddr2\[1\] _05974_ _05975_ _05978_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_100_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_100_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_132_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13104_ _06995_ cpuregs.regs\[7\]\[25\] _07068_ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__mux2_1
X_10316_ cpuregs.regs\[16\]\[26\] cpuregs.regs\[17\]\[26\] cpuregs.regs\[18\]\[26\]
+ cpuregs.regs\[19\]\[26\] _04123_ _04124_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__mux4_1
X_14084_ count_instr\[31\] _07821_ _07790_ VGND VGND VPWR VPWR _07825_ sky130_fd_sc_hd__o21ai_1
X_11296_ _05913_ _05915_ _05918_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output258_A net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17912_ clknet_leaf_84_clk _01081_ VGND VGND VPWR VPWR count_cycle\[57\] sky130_fd_sc_hd__dfxtp_1
X_13035_ _07037_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_163_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10247_ net83 VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09977__S1 _04469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14502__A decoded_imm_j\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17843_ clknet_leaf_60_clk _01012_ VGND VGND VPWR VPWR reg_next_pc\[20\] sky130_fd_sc_hd__dfxtp_1
X_10178_ cpuregs.regs\[16\]\[22\] cpuregs.regs\[17\]\[22\] cpuregs.regs\[18\]\[22\]
+ cpuregs.regs\[19\]\[22\] _04281_ _04470_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__mux4_1
XANTENNA__10900__A3 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17774_ clknet_leaf_95_clk _00943_ VGND VGND VPWR VPWR count_instr\[45\] sky130_fd_sc_hd__dfxtp_1
X_14986_ _01872_ _01869_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_141_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1007 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16725_ _06991_ cpuregs.regs\[19\]\[23\] _03098_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13937_ _03336_ _07704_ _07705_ net140 VGND VGND VPWR VPWR _07723_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_167_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_167_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13868_ _07673_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__clkbuf_1
X_16656_ _03065_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12819_ _06908_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__clkbuf_1
X_15607_ cpuregs.regs\[28\]\[30\] cpuregs.regs\[29\]\[30\] cpuregs.regs\[30\]\[30\]
+ cpuregs.regs\[31\]\[30\] _01908_ _01909_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12168__S _06534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13799_ _07620_ _07625_ _07633_ _07634_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__a211oi_2
X_16587_ _06989_ cpuregs.regs\[18\]\[22\] _03026_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__mux2_1
XANTENNA__16863__S _03174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18326_ clknet_leaf_39_clk _01394_ VGND VGND VPWR VPWR prefetched_high_word sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ _02370_ _02371_ _03653_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__mux2_1
XANTENNA__09282__A2 _04016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09901__S1 _04218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15469_ cpuregs.regs\[24\]\[22\] cpuregs.regs\[25\]\[22\] cpuregs.regs\[26\]\[22\]
+ cpuregs.regs\[27\]\[22\] _02069_ _02070_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18257_ clknet_leaf_31_clk _01328_ VGND VGND VPWR VPWR decoded_imm\[15\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_114_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17208_ clknet_leaf_176_clk _00382_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18188_ clknet_leaf_43_clk _01259_ VGND VGND VPWR VPWR instr_bgeu sky130_fd_sc_hd__dfxtp_1
Xmax_cap300 net301 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__buf_4
XFILLER_0_40_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17139_ clknet_leaf_109_clk _00313_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14315__B1 _03364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09961_ _04542_ _04599_ _04676_ _04678_ _04680_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__o311a_1
XANTENNA__15512__C1 _01969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11129__B1 _05357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08912_ _03639_ _03655_ _03676_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09892_ cpuregs.regs\[4\]\[14\] cpuregs.regs\[5\]\[14\] cpuregs.regs\[6\]\[14\] cpuregs.regs\[7\]\[14\]
+ _04290_ _04276_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08843_ net99 VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08410__A net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08774_ _03534_ _03538_ _03539_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_158_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_158_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15579__C1 _02004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09326_ cpuregs.regs\[28\]\[1\] cpuregs.regs\[29\]\[1\] cpuregs.regs\[30\]\[1\] cpuregs.regs\[31\]\[1\]
+ _04057_ _04060_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__mux4_1
XFILLER_0_164_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11604__A1 alu_out_q\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15897__B is_alu_reg_imm VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13698__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09257_ _03891_ _03862_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_895 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11710__S _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09188_ _03763_ _03928_ _03936_ _03869_ _03810_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09430__C1 _04049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11150_ _05286_ net107 _04745_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__mux2_1
XANTENNA__10591__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10101_ reg_pc\[16\] decoded_imm\[16\] _04715_ _04816_ VGND VGND VPWR VPWR _04817_
+ sky130_fd_sc_hd__a31o_1
X_11081_ _05744_ _05751_ _05757_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__or3_1
XANTENNA__12541__S _06752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09416__A _04149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10032_ _04714_ _04718_ _04749_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__and3_1
XANTENNA__14609__A1 _08071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18729__A net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14840_ count_cycle\[48\] _01777_ _01723_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_69_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14976__B _01865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ _01732_ _08350_ _01733_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__and3b_1
XANTENNA__13293__A0 _06980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10996__S _05323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_149_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_149_clk sky130_fd_sc_hd__clkbuf_2
X_11983_ _06443_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__clkbuf_1
X_13722_ _03276_ _07558_ _07559_ _07564_ VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__a31o_1
X_16510_ cpuregs.regs\[17\]\[18\] _06571_ _02979_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__mux2_1
X_10934_ instr_sll instr_slli _05226_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__o21a_2
XFILLER_0_169_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17490_ clknet_leaf_142_clk _00659_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16231__A0 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13653_ net79 decoded_imm\[20\] VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__or2_1
X_16441_ _02951_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10865_ _03495_ _05440_ _05357_ _03496_ _05555_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__o221a_1
XFILLER_0_128_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16683__S _03076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12604_ _06791_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__clkbuf_1
X_16372_ _06978_ cpuregs.regs\[16\]\[17\] _02907_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__mux2_1
X_13584_ _07432_ _07433_ _07434_ _03311_ VGND VGND VPWR VPWR _07436_ sky130_fd_sc_hd__a31o_1
XFILLER_0_171_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10796_ _05478_ _05487_ _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_30_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18111_ clknet_leaf_81_clk _01215_ VGND VGND VPWR VPWR timer\[26\] sky130_fd_sc_hd__dfxtp_1
X_15323_ cpuregs.regs\[0\]\[14\] cpuregs.regs\[1\]\[14\] cpuregs.regs\[2\]\[14\] cpuregs.regs\[3\]\[14\]
+ _01973_ _01974_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12535_ cpuregs.regs\[2\]\[2\] _06538_ _06752_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12716__S _06847_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18042_ clknet_leaf_78_clk _00019_ VGND VGND VPWR VPWR irq_pending\[26\] sky130_fd_sc_hd__dfxtp_1
X_15254_ cpuregs.regs\[24\]\[10\] cpuregs.regs\[25\]\[10\] cpuregs.regs\[26\]\[10\]
+ cpuregs.regs\[27\]\[10\] _01990_ _01992_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_476 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14545__B1 _07998_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12466_ _06105_ cpuregs.regs\[28\]\[2\] _06715_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09016__A2 _03763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14205_ reg_next_pc\[3\] _03189_ _07900_ _07910_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_117_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11417_ _03215_ _03879_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__nor2_1
X_15185_ _02019_ _02026_ _02027_ _02038_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_134_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12397_ cpuregs.regs\[27\]\[2\] _06538_ _06678_ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output85_A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14136_ _07860_ _07861_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__nor2_1
X_11348_ _03748_ _03790_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__nand2_1
X_14067_ count_instr\[26\] _07811_ _07775_ VGND VGND VPWR VPWR _07813_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15328__A _02066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12451__S _06700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11279_ reg_next_pc\[20\] reg_out\[20\] _05898_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__mux2_2
X_13018_ _07028_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16858__S _03163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17826_ clknet_leaf_21_clk _00995_ VGND VGND VPWR VPWR reg_next_pc\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09760__S _04121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17757_ clknet_leaf_82_clk _00926_ VGND VGND VPWR VPWR count_instr\[28\] sky130_fd_sc_hd__dfxtp_1
X_14969_ _08335_ _01861_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11591__A _06156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16708_ _06974_ cpuregs.regs\[19\]\[15\] _03087_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__mux2_1
X_08490_ _03226_ _03238_ _03251_ _03273_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17688_ clknet_leaf_115_clk _00857_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16639_ _03056_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15120__S1 _01974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16593__S _03026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13587__A1 _04611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_922 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09111_ _03865_ _03870_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18309_ clknet_leaf_35_clk _01377_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dfxtp_1
XANTENNA__16525__A1 _06586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10935__A _05244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09660__C1 _04388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12626__S _06799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13339__A1 _04054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09042_ mem_16bit_buffer\[4\] _03803_ _03728_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__mux2_2
XFILLER_0_60_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09638__S0 _04290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10146__S _04211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10022__B1 _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09935__S _04320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09944_ latched_is_lb latched_is_lh VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__or2_1
XANTENNA__12361__S _06652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08518__A1 _03298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13511__A1 _04611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11485__B _03428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09875_ reg_pc\[13\] decoded_imm\[13\] VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__or2_1
XANTENNA__10325__A1 _04068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ net119 VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09191__B2 _03888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10420__S1 _04478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16461__A0 _06999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08757_ net126 net94 VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13192__S _07118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11705__S _06258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08688_ net116 net84 VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__and2_1
XANTENNA__09494__A2 _04224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_963 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14775__B1 _01723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10650_ _05350_ _05351_ _05246_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09309_ reg_next_pc\[0\] decoded_imm\[0\] VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10581_ _05242_ _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__or2_1
XANTENNA__10487__S1 _04277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12320_ _06638_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14527__B1 decoded_imm_j\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12251_ _06600_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10056__S _04121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11202_ reg_next_pc\[6\] reg_out\[6\] _05834_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__mux2_1
XANTENNA__09954__B1 _04664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12182_ _06174_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10564__A1 _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15178__S1 _02031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11133_ _05591_ _05621_ _05690_ _05601_ _05805_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__a221oi_2
XANTENNA__12271__S _06604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16990_ clknet_leaf_170_clk _00164_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13502__A1 _07304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11064_ _05225_ _05740_ _05741_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__and3_1
X_15941_ mem_rdata_q\[28\] mem_rdata_q\[25\] _02632_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__or3_1
XANTENNA__11513__A0 _06078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13891__A _06053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10015_ _04732_ _04733_ _04064_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__mux2_1
X_15872_ _02612_ _02613_ _03940_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__and3_1
X_17611_ clknet_leaf_127_clk _00780_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_14823_ _01768_ _01769_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__nor2_1
X_18591_ clknet_leaf_185_clk _01656_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output123_A net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17542_ clknet_leaf_166_clk _00711_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_14754_ count_cycle\[19\] count_cycle\[20\] count_cycle\[21\] _01715_ VGND VGND VPWR
+ VPWR _01722_ sky130_fd_sc_hd__and4_2
X_11966_ _06434_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_158_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13705_ _07513_ _07526_ _07544_ VGND VGND VPWR VPWR _07548_ sky130_fd_sc_hd__or3_1
X_10917_ _03483_ _05213_ _05334_ _05226_ _05604_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__a221o_1
X_17473_ clknet_leaf_17_clk _00642_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_14685_ _08330_ _08331_ _08097_ VGND VGND VPWR VPWR _08332_ sky130_fd_sc_hd__a21oi_1
X_11897_ _06397_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13636_ _04642_ _04945_ _07236_ VGND VGND VPWR VPWR _07484_ sky130_fd_sc_hd__mux2_1
X_16424_ _02942_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10848_ _05292_ _05539_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08924__S _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13567_ _07418_ _07419_ VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16355_ _06961_ cpuregs.regs\[16\]\[9\] _02896_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_171_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10779_ _05273_ _05276_ _05331_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14227__A _07905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08996__A1 _03756_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15306_ _01982_ _02150_ _02152_ _02018_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__o211a_1
X_12518_ _06312_ cpuregs.regs\[28\]\[27\] _06737_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__mux2_1
X_16286_ _06961_ cpuregs.regs\[15\]\[9\] _02859_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13498_ _03275_ _07354_ _07355_ VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10474__B decoded_imm\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18025_ clknet_leaf_64_clk _00032_ VGND VGND VPWR VPWR irq_pending\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15237_ _02005_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__clkbuf_8
X_12449_ cpuregs.regs\[27\]\[27\] _06590_ _06700_ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12970__A _06319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09755__S _04078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15168_ _01936_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__buf_6
XFILLER_0_50_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13277__S _07165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14119_ _07843_ _07848_ VGND VGND VPWR VPWR _07849_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11586__A reg_pc\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15058__A _03670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15099_ _05286_ _01906_ _01956_ _01957_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__o22a_1
XANTENNA__15494__A1 _01959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15494__B2 decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14897__A _03196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09660_ _03680_ _04360_ _04363_ _03225_ _04388_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_2_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08611_ _03277_ _03249_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__nand2_1
XANTENNA__15246__B2 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17809_ clknet_leaf_62_clk _00978_ VGND VGND VPWR VPWR reg_pc\[17\] sky130_fd_sc_hd__dfxtp_2
X_09591_ _04320_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15341__S1 _02086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08542_ irq_mask\[6\] irq_pending\[6\] VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__and2b_2
XANTENNA__12210__A _06247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08473_ instr_auipc instr_lui VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09633__C1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10794__A1 _05287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11991__A0 _06266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09025_ _03213_ _03206_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__or2b_1
XFILLER_0_130_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13732__A1 _04959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09936__B1 _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11743__B1 _06101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12091__S _06496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14303__C irq_pending\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15485__B2 _03692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09927_ cpuregs.regs\[24\]\[15\] cpuregs.regs\[25\]\[15\] cpuregs.regs\[26\]\[15\]
+ cpuregs.regs\[27\]\[15\] _04085_ _04087_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__mux4_1
XANTENNA__12299__A1 _06578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16498__S _02979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10849__A2 _05398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09858_ _04578_ _04580_ _04575_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__mux2_1
XANTENNA__08911__A1 _03657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08809_ net80 VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__inv_2
X_09789_ cpuregs.regs\[0\]\[11\] cpuregs.regs\[1\]\[11\] cpuregs.regs\[2\]\[11\] cpuregs.regs\[3\]\[11\]
+ _04512_ _04513_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__mux4_1
XANTENNA__15332__S1 _02075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 _04754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11820_ _06355_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_114 net196 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_125 net202 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_136 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_147 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11751_ reg_pc\[26\] _06291_ _06093_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_80_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10702_ _05401_ _05342_ _05231_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__mux2_1
XANTENNA__14748__B1 _01717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14470_ _07898_ _07934_ _08134_ VGND VGND VPWR VPWR _08135_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11682_ _03409_ _03336_ _06066_ _06237_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13421_ _07283_ VGND VGND VPWR VPWR _07284_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11026__A2 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ _05275_ _05334_ _05309_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10234__B1 _04673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08978__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16140_ net294 net256 _02786_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__mux2_1
X_13352_ _07191_ _07212_ _07214_ _07218_ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__a211o_1
X_10564_ _04848_ _04880_ _05264_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12303_ cpuregs.regs\[25\]\[23\] _06582_ _06626_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13886__A _07675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16071_ _02633_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_114_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13283_ _06970_ cpuregs.regs\[5\]\[13\] _07165_ VGND VGND VPWR VPWR _07169_ sky130_fd_sc_hd__mux2_1
X_10495_ _05187_ _05191_ _04100_ _05199_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__a211o_4
XFILLER_0_133_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15022_ _03303_ _04022_ _04842_ _01893_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12234_ _06589_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10537__A1 _04262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11734__B1 reg_pc\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08699__B net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12165_ cpuregs.regs\[24\]\[4\] _06542_ _06534_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15476__A1 decoded_imm\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14279__A2 _07906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11116_ _05174_ _05143_ _05324_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__mux2_1
XANTENNA_output240_A net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12096_ _06503_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__clkbuf_1
X_16973_ clknet_leaf_101_clk _00147_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15571__S1 _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11047_ _05716_ _05719_ _05725_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__or3_1
X_15924_ instr_sltu _02617_ _02644_ _02653_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__a22o_1
XANTENNA__15228__A1 decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 irq[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18643_ clknet_leaf_163_clk _01703_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_15855_ _03305_ _02614_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__and2_1
XANTENNA__15779__A2 _07899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15323__S1 _01974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14806_ count_cycle\[37\] _01756_ _01717_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13334__S0 _04758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18574_ clknet_leaf_107_clk _01639_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_15786_ _03410_ _02575_ _02573_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__or3b_1
XANTENNA__10148__S0 _04758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12998_ cpuregs.regs\[3\]\[7\] _06548_ _07010_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17525_ clknet_leaf_105_clk _00694_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14737_ count_cycle\[16\] _08365_ _07826_ VGND VGND VPWR VPWR _08367_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_28_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11949_ _06096_ cpuregs.regs\[21\]\[1\] _06424_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_71_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_129_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15087__S0 _01936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17456_ clknet_leaf_133_clk _00625_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14668_ _08232_ _07969_ VGND VGND VPWR VPWR _08316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14203__A2 _07906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16407_ _06945_ cpuregs.regs\[29\]\[1\] _02932_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__mux2_1
X_13619_ _07191_ _07464_ _07466_ _07467_ _07468_ VGND VGND VPWR VPWR _07469_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_41_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17387_ clknet_leaf_130_clk _00556_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16871__S _03174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15951__A2 _02617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14599_ _08253_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10225__B1 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16338_ _02897_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10320__S0 _04123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13796__A _05174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16269_ _02860_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18008_ clknet_leaf_78_clk _01145_ VGND VGND VPWR VPWR irq_mask\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__14911__A0 net221 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11725__B1 _06093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08402__B latched_store VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08827__A_N net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13478__A0 _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13735__S _07224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09712_ cpuregs.regs\[28\]\[9\] cpuregs.regs\[29\]\[9\] cpuregs.regs\[30\]\[9\] cpuregs.regs\[31\]\[9\]
+ _04217_ _04219_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__mux4_1
XANTENNA__10387__S0 _04273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09514__A reg_pc\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09643_ _04289_ _04366_ _04371_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_171_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13325__S0 _04282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09574_ _04289_ _04304_ _04225_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_180_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08525_ _03304_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_62_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08456_ _03239_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16195__A2 net260 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11008__A2 _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12205__A1 _06569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10311__S0 _04084_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11003__B _05398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15155__B1 _01963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15250__S0 _01970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09008_ _03769_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_76_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10280_ count_instr\[57\] _04016_ _04105_ count_cycle\[57\] VGND VGND VPWR VPWR _04991_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09385__A1 _03226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15458__B2 _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_133_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15553__S1 _01974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13970_ _03354_ _07727_ _07728_ net151 VGND VGND VPWR VPWR _07746_ sky130_fd_sc_hd__a22o_1
XANTENNA__12141__A0 _06320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09688__A2 _04308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12921_ _06192_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__buf_2
X_15640_ _03379_ _07994_ _03364_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_148_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12852_ _06925_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15630__A1 _02458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14433__A2 _07947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11803_ cpuregs.waddr\[1\] cpuregs.waddr\[0\] VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__and2_1
X_12783_ _06888_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__clkbuf_1
X_15571_ _02399_ _02400_ _02401_ _02402_ _02111_ _02005_ VGND VGND VPWR VPWR _02403_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_53_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_2
X_17310_ clknet_leaf_166_clk _00484_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11734_ reg_pc\[23\] reg_pc\[22\] _06260_ reg_pc\[24\] VGND VGND VPWR VPWR _06284_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14522_ _07998_ _08162_ VGND VGND VPWR VPWR _08183_ sky130_fd_sc_hd__or2_1
X_18290_ clknet_leaf_5_clk _01358_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17241_ clknet_leaf_15_clk _00415_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11665_ _06186_ reg_next_pc\[16\] _06220_ _06222_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__a211o_4
XANTENNA__16691__S _03076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14453_ _07930_ _07932_ _08092_ VGND VGND VPWR VPWR _08119_ sky130_fd_sc_hd__and3_2
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10616_ _05315_ _05318_ _05309_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__mux2_1
X_13404_ _07232_ _07264_ _07266_ _07267_ VGND VGND VPWR VPWR _07268_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17172_ clknet_leaf_120_clk _00346_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_14384_ _08038_ _08041_ _08054_ _08055_ VGND VGND VPWR VPWR _08056_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11596_ _06116_ reg_next_pc\[9\] _06160_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output288_A net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16123_ net274 _05286_ _02771_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__mux2_1
X_13335_ _07200_ _07201_ _04211_ VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10547_ _03530_ _05250_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_12_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12724__S _06847_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15241__S0 _02069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_94_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13266_ _06953_ cpuregs.regs\[5\]\[5\] _07154_ VGND VGND VPWR VPWR _07160_ sky130_fd_sc_hd__mux2_1
X_16054_ _03402_ decoded_imm_j\[15\] _03403_ mem_rdata_q\[15\] VGND VGND VPWR VPWR
+ _02740_ sky130_fd_sc_hd__a22o_1
X_10478_ count_instr\[31\] _04012_ count_cycle\[31\] _04165_ _05182_ VGND VGND VPWR
+ VPWR _05183_ sky130_fd_sc_hd__a221o_1
XANTENNA__08503__A mem_do_wdata VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15005_ _04592_ _01869_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12217_ _06265_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__buf_2
XFILLER_0_121_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13197_ _07123_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08584__C1 decoder_trigger VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12148_ _06530_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10930__A1 _04708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15544__S1 _03642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12079_ _06343_ cpuregs.regs\[22\]\[31\] _06459_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__mux2_1
X_16956_ clknet_leaf_10_clk _00130_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09334__A _04068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15907_ mem_rdata_q\[28\] mem_rdata_q\[25\] mem_rdata_q\[26\] mem_rdata_q\[27\] VGND
+ VGND VPWR VPWR _02646_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16887_ clknet_leaf_43_clk _00083_ VGND VGND VPWR VPWR mem_wordsize\[2\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_144_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18626_ clknet_leaf_179_clk _01686_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_15838_ _03739_ _03869_ _02600_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__and3_1
XANTENNA__15082__C1 _00067_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11238__A2 _05864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18557_ clknet_leaf_184_clk _01622_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12435__A1 _06575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15769_ timer\[29\] _02561_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_44_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_170_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17508_ clknet_leaf_7_clk _00677_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_09290_ _04026_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18488_ clknet_leaf_3_clk _01553_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_14 _02412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17439_ clknet_leaf_169_clk _00608_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_25 _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15924__A2 _02617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 _05342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_47 _07154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15480__S0 _01995_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_69 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12634__S _06799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15232__S0 _01973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_963 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09509__A _04240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput110 net110 VGND VGND VPWR VPWR cpi_rs2[1] sky130_fd_sc_hd__buf_1
Xoutput121 net121 VGND VGND VPWR VPWR cpi_rs2[2] sky130_fd_sc_hd__buf_1
Xoutput132 net132 VGND VGND VPWR VPWR eoi[10] sky130_fd_sc_hd__buf_1
XFILLER_0_113_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput143 net143 VGND VGND VPWR VPWR eoi[20] sky130_fd_sc_hd__clkbuf_1
Xoutput154 net154 VGND VGND VPWR VPWR eoi[30] sky130_fd_sc_hd__buf_1
XFILLER_0_100_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14360__B2 _08033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11174__A1 _04038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput165 net165 VGND VGND VPWR VPWR mem_addr[12] sky130_fd_sc_hd__buf_1
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11174__B2 _03297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput176 net176 VGND VGND VPWR VPWR mem_addr[23] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput187 net187 VGND VGND VPWR VPWR mem_addr[4] sky130_fd_sc_hd__buf_1
Xoutput198 net198 VGND VGND VPWR VPWR mem_la_addr[14] sky130_fd_sc_hd__buf_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11774__A _06319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16776__S _03127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09626_ _04355_ VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15612__A1 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09557_ _04279_ _04286_ _04287_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_2
X_08508_ _03239_ _03282_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__nor2_2
XFILLER_0_65_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09488_ cpuregs.regs\[20\]\[4\] cpuregs.regs\[21\]\[4\] cpuregs.regs\[22\]\[4\] cpuregs.regs\[23\]\[4\]
+ _04217_ _04219_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08439_ _03224_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_136_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15471__S0 _01999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11450_ _06041_ irq_pending\[13\] _06043_ net5 VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10401_ instr_retirq _05107_ _05108_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11381_ _05990_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__inv_2
XANTENNA__10853__A _05292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13120_ _06941_ cpuregs.regs\[4\]\[0\] _07082_ VGND VGND VPWR VPWR _07083_ sky130_fd_sc_hd__mux2_1
X_10332_ count_cycle\[26\] _04165_ _05041_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14044__B _07778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13051_ _07045_ VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__buf_6
X_10263_ cpuregs.regs\[16\]\[24\] cpuregs.regs\[17\]\[24\] cpuregs.regs\[18\]\[24\]
+ cpuregs.regs\[19\]\[24\] _04071_ _04073_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11165__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16540__A _03003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12002_ _06453_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09853__S _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10194_ _04296_ _04894_ _04898_ _04907_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__a31o_2
XANTENNA__15526__S1 _02075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11684__A _06239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16810_ _03147_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__clkbuf_1
X_17790_ clknet_leaf_84_clk _00959_ VGND VGND VPWR VPWR count_instr\[61\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12114__A0 _06216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16741_ _07007_ cpuregs.regs\[19\]\[31\] _03075_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__mux2_1
X_13953_ _07734_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_161_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12904_ _06956_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__clkbuf_1
X_16672_ _03073_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__clkbuf_1
X_13884_ _07686_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__clkbuf_1
X_18411_ clknet_leaf_124_clk _01476_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_15623_ _02450_ _02451_ _03709_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12835_ _06916_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output203_A net203 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_26_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18342_ clknet_leaf_37_clk _01410_ VGND VGND VPWR VPWR mem_16bit_buffer\[13\] sky130_fd_sc_hd__dfxtp_1
X_15554_ cpuregs.regs\[0\]\[27\] cpuregs.regs\[1\]\[27\] cpuregs.regs\[2\]\[27\] cpuregs.regs\[3\]\[27\]
+ _02085_ _02086_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__mux4_1
X_12766_ _06879_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14505_ _08148_ _08153_ VGND VGND VPWR VPWR _08167_ sky130_fd_sc_hd__and2_1
X_11717_ reg_pc\[22\] _06260_ _06101_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18273_ clknet_leaf_25_clk _01344_ VGND VGND VPWR VPWR decoded_imm\[31\] sky130_fd_sc_hd__dfxtp_2
X_12697_ _06208_ cpuregs.regs\[12\]\[14\] _06836_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15485_ _02316_ _02318_ _02321_ _03692_ _01968_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15462__S0 _01979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17224_ clknet_leaf_133_clk _00398_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11648_ _06207_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__buf_2
X_14436_ _07930_ _08092_ _07986_ VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput12 irq[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput23 irq[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
Xinput34 mem_rdata[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_108_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput45 mem_rdata[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17155_ clknet_leaf_134_clk _00329_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14367_ _08038_ _08039_ VGND VGND VPWR VPWR _08040_ sky130_fd_sc_hd__nand2_1
X_11579_ reg_pc\[7\] _06137_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__and2_1
Xinput56 mem_rdata[30] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
XFILLER_0_13_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16867__A0 _06582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16106_ _02767_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__clkbuf_1
X_13318_ _07005_ cpuregs.regs\[5\]\[30\] _07153_ VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__mux2_1
XANTENNA__09329__A _04063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14298_ irq_pending\[28\] irq_pending\[29\] irq_pending\[30\] irq_pending\[31\] VGND
+ VGND VPWR VPWR _07975_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17086_ clknet_leaf_172_clk _00260_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16037_ decoded_imm\[7\] _02711_ _02730_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13249_ _07150_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11156__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09444__S1 _04086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15517__S1 _02031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16095__A1 _03309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13285__S _07165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08790_ _03500_ net69 _03516_ _03549_ _03555_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__a221o_1
X_17988_ clknet_leaf_105_clk _01125_ VGND VGND VPWR VPWR irq_mask\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15842__A1 instr_lui VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16939_ clknet_leaf_110_clk _00120_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08955__S0 _03649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10131__A2 _04014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09411_ _04011_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__clkbuf_4
X_18609_ clknet_leaf_165_clk _01674_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_17_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09342_ _04063_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09273_ _04009_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15453__S0 _02069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14030__B1 _07759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14581__A1 _07952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10198__A2 _04890_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11395__A1 _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_950 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15530__B1 _02197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11147__A1 _03407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11147__B2 _04422_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08797__B net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08988_ _03739_ _03749_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__nand2_1
XANTENNA__15833__A1 decoded_imm_j\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09512__A1 _04010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10950_ _03481_ _05397_ _05213_ _03480_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_168_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09609_ _04105_ count_cycle\[38\] _04009_ _04338_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_104_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15597__B1 _02427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10881_ net72 _04602_ _05264_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10848__A _05292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10673__A3 _04466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12539__S _06752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12620_ _06175_ cpuregs.regs\[30\]\[10\] _06799_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Left_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12551_ _06751_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11502_ _06071_ _06075_ reg_next_pc\[0\] VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__o21a_1
X_15270_ net100 _02081_ _02118_ _02119_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__o22a_1
X_12482_ _06714_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__buf_6
XANTENNA__14021__B1 _07759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09579__A1 _04271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14221_ _07901_ VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__clkbuf_4
X_11433_ irq_mask\[6\] _06030_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09674__S1 _04091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14152_ count_instr\[51\] _07869_ _07834_ VGND VGND VPWR VPWR _07873_ sky130_fd_sc_hd__o21ai_1
X_11364_ _05969_ _03634_ _03874_ _05977_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15585__S _01907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13103_ _07073_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__clkbuf_1
X_10315_ cpuregs.regs\[20\]\[26\] cpuregs.regs\[21\]\[26\] cpuregs.regs\[22\]\[26\]
+ cpuregs.regs\[23\]\[26\] _04123_ _04124_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__mux4_1
X_14083_ count_instr\[31\] count_instr\[30\] count_instr\[29\] _07818_ VGND VGND VPWR
+ VPWR _07824_ sky130_fd_sc_hd__and4_2
X_11295_ _05913_ _05915_ _05918_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11138__A1 _04040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_168_Left_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17911_ clknet_leaf_85_clk _01080_ VGND VGND VPWR VPWR count_cycle\[56\] sky130_fd_sc_hd__dfxtp_1
X_13034_ cpuregs.regs\[3\]\[24\] _06584_ _07032_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__mux2_1
X_10246_ _04954_ _04957_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__xor2_1
XANTENNA__09200__A0 mem_rdata_q\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16077__A1 decoded_imm\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16077__B2 mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17842_ clknet_leaf_60_clk _01011_ VGND VGND VPWR VPWR reg_next_pc\[19\] sky130_fd_sc_hd__dfxtp_1
X_10177_ cpuregs.regs\[20\]\[22\] cpuregs.regs\[21\]\[22\] cpuregs.regs\[22\]\[22\]
+ cpuregs.regs\[23\]\[22\] _04281_ _04470_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17773_ clknet_leaf_95_clk _00942_ VGND VGND VPWR VPWR count_instr\[44\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_124_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14985_ _04227_ _04298_ _04306_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__or3_4
XANTENNA__10649__A0 _04342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15614__A _03709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16724_ _03101_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13936_ _07722_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08927__S _03664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_1019 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_46 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09612__A net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16655_ cpuregs.regs\[1\]\[22\] _06273_ _03062_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__mux2_1
X_13867_ cpuregs.regs\[0\]\[30\] VGND VGND VPWR VPWR _07673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12449__S _06700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15606_ _02434_ _02435_ _02110_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__mux2_1
X_12818_ _06096_ cpuregs.regs\[6\]\[1\] _06906_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16586_ _03028_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13798_ _07633_ _07634_ _07620_ _07625_ VGND VGND VPWR VPWR _07635_ sky130_fd_sc_hd__o211a_1
XANTENNA__09806__A2 _04165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18325_ clknet_leaf_39_clk _01393_ VGND VGND VPWR VPWR mem_la_secondword sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15537_ cpuregs.regs\[0\]\[26\] cpuregs.regs\[1\]\[26\] cpuregs.regs\[2\]\[26\] cpuregs.regs\[3\]\[26\]
+ _02046_ _02047_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12749_ cpuregs.regs\[9\]\[1\] _06536_ _06869_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12973__A _06327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15435__S0 _01918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18256_ clknet_leaf_25_clk _01327_ VGND VGND VPWR VPWR decoded_imm\[14\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08490__A1 _03226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15468_ _01984_ _02305_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17207_ clknet_leaf_155_clk _00381_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_14419_ _08084_ _08086_ VGND VGND VPWR VPWR _08088_ sky130_fd_sc_hd__nand2_1
X_18187_ clknet_leaf_43_clk _01258_ VGND VGND VPWR VPWR instr_bltu sky130_fd_sc_hd__dfxtp_1
XANTENNA__12184__S _06555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15399_ _02235_ _02237_ _02240_ _02017_ _01968_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__a221o_2
Xmax_cap301 _04099_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__buf_4
XFILLER_0_25_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17138_ clknet_leaf_113_clk _00312_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15495__S _03272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14315__A1 decoder_trigger VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09960_ reg_pc\[15\] decoded_imm\[15\] _04679_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12912__S _06943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17069_ clknet_leaf_120_clk _00243_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_6_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_2
X_08911_ _03657_ _03665_ _03668_ _03673_ _03675_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__a221o_1
X_09891_ _04420_ _04612_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__or2_2
XFILLER_0_97_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08842_ _03606_ _03607_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__nor2_1
XANTENNA__12213__A _06256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08773_ net121 net89 VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__and2b_1
XFILLER_0_68_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12359__S _06652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09258__B1 _03763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14251__B1 _07942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09325_ _04059_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09353__S0 _04085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12801__A1 _06588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15897__C _02610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09256_ mem_rdata_q\[29\] _03994_ _03757_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__mux2_1
XANTENNA__13698__B decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09187_ _03775_ _03916_ _03934_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__or3_1
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09430__B1 _04163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09981__A1 _04231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12822__S _06906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16090__A _03228_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10591__A2 _03518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10100_ reg_pc\[17\] decoded_imm\[17\] VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11080_ _05218_ _05756_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08601__A instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16059__A1 decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10031_ reg_pc\[18\] decoded_imm\[18\] VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09733__A1 _03385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15267__C1 _01969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ count_cycle\[25\] _01729_ count_cycle\[26\] VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_86_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11982_ _06232_ cpuregs.regs\[21\]\[17\] _06435_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11039__A2_N _05367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13721_ _07232_ _07562_ _07563_ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__o21a_1
XANTENNA__09432__A _03253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10933_ net107 net75 VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10578__A _05251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12269__S _06604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15034__A2 _01865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16440_ _06978_ cpuregs.regs\[29\]\[17\] _02943_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__mux2_1
X_10864_ _03494_ _05367_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__or2_1
X_13652_ net79 decoded_imm\[20\] VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13889__A _07675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12603_ _06105_ cpuregs.regs\[30\]\[2\] _06788_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16371_ _02914_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__clkbuf_1
X_10795_ _03513_ _05367_ _05357_ _03515_ _05489_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__o221a_1
X_13583_ _07432_ _07433_ _07434_ VGND VGND VPWR VPWR _07435_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18110_ clknet_leaf_81_clk _01214_ VGND VGND VPWR VPWR timer\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11901__S _06398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15322_ cpuregs.regs\[4\]\[14\] cpuregs.regs\[5\]\[14\] cpuregs.regs\[6\]\[14\] cpuregs.regs\[7\]\[14\]
+ _01979_ _01980_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12534_ _06754_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18041_ clknet_leaf_78_clk _00018_ VGND VGND VPWR VPWR irq_pending\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__14545__A1 _07943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15253_ _01982_ _02100_ _02102_ _02018_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12465_ _06717_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14204_ _03188_ _06107_ VGND VGND VPWR VPWR _07910_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_117_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11416_ cpuregs.raddr1\[3\] _06006_ _06020_ _06022_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__o22a_1
X_12396_ _06680_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__clkbuf_1
X_15184_ _02029_ _02033_ _02036_ _02037_ _01969_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08775__A2 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14135_ count_instr\[46\] _07859_ _07834_ VGND VGND VPWR VPWR _07861_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11347_ _03748_ _03879_ _03844_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output78_A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14066_ _07811_ _07812_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__nor2_1
X_11278_ _03475_ _05829_ _05905_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__o21ai_4
XANTENNA__08511__A _03293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09724__A1 _04010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10229_ irq_mask\[23\] _04308_ timer\[23\] instr_timer _04026_ VGND VGND VPWR VPWR
+ _04942_ sky130_fd_sc_hd__a221o_1
X_13017_ cpuregs.regs\[3\]\[16\] _06567_ _07021_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__mux2_1
X_17825_ clknet_leaf_22_clk _00994_ VGND VGND VPWR VPWR reg_next_pc\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13563__S _07374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15344__A _02066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17756_ clknet_leaf_82_clk _00925_ VGND VGND VPWR VPWR count_instr\[27\] sky130_fd_sc_hd__dfxtp_1
X_14968_ irq_active _01860_ _01859_ _04150_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10098__A1 _04391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16707_ _03092_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09342__A _04063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13919_ _07691_ _07710_ VGND VGND VPWR VPWR _07711_ sky130_fd_sc_hd__and2_1
XANTENNA__11295__B1 _05918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09583__S0 _04217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17687_ clknet_leaf_164_clk _00856_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14899_ _01821_ _01822_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__nand2_2
XFILLER_0_159_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16638_ cpuregs.regs\[1\]\[14\] _06207_ _03051_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13036__A1 _06586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13587__A2 _05259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09996__B decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16569_ _03019_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11598__A1 reg_pc\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11811__S _06348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09110_ _03736_ _03869_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_44_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18308_ clknet_leaf_35_clk _01376_ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09660__B1 _04363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10270__A1 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09041_ _03801_ _03802_ _03203_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18239_ clknet_leaf_23_clk _01310_ VGND VGND VPWR VPWR cpuregs.raddr2\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__14536__A1 _08071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09638__S1 _04276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09412__B1 _04017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09943_ _04660_ _04661_ _04663_ _04268_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08518__A2 _03276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09874_ reg_pc\[13\] decoded_imm\[13\] VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__nand2_1
XANTENNA__11522__A1 _06066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _03453_ _03456_ _03582_ _03590_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__o31a_1
X_08756_ _03521_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11286__B1 _05911_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12089__S _06496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08687_ _03449_ _03452_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__nand2_1
XANTENNA__16784__S _03127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16213__A1 _03218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_975 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09326__S0 _04057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09308_ reg_next_pc\[0\] decoded_imm\[0\] VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10580_ _05231_ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__or2b_1
XFILLER_0_134_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09651__B1 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14527__A1 _07942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09239_ _03959_ _03978_ _03960_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12250_ _06083_ _06422_ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09403__B1 _04068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11210__A0 _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11201_ _05842_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__buf_4
XANTENNA__09954__A1 _03638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09954__B2 _03302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12181_ _06553_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12552__S _06763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11132_ _05413_ _05803_ _05804_ _05251_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_112_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ _03452_ _05739_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__or2_1
XANTENNA__13502__A2 _04447_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15940_ instr_rdcycle _02650_ _02659_ _02665_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__a22o_1
XANTENNA__12710__A0 _06257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10014_ cpuregs.regs\[8\]\[17\] cpuregs.regs\[9\]\[17\] cpuregs.regs\[10\]\[17\]
+ cpuregs.regs\[11\]\[17\] _04280_ _04059_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__mux4_1
X_15871_ instr_bltu _02618_ _02622_ _02626_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__a22o_1
X_17610_ clknet_leaf_175_clk _00779_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_14822_ count_cycle\[42\] _01765_ _01723_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15164__A _02017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18590_ clknet_leaf_173_clk _01655_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17541_ clknet_leaf_1_clk _00710_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_14753_ _01721_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11965_ _06166_ cpuregs.regs\[21\]\[9\] _06424_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output116_A net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _04945_ _07271_ _07541_ _07547_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__o22a_1
XFILLER_0_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10916_ _03484_ _05398_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__nor2_1
X_17472_ clknet_leaf_176_clk _00641_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14684_ _08232_ _07971_ VGND VGND VPWR VPWR _08331_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11896_ _06166_ cpuregs.regs\[20\]\[9\] _06387_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16423_ _06961_ cpuregs.regs\[29\]\[9\] _02932_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__mux2_1
X_13635_ _04754_ _05261_ _07451_ _07279_ VGND VGND VPWR VPWR _07483_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10847_ _05331_ _05276_ _05423_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16354_ _02905_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__clkbuf_1
X_13566_ net72 decoded_imm\[14\] VGND VGND VPWR VPWR _07419_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10778_ _05298_ _05471_ _05473_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_136_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09642__B1 _04237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15305_ _01989_ _02151_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__or2_1
X_12517_ _06744_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16285_ _02868_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__clkbuf_1
X_13497_ _07352_ _07353_ VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18024_ clknet_leaf_104_clk _00031_ VGND VGND VPWR VPWR irq_pending\[8\] sky130_fd_sc_hd__dfxtp_1
X_15236_ cpuregs.regs\[0\]\[9\] cpuregs.regs\[1\]\[9\] cpuregs.regs\[2\]\[9\] cpuregs.regs\[3\]\[9\]
+ _02085_ _02086_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12448_ _06707_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15167_ cpuregs.regs\[28\]\[6\] cpuregs.regs\[29\]\[6\] cpuregs.regs\[30\]\[6\] cpuregs.regs\[31\]\[6\]
+ _01990_ _01992_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__mux4_1
XANTENNA__12462__S _06715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12379_ _06670_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11752__A1 reg_pc\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14118_ count_instr\[42\] count_instr\[41\] count_instr\[40\] VGND VGND VPWR VPWR
+ _07848_ sky130_fd_sc_hd__and3_1
XANTENNA__09337__A _04071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15098_ is_slli_srli_srai cpuregs.raddr2\[1\] decoded_imm\[1\] _01933_ _01934_ VGND
+ VGND VPWR VPWR _01957_ sky130_fd_sc_hd__a221o_1
XANTENNA__16869__S _03174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14049_ count_instr\[20\] _07799_ VGND VGND VPWR VPWR _07801_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14897__B net299 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_105_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13293__S _07165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08610_ _03384_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__buf_4
XANTENNA__15074__A _03277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17808_ clknet_leaf_62_clk _00977_ VGND VGND VPWR VPWR reg_pc\[16\] sky130_fd_sc_hd__dfxtp_2
X_09590_ _04063_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08541_ irq_mask\[22\] irq_pending\[22\] VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__and2b_2
X_17739_ clknet_leaf_96_clk _00908_ VGND VGND VPWR VPWR count_instr\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08472_ instr_lh instr_jalr instr_jal _03255_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__or4_1
XFILLER_0_147_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11440__B1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09024_ _03779_ _03785_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11777__A reg_pc\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09936__A1 _04053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12372__S _06663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11743__A1 reg_pc\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12940__A0 _06980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09926_ cpuregs.regs\[28\]\[15\] cpuregs.regs\[29\]\[15\] cpuregs.regs\[30\]\[15\]
+ cpuregs.regs\[31\]\[15\] _04477_ _04478_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_123_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09857_ cpuregs.regs\[24\]\[13\] cpuregs.regs\[25\]\[13\] cpuregs.regs\[26\]\[13\]
+ cpuregs.regs\[27\]\[13\] _04579_ _04284_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14600__B _07959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08808_ _03461_ _03462_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__nand2_1
X_09788_ _04283_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__clkbuf_8
X_08739_ net100 net68 VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__nor2_1
XANTENNA__14996__A1 _03303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_104 _04758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 net196 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_137 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15712__A _02484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_148 net203 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11750_ _06298_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10701_ net93 net92 _03609_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11681_ reg_out\[18\] alu_out_q\[18\] _06068_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__mux2_1
XANTENNA__12547__S _06752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13420_ _07221_ VGND VGND VPWR VPWR _07283_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_153_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ instr_sra instr_srai _05205_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__o21a_4
XFILLER_0_165_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09624__B1 irq_pending\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10234__B2 _04946_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10563_ _05262_ _05265_ _05266_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__mux2_1
X_13351_ _04251_ _03313_ _07217_ _04118_ _05260_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12302_ _06629_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16070_ decoded_imm\[21\] _02650_ _02746_ mem_rdata_q\[21\] _02749_ VGND VGND VPWR
+ VPWR _01334_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_114_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13282_ _07168_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__clkbuf_1
X_10494_ _04289_ _05194_ _05198_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13184__A0 _07007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15021_ irq_mask\[20\] _01863_ _01714_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15159__A _01936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12282__S _06615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12233_ cpuregs.regs\[24\]\[26\] _06588_ _06576_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10537__A2 _04342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12931__A0 _06974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12164_ _06124_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__buf_2
XFILLER_0_102_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16689__S _03076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15476__A2 _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11115_ _05575_ _05700_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__nor2_1
XANTENNA__16673__A1 _06342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14133__C1 _07775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16972_ clknet_leaf_179_clk _00146_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_12095_ _06141_ cpuregs.regs\[23\]\[6\] _06496_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__mux2_1
X_11046_ _05723_ _05724_ _05218_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__a21oi_1
X_15923_ instr_slt _02617_ _02641_ _02653_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__a22o_1
XANTENNA__09786__S0 _04274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output233_A net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15228__A2 _02009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18642_ clknet_leaf_119_clk _01702_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_129_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _02612_ _02613_ _03940_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__nor3_1
XFILLER_0_36_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14436__B1 _07986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14805_ _01756_ _01757_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18573_ clknet_leaf_161_clk _01638_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13334__S1 _04759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15785_ _03317_ _03364_ _07984_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12997_ _07017_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16718__A _03075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10148__S1 _04759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17524_ clknet_leaf_152_clk _00693_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_14736_ _08365_ _08366_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11948_ _06425_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09863__B1 _04068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15087__S1 _03647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11670__B1 _06093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17455_ clknet_leaf_144_clk _00624_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12457__S _06677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14667_ _08288_ _08306_ _08307_ _08311_ VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__a31o_1
X_11879_ _06388_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16406_ _02933_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13618_ _07304_ _04738_ _07305_ reg_pc\[17\] _07283_ VGND VGND VPWR VPWR _07468_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17386_ clknet_leaf_182_clk _00555_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14598_ _08245_ _08252_ VGND VGND VPWR VPWR _08253_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10225__A1 _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16337_ _06941_ cpuregs.regs\[16\]\[0\] _02896_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13549_ _04566_ _07403_ _07374_ VGND VGND VPWR VPWR _07404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10320__S1 _04124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13796__B decoded_imm\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16268_ _06941_ cpuregs.regs\[15\]\[0\] _02859_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18007_ clknet_leaf_78_clk _01144_ VGND VGND VPWR VPWR irq_mask\[23\] sky130_fd_sc_hd__dfxtp_1
X_15219_ cpuregs.regs\[12\]\[8\] cpuregs.regs\[13\]\[8\] cpuregs.regs\[14\]\[8\] cpuregs.regs\[15\]\[8\]
+ _02069_ _02070_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__mux4_1
XANTENNA__15069__A _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16199_ _02814_ _02819_ _02820_ _02676_ net298 VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__a32o_1
XFILLER_0_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12922__A0 _06968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10084__S0 _04273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16599__S _03026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09711_ _04432_ _04434_ _04437_ _04206_ _04296_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__a221o_1
XANTENNA__10387__S1 _04283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09642_ _04328_ _04370_ _04237_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__a21o_1
XANTENNA__09514__B decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09573_ _04302_ _04303_ _04223_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__mux2_1
XANTENNA__13325__S1 _04285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08524_ _03277_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__buf_4
XFILLER_0_148_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08455_ _03196_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11661__B1 _06101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11008__A3 _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10311__S1 _04086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15155__A1 decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_836 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13198__S _07118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15250__S1 _01971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09007_ _03767_ _03768_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09385__A2 _04112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16655__A1 _06273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12830__S _06906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14611__A _07988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09705__A _04430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09909_ _04227_ _04630_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__or2_4
X_12920_ _06967_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10350__S _04211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12851_ _06232_ cpuregs.regs\[6\]\[17\] _06917_ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__mux2_1
X_11802_ _06344_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ cpuregs.regs\[0\]\[28\] cpuregs.regs\[1\]\[28\] cpuregs.regs\[2\]\[28\] cpuregs.regs\[3\]\[28\]
+ _01976_ _01977_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__mux4_1
XANTENNA__09845__B1 _04568_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12782_ cpuregs.regs\[9\]\[17\] _06569_ _06880_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_140_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_675 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14521_ _08180_ _08181_ _08012_ VGND VGND VPWR VPWR _08182_ sky130_fd_sc_hd__a21bo_1
X_11733_ reg_pc\[24\] reg_pc\[23\] _06268_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16040__C1 _02634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17240_ clknet_leaf_176_clk _00414_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14452_ _07898_ _07932_ _08050_ _07947_ reg_next_pc\[12\] VGND VGND VPWR VPWR _08118_
+ sky130_fd_sc_hd__a32o_1
X_11664_ _03409_ _03330_ _06066_ _06221_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__a22o_1
X_13403_ _03312_ _04360_ _05259_ _07254_ VGND VGND VPWR VPWR _07267_ sky130_fd_sc_hd__a31o_1
XFILLER_0_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15588__S _02110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10615_ _05316_ _05317_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17171_ clknet_leaf_109_clk _00345_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_14383_ _03368_ _03378_ VGND VGND VPWR VPWR _08055_ sky130_fd_sc_hd__nand2_2
X_11595_ irq_state\[1\] _03323_ _06098_ _06159_ _06118_ VGND VGND VPWR VPWR _06160_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16122_ _02778_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16343__A0 _06949_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13334_ cpuregs.regs\[0\]\[0\] cpuregs.regs\[1\]\[0\] cpuregs.regs\[2\]\[0\] cpuregs.regs\[3\]\[0\]
+ _04758_ _04759_ VGND VGND VPWR VPWR _07201_ sky130_fd_sc_hd__mux4_1
X_10546_ _05226_ _05210_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__or2_2
XFILLER_0_135_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13157__A0 _06980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15241__S1 _02070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16053_ decoded_imm\[14\] _02720_ _02736_ _02739_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13265_ _07159_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__clkbuf_1
X_10477_ count_instr\[63\] _04104_ _04105_ count_cycle\[63\] VGND VGND VPWR VPWR _05182_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15004_ irq_mask\[12\] _01880_ _01883_ _01876_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__a211o_1
X_12216_ _06577_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__clkbuf_1
X_13196_ _06951_ cpuregs.regs\[8\]\[4\] _07118_ VGND VGND VPWR VPWR _07123_ sky130_fd_sc_hd__mux2_1
XANTENNA__16646__A1 _06239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12380__A1 _06590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12147_ _06343_ cpuregs.regs\[23\]\[31\] _06495_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__mux2_1
XANTENNA__10930__A2 _04642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09759__S0 _04232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12078_ _06493_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__clkbuf_1
X_16955_ clknet_leaf_10_clk _00129_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11029_ _03469_ _03473_ _05677_ _05708_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__a31o_1
X_15906_ mem_rdata_q\[29\] mem_rdata_q\[30\] mem_rdata_q\[31\] VGND VGND VPWR VPWR
+ _02645_ sky130_fd_sc_hd__or3_1
X_16886_ clknet_leaf_39_clk _00082_ VGND VGND VPWR VPWR mem_wordsize\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18625_ clknet_leaf_18_clk _01685_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15837_ _03816_ _03916_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12976__A _06335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15352__A _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15768_ _05107_ _02486_ _02563_ _02545_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__o211a_1
X_18556_ clknet_leaf_187_clk _01621_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11238__A3 _05868_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09350__A _04084_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10446__B2 _04013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14719_ count_cycle\[10\] _08353_ _07826_ VGND VGND VPWR VPWR _08355_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11643__B1 _06093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17507_ clknet_leaf_11_clk _00676_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12187__S _06555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09931__S0 _04232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18487_ clknet_leaf_11_clk _01552_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10496__A _05200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15699_ timer\[11\] _02511_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__xor2_1
XANTENNA__10541__S1 _05244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17438_ clknet_leaf_125_clk _00607_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_15 _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_26 _04397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12199__A1 _06565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 _05864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15480__S1 _01937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _07944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17369_ clknet_leaf_100_clk _00538_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_59 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13600__A _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15232__S1 _01974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput100 net100 VGND VGND VPWR VPWR cpi_rs2[10] sky130_fd_sc_hd__buf_1
XFILLER_0_141_975 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput111 net111 VGND VGND VPWR VPWR cpi_rs2[20] sky130_fd_sc_hd__buf_1
XFILLER_0_11_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput122 net122 VGND VGND VPWR VPWR cpi_rs2[30] sky130_fd_sc_hd__clkbuf_1
Xoutput133 net133 VGND VGND VPWR VPWR eoi[11] sky130_fd_sc_hd__buf_1
XFILLER_0_3_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14360__A2 _07947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput144 net144 VGND VGND VPWR VPWR eoi[21] sky130_fd_sc_hd__buf_1
Xoutput155 net155 VGND VGND VPWR VPWR eoi[31] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11174__A2 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput166 net166 VGND VGND VPWR VPWR mem_addr[13] sky130_fd_sc_hd__clkbuf_1
XANTENNA__16098__C1 _03891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput177 net177 VGND VGND VPWR VPWR mem_addr[24] sky130_fd_sc_hd__clkbuf_1
Xoutput188 net188 VGND VGND VPWR VPWR mem_addr[5] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput199 net199 VGND VGND VPWR VPWR mem_la_addr[15] sky130_fd_sc_hd__clkbuf_1
XANTENNA__16101__A3 _03885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13320__A0 _07007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09625_ _04341_ _04346_ _04354_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__or3_1
XANTENNA__11882__A0 _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15612__A2 _01906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09556_ _04065_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10437__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08507_ _03276_ _03289_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__nand2_1
XANTENNA__09922__S0 _04281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12097__S _06496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09487_ _04218_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08438_ net66 _03223_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13387__A0 _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15471__S1 _02000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10400_ irq_mask\[28\] instr_maskirq timer\[28\] instr_timer _04025_ VGND VGND VPWR
+ VPWR _05108_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11380_ _03787_ _03770_ _05989_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__or3_2
XFILLER_0_144_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10853__B _05544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10331_ count_instr\[26\] _04145_ _04009_ _05040_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__a211o_1
XANTENNA__09419__B decoded_imm\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14887__B1 _07224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10262_ cpuregs.regs\[20\]\[24\] cpuregs.regs\[21\]\[24\] cpuregs.regs\[22\]\[24\]
+ cpuregs.regs\[23\]\[24\] _04071_ _04073_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__mux4_1
X_13050_ _06346_ _06904_ VGND VGND VPWR VPWR _07045_ sky130_fd_sc_hd__nand2_4
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11165__A2 _04710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12001_ _06304_ cpuregs.regs\[21\]\[26\] _06446_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12560__S _06763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10193_ _04133_ _04906_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__nand2_1
XANTENNA__09435__A instr_retirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15300__A1 _02020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16740_ _03109_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__clkbuf_1
X_13952_ _07714_ _07733_ VGND VGND VPWR VPWR _07734_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_161_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12903_ _06955_ cpuregs.regs\[31\]\[6\] _06943_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__mux2_1
XANTENNA__10220__S0 _04281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16671_ cpuregs.regs\[1\]\[30\] _06335_ _03039_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13883_ _07675_ _07685_ VGND VGND VPWR VPWR _07686_ sky130_fd_sc_hd__and2_1
X_15622_ cpuregs.regs\[12\]\[31\] cpuregs.regs\[13\]\[31\] cpuregs.regs\[14\]\[31\]
+ cpuregs.regs\[15\]\[31\] _03645_ _03647_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18410_ clknet_leaf_123_clk _01475_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12834_ _06166_ cpuregs.regs\[6\]\[9\] _06906_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18341_ clknet_leaf_36_clk _01409_ VGND VGND VPWR VPWR mem_16bit_buffer\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15553_ cpuregs.regs\[4\]\[27\] cpuregs.regs\[5\]\[27\] cpuregs.regs\[6\]\[27\] cpuregs.regs\[7\]\[27\]
+ _01973_ _01974_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__mux4_1
X_12765_ cpuregs.regs\[9\]\[9\] _06552_ _06869_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14504_ _08164_ _08165_ VGND VGND VPWR VPWR _08166_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11716_ reg_pc\[22\] _06260_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18272_ clknet_leaf_25_clk _01343_ VGND VGND VPWR VPWR decoded_imm\[30\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_126_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15484_ _02319_ _02320_ _03653_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12696_ _06840_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17223_ clknet_leaf_144_clk _00397_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15462__S1 _01980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14435_ _07930_ _08092_ VGND VGND VPWR VPWR _08102_ sky130_fd_sc_hd__and2_1
X_11647_ _06186_ reg_next_pc\[14\] _06204_ _06206_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__a211o_2
XFILLER_0_65_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 irq[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14516__A decoded_imm_j\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13420__A _07221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput24 irq[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17154_ clknet_leaf_185_clk _00328_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16316__A0 _06991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10287__S0 _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput35 mem_rdata[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_80_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14366_ decoded_imm_j\[5\] _07917_ VGND VGND VPWR VPWR _08039_ sky130_fd_sc_hd__or2_1
Xinput46 mem_rdata[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
XANTENNA__08514__A mem_do_wdata VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11578_ _06116_ reg_next_pc\[7\] _06144_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput57 mem_rdata[31] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_2
XFILLER_0_123_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16105_ is_alu_reg_reg _02766_ _03635_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__mux2_1
XANTENNA__10600__A1 _04040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13317_ _07186_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_168_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10529_ _04419_ _04456_ _04466_ _04532_ _05230_ _05232_ VGND VGND VPWR VPWR _05233_
+ sky130_fd_sc_hd__mux4_1
X_17085_ clknet_leaf_1_clk _00259_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[4\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_172_Right_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14297_ irq_pending\[16\] irq_pending\[17\] irq_pending\[18\] irq_pending\[19\] VGND
+ VGND VPWR VPWR _07974_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14878__B1 _03240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16036_ _02715_ decoded_imm_j\[7\] _02726_ mem_rdata_q\[27\] _02634_ VGND VGND VPWR
+ VPWR _02730_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13248_ _07003_ cpuregs.regs\[8\]\[29\] _07140_ VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16619__A1 _06131_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12470__S _06715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10364__B1 _04009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13179_ _07113_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09345__A _00073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16877__S _03174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17987_ clknet_leaf_105_clk _01124_ VGND VGND VPWR VPWR irq_mask\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16938_ clknet_leaf_161_clk _00119_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10211__S0 _04512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08955__S1 _03643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16869_ _06584_ cpuregs.regs\[14\]\[24\] _03174_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__mux2_1
XANTENNA__10762__S1 _05287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09410_ irq_mask\[2\] _04022_ timer\[2\] _04024_ _04027_ VGND VGND VPWR VPWR _04144_
+ sky130_fd_sc_hd__a221o_1
X_18608_ clknet_leaf_111_clk _01673_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09809__B1 _04507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13605__B2 _07283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09080__A _03229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09904__S0 _04290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09341_ cpuregs.regs\[16\]\[1\] cpuregs.regs\[17\]\[1\] cpuregs.regs\[18\]\[1\] cpuregs.regs\[19\]\[1\]
+ _04072_ _04074_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__mux4_1
X_18539_ clknet_leaf_119_clk _01604_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08408__B irq_state\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15358__A1 _01982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09272_ _03252_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_16_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_132_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15453__S1 _02070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12645__S _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14581__A2 _07954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09993__C1 _04712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14869__B1 _01714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_147_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15530__A1 decoded_imm\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13984__B _07755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11147__A2 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12380__S _06663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08987_ _03743_ _03748_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__or2_2
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10658__A1 _05225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09608_ count_instr\[38\] _04015_ instr_rdinstr count_instr\[6\] VGND VGND VPWR VPWR
+ _04338_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15597__A1 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10880_ _05444_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09539_ count_instr\[37\] _04016_ count_cycle\[5\] _04013_ _04269_ VGND VGND VPWR
+ VPWR _04270_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15720__A _04702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12550_ _06762_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11501_ _06074_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_109_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12481_ _06725_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14336__A _07972_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14220_ reg_pc\[7\] _07906_ _07921_ _07912_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__a22o_1
XANTENNA__09579__A2 _04307_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11432_ _06029_ irq_pending\[5\] _06033_ net28 VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13780__A0 _05086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12583__A1 _06586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14151_ count_instr\[51\] _07865_ _07868_ VGND VGND VPWR VPWR _07872_ sky130_fd_sc_hd__and3_1
XANTENNA__09984__C1 _04027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11363_ _03979_ _05976_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13102_ _06993_ cpuregs.regs\[7\]\[24\] _07068_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10314_ _04052_ _05023_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__nand2_1
X_14082_ _07823_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__clkbuf_1
X_11294_ reg_next_pc\[23\] reg_out\[23\] _05898_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__mux2_2
XFILLER_0_120_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17910_ clknet_leaf_85_clk _01079_ VGND VGND VPWR VPWR count_cycle\[55\] sky130_fd_sc_hd__dfxtp_1
X_13033_ _07036_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__clkbuf_1
X_10245_ _04955_ _04956_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__nand2_1
XANTENNA__12290__S _06615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09200__A1 _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10176_ count_instr\[22\] _04145_ count_cycle\[22\] _04013_ _04889_ VGND VGND VPWR
+ VPWR _04890_ sky130_fd_sc_hd__a221o_1
X_17841_ clknet_leaf_60_clk _01010_ VGND VGND VPWR VPWR reg_next_pc\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_output146_A net146 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15285__B1 _01963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17772_ clknet_leaf_95_clk _00941_ VGND VGND VPWR VPWR count_instr\[43\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15380__S0 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14984_ irq_mask\[4\] _01864_ _01871_ _08335_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_124_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10649__A1 _04419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12150__A_N cpuregs.waddr\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13935_ _07714_ _07721_ VGND VGND VPWR VPWR _07722_ sky130_fd_sc_hd__and2_1
X_16723_ _06989_ cpuregs.regs\[19\]\[22\] _03098_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13415__A _04198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16112__B1_N _02771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16654_ _03064_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__clkbuf_1
X_13866_ _07672_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15132__S0 _01985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15605_ cpuregs.regs\[16\]\[30\] cpuregs.regs\[17\]\[30\] cpuregs.regs\[18\]\[30\]
+ cpuregs.regs\[19\]\[30\] _02221_ _02222_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__mux4_1
X_12817_ _06907_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16585_ _06987_ cpuregs.regs\[18\]\[21\] _03026_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__mux2_1
XANTENNA__09267__A1 _03737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13797_ _05174_ decoded_imm\[30\] VGND VGND VPWR VPWR _07634_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18324_ clknet_leaf_38_clk _01392_ VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15536_ cpuregs.regs\[4\]\[26\] cpuregs.regs\[5\]\[26\] cpuregs.regs\[6\]\[26\] cpuregs.regs\[7\]\[26\]
+ _02046_ _02047_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__mux4_1
XFILLER_0_167_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12748_ _06870_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15435__S1 _01919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18255_ clknet_leaf_26_clk _01326_ VGND VGND VPWR VPWR decoded_imm\[13\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_44_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15467_ cpuregs.regs\[28\]\[22\] cpuregs.regs\[29\]\[22\] cpuregs.regs\[30\]\[22\]
+ cpuregs.regs\[31\]\[22\] _01996_ _01997_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__mux4_1
XFILLER_0_154_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12679_ _06831_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_139_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17206_ clknet_leaf_125_clk _00380_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_14418_ _08084_ _08086_ VGND VGND VPWR VPWR _08087_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18186_ clknet_leaf_43_clk _01257_ VGND VGND VPWR VPWR instr_bge sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15398_ _02238_ _02239_ _03653_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17137_ clknet_leaf_115_clk _00311_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_14349_ _08007_ _08010_ _08019_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__o21ba_1
XANTENNA__15199__S0 _03645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17068_ clknet_leaf_180_clk _00242_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15512__B2 _02037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11129__A2 _05440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12326__A1 _06536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15077__A _03669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11809__S _06348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08910_ _03674_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__buf_4
X_16019_ mem_rdata_q\[22\] _02712_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09890_ net56 _04030_ _04034_ net38 _04423_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08841_ net124 net92 VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08772_ _03535_ _03536_ _03537_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11544__S _06086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15123__S0 _01976_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15579__A1 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09324_ _04058_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09353__S1 _04087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09255_ _03754_ _03744_ _03745_ _03753_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__a22o_2
XFILLER_0_63_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15751__A1 _04979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09186_ _03783_ _03779_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__nor2_2
XFILLER_0_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09430__A1 _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09430__B2 _03226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10591__A3 _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10030_ irq_pending\[17\] _04008_ _04720_ _04748_ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__o22a_1
XANTENNA__10423__S0 _04057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16310__S _02881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11981_ _06442_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_86_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13720_ _07209_ _04979_ _07211_ reg_pc\[24\] _07221_ VGND VGND VPWR VPWR _07563_
+ sky130_fd_sc_hd__a221o_1
X_10932_ _05255_ _05321_ _05597_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__o21a_1
XFILLER_0_169_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13651_ _07191_ _07494_ _07496_ _07497_ VGND VGND VPWR VPWR _07498_ sky130_fd_sc_hd__o31a_1
XFILLER_0_169_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10863_ _05414_ _05424_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14242__A1 reg_next_pc\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12602_ _06790_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__clkbuf_1
X_16370_ _06976_ cpuregs.regs\[16\]\[16\] _02907_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13582_ _07418_ _07422_ VGND VGND VPWR VPWR _07434_ sky130_fd_sc_hd__nand2_1
XANTENNA__15990__A1 _03636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10794_ _05287_ _05311_ _05488_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15321_ net103 _02081_ _02166_ _02167_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_30_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12533_ cpuregs.regs\[2\]\[1\] _06536_ _06752_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__mux2_1
XANTENNA__10594__A _05292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18040_ clknet_leaf_78_clk _00017_ VGND VGND VPWR VPWR irq_pending\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12005__A0 _06320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15252_ _01989_ _02101_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__or2_1
X_12464_ _06096_ cpuregs.regs\[28\]\[1\] _06715_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14203_ reg_pc\[2\] _07906_ _07909_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11415_ _03892_ _05994_ _06021_ _05973_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__a211o_1
XFILLER_0_152_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10567__A0 _04959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15183_ _03692_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__clkbuf_8
X_12395_ cpuregs.regs\[27\]\[1\] _06536_ _06678_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14134_ count_instr\[46\] _07859_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11346_ _03739_ _03853_ _03926_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output263_A net263 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14065_ count_instr\[25\] _07808_ _07790_ VGND VGND VPWR VPWR _07812_ sky130_fd_sc_hd__o21ai_1
X_11277_ _03841_ _05903_ _05904_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_18_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13016_ _07027_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__clkbuf_1
X_10228_ _04940_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__inv_2
XANTENNA__09724__A2 _04429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17824_ clknet_leaf_22_clk _00993_ VGND VGND VPWR VPWR reg_next_pc\[1\] sky130_fd_sc_hd__dfxtp_1
X_10159_ _04010_ _04854_ _04873_ _04150_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17755_ clknet_leaf_89_clk _00924_ VGND VGND VPWR VPWR count_instr\[26\] sky130_fd_sc_hd__dfxtp_1
X_14967_ _07679_ _01859_ _07680_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16706_ _06972_ cpuregs.regs\[19\]\[14\] _03087_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__mux2_1
X_13918_ _03357_ _07704_ _07705_ net134 VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__a22o_1
XANTENNA__09583__S1 _04219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14898_ net224 net257 VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__or2_2
X_17686_ clknet_leaf_119_clk _00855_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16637_ _03055_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__clkbuf_1
X_13849_ cpuregs.regs\[0\]\[21\] VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16568_ _06970_ cpuregs.regs\[18\]\[13\] _03015_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12795__A1 _06582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18307_ clknet_leaf_35_clk _01375_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15519_ cpuregs.regs\[16\]\[25\] cpuregs.regs\[17\]\[25\] cpuregs.regs\[18\]\[25\]
+ cpuregs.regs\[19\]\[25\] _02085_ _02086_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__mux4_1
XANTENNA__13992__B1 _07759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09660__A1 _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16499_ _02982_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09660__B2 _03225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09040_ net45 mem_rdata_q\[20\] _03730_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__mux2_1
XANTENNA__10270__A2 _04962_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18238_ clknet_leaf_23_clk _01309_ VGND VGND VPWR VPWR cpuregs.raddr2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13744__A0 _05174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10558__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18169_ clknet_leaf_23_clk _01240_ VGND VGND VPWR VPWR decoded_imm_j\[10\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_130_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10022__A2 _04104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08702__A net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09942_ count_instr\[15\] _04145_ count_cycle\[15\] _03253_ _04662_ VGND VGND VPWR
+ VPWR _04663_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15592__S0 _01908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09873_ _04010_ _04572_ _04595_ _04150_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__o211a_1
XANTENNA__15249__B1 _02098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08824_ net118 _03583_ _03453_ _03587_ _03589_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__o221a_1
XANTENNA__09533__A _04036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08755_ _03519_ _03520_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_68_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _03450_ _03451_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_136_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14224__A1 reg_pc\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09326__S1 _04060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09307_ net33 net258 _04035_ net40 _04042_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10618__S _05292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09651__A1 _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11303__A _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09238_ _03728_ _03806_ _03808_ _03809_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__a31o_2
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13735__A0 _05013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09403__A1 _04064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09169_ _03849_ _03807_ _03805_ _03850_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16305__S _02870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11200_ _04262_ _05841_ _05827_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10644__S0 _05264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09954__A2 _04642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12180_ cpuregs.regs\[24\]\[9\] _06552_ _06534_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__mux2_1
X_11131_ _05746_ _05395_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__or2b_1
XANTENNA__15583__S0 _01908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11062_ _03452_ _05739_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__nand2_1
X_10013_ cpuregs.regs\[12\]\[17\] cpuregs.regs\[13\]\[17\] cpuregs.regs\[14\]\[17\]
+ cpuregs.regs\[15\]\[17\] _04280_ _04059_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__mux4_1
X_15870_ _02612_ _02613_ _03940_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__and3b_1
XANTENNA__10721__B1 _05215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14821_ count_cycle\[40\] count_cycle\[41\] count_cycle\[42\] _01762_ VGND VGND VPWR
+ VPWR _01768_ sky130_fd_sc_hd__and4_2
XFILLER_0_116_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14752_ _01719_ _08350_ _01720_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__and3b_1
X_17540_ clknet_leaf_10_clk _00709_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11964_ _06433_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13703_ _03631_ _07546_ _07271_ VGND VGND VPWR VPWR _07547_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_158_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ _05292_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__nor2_2
X_17471_ clknet_leaf_177_clk _00640_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14683_ _08315_ _08318_ _08316_ _08309_ VGND VGND VPWR VPWR _08330_ sky130_fd_sc_hd__o211a_1
XANTENNA__09890__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11895_ _06396_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output109_A net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09890__B2 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13634_ _07482_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16422_ _02941_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10846_ _05234_ _05267_ _05270_ _05273_ _05413_ _05414_ VGND VGND VPWR VPWR _05538_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__15963__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16353_ _06959_ cpuregs.regs\[16\]\[8\] _02896_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13565_ net72 decoded_imm\[14\] VGND VGND VPWR VPWR _07418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10777_ _03511_ _05440_ _05357_ _03512_ _05472_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__o221a_1
XANTENNA__10788__A0 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09642__A1 _04328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15304_ cpuregs.regs\[8\]\[13\] cpuregs.regs\[9\]\[13\] cpuregs.regs\[10\]\[13\]
+ cpuregs.regs\[11\]\[13\] _02013_ _02014_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_171_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12516_ _06304_ cpuregs.regs\[28\]\[26\] _06737_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16284_ _06959_ cpuregs.regs\[15\]\[8\] _02859_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13496_ _07352_ _07353_ VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15235_ _01919_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__buf_8
X_18023_ clknet_leaf_104_clk _00030_ VGND VGND VPWR VPWR irq_pending\[7\] sky130_fd_sc_hd__dfxtp_1
X_12447_ cpuregs.regs\[27\]\[26\] _06588_ _06700_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__mux2_1
XANTENNA__12743__S _06863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14524__A _07943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output90_A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15166_ _03639_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__buf_6
XFILLER_0_151_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08522__A _03301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12378_ cpuregs.regs\[26\]\[26\] _06588_ _06663_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_26_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14117_ count_instr\[41\] _07845_ _07847_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__a21oi_1
X_11329_ reg_next_pc\[29\] _05928_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16140__A1 net256 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15097_ _03388_ _01955_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__nor2_1
X_14048_ _07799_ _07800_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__nor2_1
XANTENNA__12979__A _06342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15326__S0 _01982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17807_ clknet_leaf_61_clk _00976_ VGND VGND VPWR VPWR reg_pc\[15\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__15074__B _03301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15999_ decoded_rd\[4\] _05974_ _03763_ _02706_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_173_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08540_ decoder_trigger do_waitirq instr_waitirq VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__o21a_2
XFILLER_0_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17738_ clknet_leaf_96_clk _00907_ VGND VGND VPWR VPWR count_instr\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08471_ instr_sltu instr_slt instr_sltiu instr_slti VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__or4_2
XFILLER_0_49_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17669_ clknet_leaf_19_clk _00838_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12768__A1 _06554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13322__B _03274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09023_ _03782_ _03784_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12653__S _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16125__S _02771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09397__B1 _04080_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11777__B reg_pc\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16131__A1 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10951__B1 _05334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14142__B1 _07834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09925_ _04483_ _04645_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09856_ _04487_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__buf_8
X_08807_ net111 VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09787_ _04273_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__buf_8
XANTENNA__16795__S _03138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14445__A1 reg_next_pc\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14445__B2 _08033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08738_ _03502_ _03503_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__nor2_2
XANTENNA_105 _05591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14996__A2 _04022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10467__C1 _03302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_138 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08669_ net122 net90 VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__nor2_1
XANTENNA_149 net203 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09872__A1 _04168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12828__S _06906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10700_ _05244_ _05399_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__nand2_1
X_11680_ _06234_ _06118_ _06235_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__and3b_1
XFILLER_0_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10631_ _05272_ _05274_ _05309_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10234__A2 _04945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13350_ _07216_ VGND VGND VPWR VPWR _07217_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10562_ _05235_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__buf_4
XFILLER_0_107_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12301_ cpuregs.regs\[25\]\[22\] _06580_ _06626_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13281_ _06968_ cpuregs.regs\[5\]\[12\] _07165_ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__mux2_1
XANTENNA__10872__A _05287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10493_ _04328_ _05197_ _04237_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15020_ irq_mask\[19\] _01880_ _01892_ _01891_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12232_ _06303_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_131_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10537__A3 _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12163_ _06541_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15556__S0 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11114_ _03438_ _05787_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__xnor2_1
X_16971_ clknet_leaf_153_clk _00145_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_12094_ _06502_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15175__A _02012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11907__S _06398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11045_ _03456_ _05722_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__or2_1
X_15922_ instr_sll _02617_ _02620_ _02653_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__a22o_1
XANTENNA__15308__S0 _02022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09786__S1 _04317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09173__A _03781_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18641_ clknet_leaf_99_clk _01701_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_129_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ mem_rdata_q\[13\] VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_output226_A net226 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14804_ count_cycle\[36\] _01752_ _01723_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__o21ai_1
X_18572_ clknet_leaf_110_clk _01637_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_15784_ _03630_ is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__or2b_1
X_12996_ cpuregs.regs\[3\]\[6\] _06546_ _07010_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17523_ clknet_leaf_154_clk _00692_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14735_ count_cycle\[15\] _08362_ _07877_ VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__o21ai_1
X_11947_ _06078_ cpuregs.regs\[21\]\[0\] _06424_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09863__A1 _04320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ clknet_leaf_137_clk _00623_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14666_ reg_next_pc\[29\] _07948_ _08305_ _08314_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11878_ _06078_ cpuregs.regs\[20\]\[0\] _06387_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13617_ _04708_ _05260_ _07425_ _07238_ VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__o211a_1
X_16405_ _06941_ cpuregs.regs\[29\]\[0\] _02932_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__mux2_1
X_10829_ _03501_ _05220_ _05301_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09615__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14597_ reg_next_pc\[23\] _07903_ _08250_ _03378_ _08251_ VGND VGND VPWR VPWR _08252_
+ sky130_fd_sc_hd__a221o_1
X_17385_ clknet_leaf_183_clk _00554_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09615__B2 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13548_ _07391_ _07392_ _07401_ _07402_ VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__a22o_1
X_16336_ _02895_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08951__S _03713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16267_ _02858_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__buf_6
X_13479_ _07338_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18006_ clknet_leaf_80_clk _01143_ VGND VGND VPWR VPWR irq_mask\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15218_ _01991_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__buf_8
XFILLER_0_11_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11597__B reg_pc\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16198_ net298 _01822_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11186__A0 reg_next_pc\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16113__A1 _05829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15149_ _03675_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__buf_6
XANTENNA__10084__S1 _04283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16113__B2 net193 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14124__B1 _07834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09710_ _04435_ _04436_ _04321_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__mux2_1
XANTENNA__11817__S _06348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12686__A0 _06166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09641_ _04367_ _04368_ _04369_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09572_ cpuregs.regs\[16\]\[5\] cpuregs.regs\[17\]\[5\] cpuregs.regs\[18\]\[5\] cpuregs.regs\[19\]\[5\]
+ _04217_ _04219_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08523_ _03302_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14429__A instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13650__A2 _04842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08454_ mem_do_prefetch _03237_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15927__A1 _02625_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15155__A2 _02009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09006_ _03743_ _03747_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__or2_2
XFILLER_0_104_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08593__A1 _03277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08593__B2 _03298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09908_ _04082_ _04617_ _04621_ _04625_ _04629_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__a32o_1
X_09839_ irq_mask\[12\] _04308_ timer\[12\] instr_timer _04026_ VGND VGND VPWR VPWR
+ _04563_ sky130_fd_sc_hd__a221o_1
X_12850_ _06924_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09721__A _04308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11801_ _06343_ cpuregs.regs\[10\]\[31\] _06085_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11101__A0 _05143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12781_ _06887_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12558__S _06763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10867__A _05288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09845__B2 _03225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14339__A _07998_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14520_ _08176_ _08179_ VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__nand2_1
X_11732_ _06282_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_25_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14451_ _08115_ _08116_ VGND VGND VPWR VPWR _08117_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11663_ reg_out\[16\] alu_out_q\[16\] _06067_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__mux2_1
XANTENNA__10078__S _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13402_ _03399_ _07265_ VGND VGND VPWR VPWR _07266_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10614_ _05263_ _05205_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__or2b_1
X_17170_ clknet_leaf_114_clk _00344_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14382_ _08052_ _08053_ VGND VGND VPWR VPWR _08054_ sky130_fd_sc_hd__nand2_1
X_11594_ reg_out\[9\] alu_out_q\[9\] _06067_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16121_ net263 _05324_ _02771_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13333_ cpuregs.regs\[4\]\[0\] cpuregs.regs\[5\]\[0\] cpuregs.regs\[6\]\[0\] cpuregs.regs\[7\]\[0\]
+ _04758_ _04759_ VGND VGND VPWR VPWR _07200_ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10545_ _05248_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_130_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_130_clk sky130_fd_sc_hd__clkbuf_2
X_16052_ _03402_ decoded_imm_j\[14\] _03403_ _03940_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__a22o_1
X_13264_ _06951_ cpuregs.regs\[5\]\[4\] _07154_ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10476_ _05146_ _05178_ _05179_ _04156_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__a31o_1
XANTENNA__11168__B1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15003_ _04561_ _01869_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output176_A net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12215_ cpuregs.regs\[24\]\[20\] _06575_ _06576_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13195_ _07122_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08584__A1 _03340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12146_ _06529_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_166_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08800__A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13418__A _07209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10930__A3 _04611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12668__A0 _06078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16954_ clknet_leaf_190_clk _00128_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12077_ _06336_ cpuregs.regs\[22\]\[30\] _06459_ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__mux2_1
XANTENNA__09759__S1 _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11028_ _03468_ _03471_ _03467_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__a21boi_1
X_15905_ instr_sw _02635_ _02639_ is_sb_sh_sw VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__a22o_1
X_16885_ clknet_leaf_41_clk _00081_ VGND VGND VPWR VPWR mem_wordsize\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12745__B_N _06081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18624_ clknet_leaf_1_clk _01684_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_15836_ _08232_ _05987_ _03756_ _02587_ _02596_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__a221o_1
XANTENNA__15082__A1 _03709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09631__A _03518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18555_ clknet_leaf_182_clk _01620_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_15767_ timer\[28\] _02560_ _02562_ _02488_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__a211o_1
XANTENNA__09836__A1 _04328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12468__S _06715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12979_ _06342_ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__buf_2
X_17506_ clknet_leaf_188_clk _00675_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10446__A2 _04012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14718_ _08353_ _08354_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18486_ clknet_leaf_189_clk _01551_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09931__S1 _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15698_ _07371_ _02486_ _02510_ _02511_ _06026_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__o221a_1
XFILLER_0_87_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17437_ clknet_leaf_114_clk _00606_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14649_ _03293_ _07967_ _07995_ _07904_ reg_next_pc\[28\] VGND VGND VPWR VPWR _08299_
+ sky130_fd_sc_hd__a32o_1
XANTENNA_16 _03351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_27 _04483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_38 _05864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 decoded_imm\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17368_ clknet_leaf_164_clk _00537_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13600__B _05227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16319_ _02886_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_121_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_121_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__08811__A2 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17299_ clknet_leaf_166_clk _00473_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput101 net101 VGND VGND VPWR VPWR cpi_rs2[11] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09447__S0 _04055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14896__A1 _05205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput112 net112 VGND VGND VPWR VPWR cpi_rs2[21] sky130_fd_sc_hd__buf_1
XFILLER_0_141_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput123 net123 VGND VGND VPWR VPWR cpi_rs2[31] sky130_fd_sc_hd__buf_1
Xoutput134 net134 VGND VGND VPWR VPWR eoi[12] sky130_fd_sc_hd__clkbuf_1
XANTENNA__12931__S _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput145 net145 VGND VGND VPWR VPWR eoi[22] sky130_fd_sc_hd__buf_1
XANTENNA__14712__A _03304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput156 net156 VGND VGND VPWR VPWR eoi[3] sky130_fd_sc_hd__buf_1
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput167 net167 VGND VGND VPWR VPWR mem_addr[14] sky130_fd_sc_hd__clkbuf_1
Xoutput178 net178 VGND VGND VPWR VPWR mem_addr[25] sky130_fd_sc_hd__clkbuf_1
XANTENNA__08710__A net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput189 net189 VGND VGND VPWR VPWR mem_addr[6] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_54_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12659__A0 _06328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13328__A _04272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12232__A _06303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09524__B1 _04008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_188_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_188_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09624_ cpu_state\[3\] _04351_ _04353_ irq_pending\[6\] _04266_ VGND VGND VPWR VPWR
+ _04354_ sky130_fd_sc_hd__a32o_1
XANTENNA__09541__A _04054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09555_ cpuregs.regs\[8\]\[5\] cpuregs.regs\[9\]\[5\] cpuregs.regs\[10\]\[5\] cpuregs.regs\[11\]\[5\]
+ _04282_ _04285_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__mux4_1
XANTENNA__12378__S _06663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08506_ _03281_ _03285_ _03288_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09922__S1 _04470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09486_ _04124_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__buf_4
XFILLER_0_93_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08437_ _03187_ _03215_ _03217_ _03222_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13387__A1 _04198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_112_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_112_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__10070__B1 _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13002__S _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10330_ count_instr\[58\] _04015_ instr_rdcycleh count_cycle\[58\] VGND VGND VPWR
+ VPWR _05040_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12841__S _06917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10261_ _04971_ _04972_ _04222_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12000_ _06452_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10192_ _04900_ _04902_ _04905_ _04052_ _04095_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__a221o_1
XANTENNA__15836__B1 _03756_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13951_ _03320_ _07727_ _07728_ net145 VGND VGND VPWR VPWR _07733_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_179_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_179_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__10125__A1 _04272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12902_ _06140_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__buf_2
XFILLER_0_88_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13882_ _03351_ _07678_ _07682_ net142 VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__a22o_1
X_16670_ _03072_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10220__S1 _04470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12833_ _06915_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__clkbuf_1
X_15621_ cpuregs.regs\[8\]\[31\] cpuregs.regs\[9\]\[31\] cpuregs.regs\[10\]\[31\]
+ cpuregs.regs\[11\]\[31\] _03645_ _01991_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__mux4_1
XANTENNA__12288__S _06615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18340_ clknet_leaf_38_clk _01408_ VGND VGND VPWR VPWR mem_16bit_buffer\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12822__A0 _06114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12764_ _06878_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15552_ cpuregs.regs\[16\]\[27\] cpuregs.regs\[17\]\[27\] cpuregs.regs\[18\]\[27\]
+ cpuregs.regs\[19\]\[27\] _02030_ _02031_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__mux4_1
XFILLER_0_83_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14503_ decoded_imm_j\[16\] _07941_ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__nor2_1
X_11715_ _06267_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15900__B _02613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15483_ cpuregs.regs\[16\]\[23\] cpuregs.regs\[17\]\[23\] cpuregs.regs\[18\]\[23\]
+ cpuregs.regs\[19\]\[23\] _02046_ _02047_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__mux4_1
X_18271_ clknet_leaf_25_clk _01342_ VGND VGND VPWR VPWR decoded_imm\[29\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12695_ _06201_ cpuregs.regs\[12\]\[13\] _06836_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11920__S _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09597__S _04223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17222_ clknet_leaf_137_clk _00396_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11646_ _03409_ _03353_ _06066_ _06205_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__a22o_1
X_14434_ _07899_ _07928_ _08050_ _08101_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14516__B _07943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 irq[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput25 irq[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17153_ clknet_leaf_184_clk _00327_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_14365_ decoded_imm_j\[5\] _07917_ VGND VGND VPWR VPWR _08038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 mem_rdata[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_103_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_103_clk sky130_fd_sc_hd__clkbuf_2
X_11577_ _06072_ _03349_ _06098_ _06143_ _06118_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__a221o_1
XANTENNA__10287__S1 _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput47 mem_rdata[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
XFILLER_0_135_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08514__B net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput58 mem_rdata[3] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_1
X_13316_ _07003_ cpuregs.regs\[5\]\[29\] _07176_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16104_ _06023_ _02764_ _02765_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10600__A2 _05286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10528_ _05231_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17084_ clknet_leaf_3_clk _00258_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_14296_ irq_pending\[20\] irq_pending\[21\] irq_pending\[22\] irq_pending\[23\] VGND
+ VGND VPWR VPWR _07973_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13247_ _07149_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__clkbuf_1
X_16035_ decoded_imm\[6\] _02711_ _02729_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__o21a_1
X_10459_ cpuregs.regs\[8\]\[30\] cpuregs.regs\[9\]\[30\] cpuregs.regs\[10\]\[30\]
+ cpuregs.regs\[11\]\[30\] _04280_ _04059_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__mux4_1
XANTENNA__12751__S _06869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13178_ _07001_ cpuregs.regs\[4\]\[28\] _07104_ VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__mux2_1
XANTENNA__08530__A _03237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15827__B1 _03891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12129_ _06274_ cpuregs.regs\[23\]\[22\] _06518_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__mux2_1
X_17986_ clknet_leaf_103_clk _01123_ VGND VGND VPWR VPWR irq_mask\[2\] sky130_fd_sc_hd__dfxtp_4
XANTENNA__09506__B1 _04237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16937_ clknet_leaf_164_clk _00118_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09601__S0 _04329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_56 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10211__S1 _04513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16868_ _03178_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__clkbuf_1
X_18607_ clknet_leaf_164_clk _01672_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_15819_ _03867_ _06016_ _02586_ _04000_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16799_ _06582_ cpuregs.regs\[13\]\[23\] _03138_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__mux2_1
X_09340_ cpuregs.regs\[20\]\[1\] cpuregs.regs\[21\]\[1\] cpuregs.regs\[22\]\[1\] cpuregs.regs\[23\]\[1\]
+ _04072_ _04074_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18538_ clknet_leaf_98_clk _01603_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09904__S1 _04276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09271_ _04007_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18469_ clknet_leaf_132_clk _01534_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09690__C1 _04149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11830__S _06359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08705__A net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09993__B1 _04202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15530__A2 _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16133__S _02771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08986_ _03747_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16243__A0 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09607_ irq_mask\[6\] _04021_ timer\[6\] _04187_ _04188_ VGND VGND VPWR VPWR _04337_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__15597__A2 _01906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09538_ count_instr\[5\] _04011_ _04017_ count_cycle\[37\] VGND VGND VPWR VPWR _04269_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_955 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09469_ _04048_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15720__B _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11740__S _06258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11500_ _03195_ _06065_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13521__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14557__B1 _08055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12480_ _06166_ cpuregs.regs\[28\]\[9\] _06715_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10864__B _05367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08615__A is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11431_ irq_mask\[5\] _06030_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__or2_1
XFILLER_0_163_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14150_ _07871_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11362_ _03228_ _03633_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__nand2_2
XFILLER_0_81_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13101_ _07072_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10313_ _05021_ _05022_ _04077_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14081_ _07821_ _07815_ _07822_ VGND VGND VPWR VPWR _07823_ sky130_fd_sc_hd__and3b_1
XFILLER_0_132_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11293_ _05917_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_2
X_13032_ cpuregs.regs\[3\]\[23\] _06582_ _07032_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__mux2_1
X_10244_ reg_pc\[24\] decoded_imm\[24\] VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_163_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17840_ clknet_leaf_61_clk _01009_ VGND VGND VPWR VPWR reg_next_pc\[17\] sky130_fd_sc_hd__dfxtp_1
X_10175_ count_instr\[54\] _04015_ _04017_ count_cycle\[54\] VGND VGND VPWR VPWR _04889_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15285__A1 decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17771_ clknet_leaf_95_clk _00940_ VGND VGND VPWR VPWR count_instr\[42\] sky130_fd_sc_hd__dfxtp_1
X_14983_ _04240_ _01869_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__nor2_1
XANTENNA__15380__S1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11915__S _06398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15183__A _03692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16722_ _03100_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__clkbuf_1
X_13934_ _03348_ _07704_ _07705_ net139 VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__a22o_1
XANTENNA__10649__A2 _03518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16653_ cpuregs.regs\[1\]\[21\] _06265_ _03062_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__mux2_1
X_13865_ cpuregs.regs\[0\]\[29\] VGND VGND VPWR VPWR _07672_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15132__S1 _01986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15911__A _02611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15604_ cpuregs.regs\[20\]\[30\] cpuregs.regs\[21\]\[30\] cpuregs.regs\[22\]\[30\]
+ cpuregs.regs\[23\]\[30\] _02221_ _02222_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14796__B1 _01717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12816_ _06078_ cpuregs.regs\[6\]\[0\] _06906_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__mux2_1
X_16584_ _03027_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__clkbuf_1
X_13796_ _05174_ decoded_imm\[30\] VGND VGND VPWR VPWR _07633_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18323_ clknet_leaf_38_clk _01391_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15535_ _03719_ _02368_ _00068_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16537__A1 _06598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12747_ cpuregs.regs\[9\]\[0\] _06531_ _06869_ VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18254_ clknet_leaf_26_clk _01325_ VGND VGND VPWR VPWR decoded_imm\[12\] sky130_fd_sc_hd__dfxtp_4
X_15466_ _02300_ _02301_ _02302_ _02303_ _02111_ _02004_ VGND VGND VPWR VPWR _02304_
+ sky130_fd_sc_hd__mux4_1
X_12678_ _06132_ cpuregs.regs\[12\]\[5\] _06825_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08525__A _03304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_578 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17205_ clknet_leaf_115_clk _00379_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11629_ _03409_ _03357_ _06066_ _06190_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14417_ _08060_ _08064_ _08085_ _08073_ VGND VGND VPWR VPWR _08086_ sky130_fd_sc_hd__a31o_1
X_18185_ clknet_leaf_43_clk _01256_ VGND VGND VPWR VPWR instr_blt sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15397_ cpuregs.regs\[0\]\[18\] cpuregs.regs\[1\]\[18\] cpuregs.regs\[2\]\[18\] cpuregs.regs\[3\]\[18\]
+ _02046_ _02047_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17136_ clknet_leaf_110_clk _00310_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14348_ reg_next_pc\[3\] _07948_ _08015_ _08022_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15199__S1 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17067_ clknet_leaf_178_clk _00241_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_14279_ reg_pc\[25\] _07906_ _07962_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13523__A1 _04466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09356__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16018_ decoded_imm\[1\] _02711_ _02714_ _02717_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11534__A0 _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10337__B2 _05046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09822__S0 _04085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08840_ _03530_ net92 VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09790__S _04321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08771_ net110 net78 VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__or2b_1
XANTENNA__13287__A0 _06974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17969_ clknet_leaf_4_clk _01106_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dfxtp_1
XANTENNA__15805__B _03763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13604__A1_N _03387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11825__S _06348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16225__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15123__S1 _01977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09323_ _00070_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14437__A decoded_imm_j\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09254_ _03838_ _03988_ _03993_ _03888_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09185_ mem_rdata_q\[13\] _03747_ _03227_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13762__A1 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10576__A1 _05255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09430__A2 _04160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10576__B2 _03630_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09718__B1 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10423__S1 _04060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14900__A _01823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15267__B2 _02037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08969_ net36 mem_rdata_q\[12\] _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__mux2_1
XANTENNA__15207__S _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11980_ _06224_ cpuregs.regs\[21\]\[16\] _06435_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10187__S0 _04280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10931_ _05617_ _05561_ _05395_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__mux2_1
XANTENNA__11036__A _05287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10862_ _03496_ _05552_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__xor2_1
X_13650_ _07281_ _04842_ _07282_ reg_pc\[20\] _07283_ VGND VGND VPWR VPWR _07497_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _06096_ cpuregs.regs\[30\]\[1\] _06788_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11056__A2 _05357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13581_ net73 decoded_imm\[15\] VGND VGND VPWR VPWR _07433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16519__A1 _06580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10793_ _03530_ _05291_ _05228_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12566__S _06763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15990__A2 _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15320_ decoded_imm\[13\] _02009_ _01963_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__a21o_1
X_12532_ _06753_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15877__S _03635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15251_ cpuregs.regs\[8\]\[10\] cpuregs.regs\[9\]\[10\] cpuregs.regs\[10\]\[10\]
+ cpuregs.regs\[11\]\[10\] _02013_ _02014_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__mux4_1
X_12463_ _06716_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10016__B1 _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14202_ _06860_ _07908_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__nor2_1
X_11414_ _03215_ _03918_ _06002_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__and3_1
X_15182_ _02034_ _02035_ _02002_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12394_ _06679_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10567__A1 _05013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10111__S0 _04275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14133_ _07857_ _07855_ _07859_ _07775_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_134_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11345_ _03228_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_134_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15050__S0 _01908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14064_ count_instr\[25\] count_instr\[24\] count_instr\[23\] _07805_ VGND VGND VPWR
+ VPWR _07811_ sky130_fd_sc_hd__and4_2
XANTENNA__09176__A _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11276_ _05896_ _05899_ _05902_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__and3_1
XANTENNA_output256_A net256 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11516__B1 _03351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13015_ cpuregs.regs\[3\]\[15\] _06565_ _07021_ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__mux2_1
XANTENNA__09185__A1 _03747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10227_ _04927_ _04931_ _04939_ _04100_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__a211o_2
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15906__A mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17823_ clknet_leaf_68_clk _00992_ VGND VGND VPWR VPWR reg_pc\[31\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10158_ _04168_ _04871_ _04872_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_131_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17754_ clknet_leaf_85_clk _00923_ VGND VGND VPWR VPWR count_instr\[25\] sky130_fd_sc_hd__dfxtp_1
X_10089_ _04805_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__inv_2
X_14966_ _06186_ _03298_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10178__S0 _04281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16705_ _03091_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__clkbuf_1
X_13917_ _07709_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11295__A2 _05915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17685_ clknet_leaf_97_clk _00854_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14897_ _03196_ net299 VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__nor2_2
X_16636_ cpuregs.regs\[1\]\[13\] _06200_ _03051_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_146_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13848_ _07663_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16567_ _03018_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12476__S _06715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13779_ _03275_ _07611_ _07612_ _07616_ _07617_ VGND VGND VPWR VPWR _07618_ sky130_fd_sc_hd__a32o_1
XANTENNA__14257__A _07947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13161__A _07081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18306_ clknet_leaf_35_clk _01374_ VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dfxtp_1
X_15518_ cpuregs.regs\[20\]\[25\] cpuregs.regs\[21\]\[25\] cpuregs.regs\[22\]\[25\]
+ cpuregs.regs\[23\]\[25\] _01973_ _01974_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_44_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16498_ cpuregs.regs\[17\]\[12\] _06559_ _02979_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__mux2_1
XANTENNA__09660__A2 _04360_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18237_ clknet_leaf_23_clk _01308_ VGND VGND VPWR VPWR cpuregs.raddr2\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_1001 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_61_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15449_ cpuregs.regs\[8\]\[21\] cpuregs.regs\[9\]\[21\] cpuregs.regs\[10\]\[21\]
+ cpuregs.regs\[11\]\[21\] _02085_ _02086_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16472__A _02967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09785__S _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13744__A1 _04913_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09948__B1 _04668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18168_ clknet_leaf_23_clk _01239_ VGND VGND VPWR VPWR decoded_imm_j\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10558__A1 _04744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09412__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14704__B _07815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17119_ clknet_leaf_179_clk _00293_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08620__B1 _03394_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18099_ clknet_leaf_91_clk _01203_ VGND VGND VPWR VPWR timer\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08702__B net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13100__S _07068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09941_ count_instr\[47\] _04015_ _04017_ count_cycle\[47\] VGND VGND VPWR VPWR _04662_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15592__S1 _01909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10025__A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09872_ _04168_ _04593_ _04594_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__a21o_1
XANTENNA__16411__S _02932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15249__A1 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08823_ _03449_ _03588_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__nand2_1
X_08754_ net127 net95 VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ net117 net85 VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11286__A2 _05906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14224__A2 _07906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12386__S _06640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10695__A _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09306_ _04037_ _04038_ _04041_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09237_ mem_rdata_q\[27\] _03977_ _03227_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15185__B1 _02027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_863 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15280__S0 _01999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14932__A0 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09168_ _03908_ _03919_ _03917_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__o21a_1
XFILLER_0_161_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09099_ _03835_ _03858_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11130_ _05205_ _05174_ _05143_ _05086_ _05324_ _05286_ VGND VGND VPWR VPWR _05803_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15583__S1 _01909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11061_ _05736_ _05738_ _05322_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ _04729_ _04730_ _04121_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__mux2_1
X_14820_ _01767_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14751_ count_cycle\[19\] _01715_ count_cycle\[20\] VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__a21o_1
X_11963_ _06157_ cpuregs.regs\[21\]\[8\] _06424_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_2
X_13702_ _07544_ _07545_ VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10914_ instr_sll instr_slli _05226_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__o21ai_2
X_17470_ clknet_leaf_128_clk _00639_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11894_ _06157_ cpuregs.regs\[20\]\[8\] _06387_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__mux2_1
X_14682_ _03195_ _03363_ _07971_ _08050_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__o31a_1
XFILLER_0_168_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16421_ _06959_ cpuregs.regs\[29\]\[8\] _02932_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__mux2_1
X_10845_ _03499_ _05535_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__or2_1
X_13633_ _04754_ _07481_ _07374_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16352_ _02904_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13564_ _07417_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__clkbuf_1
X_10776_ _03509_ _05301_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__nand2_1
XANTENNA__10788__A1 _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15303_ cpuregs.regs\[12\]\[13\] cpuregs.regs\[13\]\[13\] cpuregs.regs\[14\]\[13\]
+ cpuregs.regs\[15\]\[13\] _01970_ _01971_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11213__B _05848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12515_ _06743_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_171_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13495_ _03510_ decoded_imm\[8\] _07347_ VGND VGND VPWR VPWR _07353_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16283_ _02867_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15271__S0 _01970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18022_ clknet_leaf_105_clk _00029_ VGND VGND VPWR VPWR irq_pending\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_124_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12446_ _06706_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__clkbuf_1
X_15234_ _01918_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__buf_12
XFILLER_0_125_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08803__A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09618__B decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15165_ _01989_ _02011_ _02016_ _02018_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__o211a_1
X_12377_ _06669_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output83_A net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11328_ _05938_ _05943_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__and2_1
X_14116_ count_instr\[41\] _07845_ _07675_ VGND VGND VPWR VPWR _07847_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15096_ _03679_ _01954_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__nand2_2
XFILLER_0_157_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09158__A1 _03878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14047_ count_instr\[19\] _07796_ _07790_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__o21ai_1
X_11259_ _05888_ _05889_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15326__S1 _03639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17806_ clknet_leaf_62_clk _00975_ VGND VGND VPWR VPWR reg_pc\[14\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_2_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13337__S0 _04579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15998_ decoded_rd\[3\] _05987_ _03892_ _02706_ _02710_ VGND VGND VPWR VPWR _01301_
+ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_167_Right_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17737_ clknet_leaf_96_clk _00906_ VGND VGND VPWR VPWR count_instr\[8\] sky130_fd_sc_hd__dfxtp_1
X_14949_ net209 net178 _01846_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_74_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10476__B1 _04156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08470_ _03252_ instr_rdcycle _03253_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__or3b_4
X_17668_ clknet_leaf_2_clk _00837_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16619_ cpuregs.regs\[1\]\[5\] _06131_ _03040_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17599_ clknet_leaf_163_clk _00768_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09633__A2 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10323__S0 _04055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12934__S _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15262__S0 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09022_ _03783_ _03213_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09397__A1 _04052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09528__B decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14544__B1_N _07972_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12235__A _06311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09149__A1 _03763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10951__B2 _05254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09924_ _04643_ _04644_ _04065_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09544__A _04274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09855_ cpuregs.regs\[28\]\[13\] cpuregs.regs\[29\]\[13\] cpuregs.regs\[30\]\[13\]
+ cpuregs.regs\[31\]\[13\] _04512_ _04513_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__mux4_1
X_08806_ net109 _03475_ _03489_ _03564_ _03571_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__o221a_1
XFILLER_0_147_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09786_ cpuregs.regs\[4\]\[11\] cpuregs.regs\[5\]\[11\] cpuregs.regs\[6\]\[11\] cpuregs.regs\[7\]\[11\]
+ _04274_ _04317_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__mux4_1
XANTENNA__15642__A1 is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14445__A2 _07947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15642__B2 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08737_ net101 net69 VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_106 _05929_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_65_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__14996__A3 _04447_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_128 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08668_ _03432_ _03433_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__nand2_2
XANTENNA_139 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09872__A2 _04593_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12208__A1 _06571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08599_ _03363_ _03293_ _03376_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__and3b_1
XFILLER_0_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13005__S _07021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10630_ _05329_ _05330_ _05331_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__mux2_1
XANTENNA__11314__A _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10561_ _04754_ _04810_ _05264_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16316__S _02881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12300_ _06628_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14905__A0 net218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13280_ _07167_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__clkbuf_1
X_10492_ _05195_ _05196_ _04222_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12231_ _06587_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12162_ cpuregs.regs\[24\]\[3\] _06540_ _06534_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10942__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15556__S1 _01997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11113_ _05363_ _05783_ _05786_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15330__B1 _02017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16970_ clknet_leaf_140_clk _00144_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12093_ _06132_ cpuregs.regs\[23\]\[5\] _06496_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_15_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11044_ _03456_ _05722_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__nand2_1
XANTENNA__09454__A instr_timer VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15921_ is_alu_reg_reg _02615_ _02656_ _02616_ _05517_ VGND VGND VPWR VPWR _01278_
+ sky130_fd_sc_hd__a32o_1
XANTENNA__15308__S1 _02023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18640_ clknet_leaf_99_clk _01700_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15852_ mem_rdata_q\[12\] VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15633__A1 mem_do_prefetch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14803_ count_cycle\[34\] count_cycle\[35\] count_cycle\[36\] _01748_ VGND VGND VPWR
+ VPWR _01756_ sky130_fd_sc_hd__and4_2
X_18571_ clknet_leaf_122_clk _01636_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12447__A1 _06588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output121_A net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15783_ _03298_ _04006_ _03389_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_2
X_12995_ _07016_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output219_A net219 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17522_ clknet_leaf_146_clk _00691_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_14734_ count_cycle\[13\] count_cycle\[14\] count_cycle\[15\] _08359_ VGND VGND VPWR
+ VPWR _08365_ sky130_fd_sc_hd__and4_2
X_11946_ _06423_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__buf_6
XFILLER_0_52_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ clknet_leaf_148_clk _00622_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_14665_ _08012_ _08312_ _08313_ _08120_ VGND VGND VPWR VPWR _08314_ sky130_fd_sc_hd__o2bb2a_1
X_11877_ _06386_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__buf_6
XFILLER_0_157_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16404_ _02931_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__buf_6
X_13616_ _04602_ _07236_ _07465_ _07217_ VGND VGND VPWR VPWR _07466_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10828_ _03504_ _05520_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__xor2_2
X_17384_ clknet_leaf_172_clk _00553_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09615__A2 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14596_ _03293_ _07958_ _07992_ VGND VGND VPWR VPWR _08251_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16335_ _06383_ _02894_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__nand2_4
X_13547_ _07394_ _07397_ _07400_ _03631_ VGND VGND VPWR VPWR _07402_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_15_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10759_ _05383_ _05423_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15244__S0 _02074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16266_ _06346_ _06823_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__nand2_2
X_13478_ _04360_ _07337_ _07225_ VGND VGND VPWR VPWR _07338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18005_ clknet_leaf_79_clk _01142_ VGND VGND VPWR VPWR irq_mask\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15217_ _01936_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__buf_8
XFILLER_0_2_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12429_ _06697_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__clkbuf_1
X_16197_ net257 net261 _01822_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15148_ _01998_ _02001_ _02002_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15321__B1 _02166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15079_ cpuregs.regs\[8\]\[1\] cpuregs.regs\[9\]\[1\] cpuregs.regs\[10\]\[1\] cpuregs.regs\[11\]\[1\]
+ _01936_ _01937_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09640_ _00071_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__buf_6
XANTENNA__16821__A0 _06536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09571_ cpuregs.regs\[20\]\[5\] cpuregs.regs\[21\]\[5\] cpuregs.regs\[22\]\[5\] cpuregs.regs\[23\]\[5\]
+ _04217_ _04219_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__mux4_1
XANTENNA__09839__C1 _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_47_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_2
X_08522_ _03301_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09811__B decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14429__B _07754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08453_ _03236_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__buf_2
XFILLER_0_93_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10449__S _04065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15483__S0 _02046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_830 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13987__C _07755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09005_ _03727_ _03764_ _03765_ _03766_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__a31o_4
XFILLER_0_170_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11177__A1 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09274__A instr_rdinstr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14666__A2 _07948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09907_ _04328_ _04628_ _04081_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_45_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09838_ _04561_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09769_ irq_mask\[10\] _04021_ timer\[10\] _04023_ _04188_ VGND VGND VPWR VPWR _04495_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__12839__S _06917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_2
X_11800_ _06342_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__buf_2
XANTENNA__11101__A1 _05086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12780_ cpuregs.regs\[9\]\[16\] _06567_ _06880_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09845__A2 _04566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _06281_ cpuregs.regs\[10\]\[23\] _06258_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16040__B2 mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09058__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14450_ _08106_ _08108_ _08104_ VGND VGND VPWR VPWR _08116_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11662_ _06218_ _06219_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_54_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13401_ _04160_ _04251_ _05257_ VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__mux2_1
X_10613_ instr_sra instr_srai _05205_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_37_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11593_ _06158_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__clkbuf_1
X_14381_ decoded_imm_j\[6\] _07919_ VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10612__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16120_ mem_state\[1\] _02775_ _02777_ _02771_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10544_ _05246_ _05247_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__or2_1
X_13332_ _04215_ _07198_ _04225_ VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16051_ decoded_imm\[13\] _02720_ _02736_ _02738_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__o22a_1
XFILLER_0_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10475_ _05146_ _05178_ _05179_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__a21oi_1
X_13263_ _07158_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11168__A1 _04038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11168__B2 _03297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15002_ irq_mask\[11\] _01880_ _01882_ _01876_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12214_ _06533_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__clkbuf_8
X_13194_ _06949_ cpuregs.regs\[8\]\[3\] _07118_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__mux2_1
XANTENNA__09781__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08584__A2 _03361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12145_ _06336_ cpuregs.regs\[23\]\[30\] _06495_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__mux2_1
XANTENNA__09781__B2 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_63_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12076_ _06492_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__clkbuf_1
X_16953_ clknet_leaf_17_clk _00127_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11027_ _05599_ _05601_ _05701_ _05704_ _05706_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__a2111o_1
X_15904_ instr_andi _02617_ _02627_ _02643_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__a22o_1
XANTENNA__15914__A _03277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16884_ _03186_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16803__A0 _06586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14409__A2 _07947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18623_ clknet_leaf_10_clk _01683_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15835_ decoded_imm_j\[19\] _05983_ _02596_ _02599_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_144_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12749__S _06869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10694__A3 _05334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_91_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18554_ clknet_leaf_171_clk _01619_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15766_ _02561_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14290__B1 _07944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08528__A irq_mask\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12978_ _07006_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__clkbuf_1
X_17505_ clknet_leaf_15_clk _00674_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_14717_ count_cycle\[9\] _08349_ _07877_ VGND VGND VPWR VPWR _08354_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11929_ _06414_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__clkbuf_1
X_18485_ clknet_leaf_14_clk _01550_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15697_ timer\[10\] _02508_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16745__A _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10851__A0 _04566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15465__S0 _02085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17436_ clknet_leaf_106_clk _00605_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09049__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14648_ _08295_ _08296_ _08297_ VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__o21a_1
XFILLER_0_172_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_17 _03428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _04570_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_39 _05885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17367_ clknet_leaf_111_clk _00536_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14265__A _07905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14579_ _07898_ _07956_ _08050_ _07904_ reg_next_pc\[22\] VGND VGND VPWR VPWR _08235_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_160_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16318_ _06993_ cpuregs.regs\[15\]\[24\] _02881_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17298_ clknet_leaf_109_clk _00472_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16249_ mem_rdata_q\[1\] _03213_ _03914_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput102 net102 VGND VGND VPWR VPWR cpi_rs2[12] sky130_fd_sc_hd__clkbuf_1
XANTENNA__09447__S1 _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput113 net113 VGND VGND VPWR VPWR cpi_rs2[22] sky130_fd_sc_hd__buf_1
Xoutput124 net124 VGND VGND VPWR VPWR cpi_rs2[3] sky130_fd_sc_hd__buf_1
XFILLER_0_3_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput135 net135 VGND VGND VPWR VPWR eoi[13] sky130_fd_sc_hd__buf_1
XFILLER_0_11_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput146 net146 VGND VGND VPWR VPWR eoi[23] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput157 net157 VGND VGND VPWR VPWR eoi[4] sky130_fd_sc_hd__buf_1
XANTENNA__11828__S _06359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15096__A _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13609__A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput168 net168 VGND VGND VPWR VPWR mem_addr[15] sky130_fd_sc_hd__clkbuf_1
XANTENNA__12108__A0 _06193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput179 net179 VGND VGND VPWR VPWR mem_addr[26] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_54_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08710__B net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08958__S0 _03661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09623_ _04352_ _04350_ _04349_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12659__S _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13344__A _07210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09554_ _04284_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_167_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14281__B1 _07942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08438__A net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09033__S _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08505_ instr_sw instr_sh instr_sb _03287_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__or4b_1
XFILLER_0_66_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10179__S _04065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09485_ _04216_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__buf_6
XFILLER_0_77_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15456__S0 _02074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09968__S _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08436_ _03198_ _03221_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11398__A1 _03867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11398__B2 _03880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10260_ cpuregs.regs\[24\]\[24\] cpuregs.regs\[25\]\[24\] cpuregs.regs\[26\]\[24\]
+ cpuregs.regs\[27\]\[24\] _04329_ _04218_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__mux4_1
XANTENNA__09212__A0 mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_148_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10191_ _04903_ _04904_ _04064_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15836__A1 _08232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08949__S0 _03661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13950_ _07732_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12901_ _06954_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_161_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13881_ _07684_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15620_ _02443_ _02445_ _02448_ _03675_ _03654_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__a221o_2
X_12832_ _06157_ cpuregs.regs\[6\]\[8\] _06906_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14272__B1 _07942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15551_ cpuregs.regs\[20\]\[27\] cpuregs.regs\[21\]\[27\] cpuregs.regs\[22\]\[27\]
+ cpuregs.regs\[23\]\[27\] _01979_ _01980_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__mux4_1
X_12763_ cpuregs.regs\[9\]\[8\] _06550_ _06869_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16013__A1 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15447__S0 _02030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14502_ decoded_imm_j\[16\] _07941_ VGND VGND VPWR VPWR _08164_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11714_ _06266_ cpuregs.regs\[10\]\[21\] _06258_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__mux2_1
X_18270_ clknet_leaf_26_clk _01341_ VGND VGND VPWR VPWR decoded_imm\[28\] sky130_fd_sc_hd__dfxtp_4
X_15482_ cpuregs.regs\[20\]\[23\] cpuregs.regs\[21\]\[23\] cpuregs.regs\[22\]\[23\]
+ cpuregs.regs\[23\]\[23\] _02046_ _02047_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__mux4_1
XFILLER_0_166_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15900__C _02612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12694_ _06839_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17221_ clknet_leaf_148_clk _00395_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14433_ reg_next_pc\[10\] _07947_ _08100_ _08033_ VGND VGND VPWR VPWR _08101_ sky130_fd_sc_hd__a22o_1
XANTENNA__10817__S _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11645_ reg_out\[14\] alu_out_q\[14\] _06068_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17152_ clknet_leaf_174_clk _00326_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09179__A _03916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput15 irq[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14364_ _07915_ _08016_ _07917_ VGND VGND VPWR VPWR _08037_ sky130_fd_sc_hd__a21oi_1
X_11576_ reg_out\[7\] alu_out_q\[7\] _06067_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__mux2_1
Xinput26 irq[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_2
XFILLER_0_80_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput37 mem_rdata[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput48 mem_rdata[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
XFILLER_0_141_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10061__A1 _04271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16103_ _02602_ _02755_ _06023_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__a21oi_1
Xinput59 mem_rdata[4] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_1
XFILLER_0_40_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13315_ _07185_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__clkbuf_1
X_10527_ net110 VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15909__A is_alu_reg_imm VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17083_ clknet_leaf_3_clk _00257_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15524__B1 _02017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10600__A3 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16504__S _02979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14295_ _06863_ _03368_ VGND VGND VPWR VPWR _07972_ sky130_fd_sc_hd__and2_2
XFILLER_0_150_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16034_ _02715_ decoded_imm_j\[6\] _02726_ mem_rdata_q\[26\] _02634_ VGND VGND VPWR
+ VPWR _02729_ sky130_fd_sc_hd__a221o_1
X_10458_ cpuregs.regs\[12\]\[30\] cpuregs.regs\[13\]\[30\] cpuregs.regs\[14\]\[30\]
+ cpuregs.regs\[15\]\[30\] _04487_ _04059_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__mux4_1
X_13246_ _07001_ cpuregs.regs\[8\]\[28\] _07140_ VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11010__B1 _05215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08411__D1 _03196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11875__C _06081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10389_ _04214_ _05096_ _04081_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__a21oi_1
X_13177_ _07112_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10364__A2 _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15827__A1 decoded_imm_j\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12128_ _06520_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__clkbuf_1
X_17985_ clknet_leaf_103_clk _01122_ VGND VGND VPWR VPWR irq_mask\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_165_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09506__A1 _04231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12059_ _06266_ cpuregs.regs\[22\]\[21\] _06482_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__mux2_1
X_16936_ clknet_leaf_120_clk _00117_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08957__S _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09601__S1 _04218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16867_ _06582_ cpuregs.regs\[14\]\[23\] _03174_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18606_ clknet_leaf_163_clk _01671_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_15818_ decoded_imm_j\[9\] _05974_ _02592_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__a21o_1
X_16798_ _03141_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09809__A2 _04049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18537_ clknet_leaf_105_clk _01602_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15749_ timer\[24\] _02547_ _02488_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16004__A1 _03635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15438__S0 _02030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09270_ _04006_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18468_ clknet_leaf_143_clk _01533_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17419_ clknet_leaf_127_clk _00588_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18399_ clknet_leaf_132_clk _01464_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08705__B net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11412__A _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_3_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15515__B1 _02349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09993__A1 _03638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09993__B2 irq_pending\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15610__S0 _01968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08721__A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08985_ mem_16bit_buffer\[13\] _03746_ _03727_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__mux2_4
XANTENNA__11304__A1 _04959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_1014 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09552__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10698__A _05397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09606_ _04051_ _04335_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14254__B1 latched_store VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09537_ _04009_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10815__B1 _05367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09468_ net58 net258 _04035_ net43 _04200_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13521__B decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08419_ mem_la_secondword _03198_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09399_ _04132_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__buf_8
XFILLER_0_81_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13013__S _07021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11430_ _06029_ irq_pending\[4\] _06032_ net27 VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__a31o_1
XANTENNA__09433__B1 _04145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_128_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11240__A0 _04566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11361_ _05969_ _03874_ _05967_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09984__B2 _04024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16324__S _02881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11791__A1 _06116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15601__S0 _03641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13100_ _06991_ cpuregs.regs\[7\]\[23\] _07068_ VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__mux2_1
X_10312_ cpuregs.regs\[24\]\[26\] cpuregs.regs\[25\]\[26\] cpuregs.regs\[26\]\[26\]
+ cpuregs.regs\[27\]\[26\] _04084_ _04086_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14080_ count_instr\[29\] _07818_ count_instr\[30\] VGND VGND VPWR VPWR _07822_ sky130_fd_sc_hd__a21o_1
X_11292_ _04913_ _05916_ _03219_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10243_ reg_pc\[24\] decoded_imm\[24\] VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__nand2_1
X_13031_ _07035_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_163_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10174_ _04875_ _04878_ _04886_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__a21o_1
XANTENNA__15285__A2 _02009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17770_ clknet_leaf_95_clk _00939_ VGND VGND VPWR VPWR count_instr\[41\] sky130_fd_sc_hd__dfxtp_1
X_14982_ irq_mask\[3\] _01864_ _01870_ _08335_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_137_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15690__C1 _06026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16721_ _06987_ cpuregs.regs\[19\]\[21\] _03098_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__mux2_1
X_13933_ _07720_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10649__A3 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12299__S _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16652_ _03063_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13048__A1 _06598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13864_ _07671_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15442__C1 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15603_ _02431_ _02432_ _02110_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12815_ _06905_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__buf_6
XANTENNA_output201_A net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16583_ _06984_ cpuregs.regs\[18\]\[20\] _03026_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__mux2_1
X_13795_ _07632_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15993__B1 _03880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18322_ clknet_leaf_38_clk _01390_ VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13712__A net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15534_ cpuregs.regs\[20\]\[26\] cpuregs.regs\[21\]\[26\] cpuregs.regs\[22\]\[26\]
+ cpuregs.regs\[23\]\[26\] _01995_ _01937_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__mux4_1
X_12746_ _06868_ VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__buf_6
XFILLER_0_57_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18253_ clknet_leaf_24_clk _01324_ VGND VGND VPWR VPWR decoded_imm\[11\] sky130_fd_sc_hd__dfxtp_4
X_15465_ cpuregs.regs\[0\]\[22\] cpuregs.regs\[1\]\[22\] cpuregs.regs\[2\]\[22\] cpuregs.regs\[3\]\[22\]
+ _02085_ _02086_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__mux4_1
XFILLER_0_154_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12677_ _06830_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_146_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17204_ clknet_leaf_113_clk _00378_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13756__C1 _07283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14416_ decoded_imm_j\[8\] _07924_ VGND VGND VPWR VPWR _08085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18184_ clknet_leaf_43_clk _01255_ VGND VGND VPWR VPWR instr_bne sky130_fd_sc_hd__dfxtp_1
X_11628_ reg_out\[12\] alu_out_q\[12\] _06067_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15396_ cpuregs.regs\[4\]\[18\] cpuregs.regs\[5\]\[18\] cpuregs.regs\[6\]\[18\] cpuregs.regs\[7\]\[18\]
+ _02046_ _02047_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17135_ clknet_leaf_124_clk _00309_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14347_ _07988_ _08016_ _08021_ _08012_ VGND VGND VPWR VPWR _08022_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11559_ reg_out\[5\] alu_out_q\[5\] _06067_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__mux2_1
XANTENNA__11782__A1 _06116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17066_ clknet_leaf_139_clk _00240_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_90_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14278_ _03293_ _07944_ _07961_ VGND VGND VPWR VPWR _07962_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16017_ _02715_ decoded_imm_j\[1\] mem_rdata_q\[8\] _02716_ _02633_ VGND VGND VPWR
+ VPWR _02717_ sky130_fd_sc_hd__a221o_1
XANTENNA__13523__A2 decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13229_ _07117_ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__buf_6
XFILLER_0_110_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09822__S1 _04087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08770_ net67 net99 VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__and2b_1
X_17968_ clknet_leaf_4_clk _01105_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16919_ clknet_leaf_18_clk _00100_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15028__A2 _01865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17899_ clknet_leaf_95_clk _01068_ VGND VGND VPWR VPWR count_cycle\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15821__B _03737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12937__S _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16409__S _02932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09322_ _04056_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__buf_8
XFILLER_0_47_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09253_ _03826_ _03894_ _03988_ _03786_ _03992_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10457__S _04121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12238__A _06319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09184_ _03840_ _03922_ _03933_ _03888_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13762__A2 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12672__S _06825_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10576__A2 _05261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11773__A1 _06116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09547__A _04277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10981__C1 _05323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09718__A1 _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10959__S0 _05237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10205__B decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08968_ _03729_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_166_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08899_ _03652_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__buf_6
XANTENNA__10187__S1 _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10930_ _04744_ _04708_ _04642_ _04611_ _05237_ _05240_ VGND VGND VPWR VPWR _05617_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_168_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10861_ _05549_ _05551_ _05363_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__mux2_1
XANTENNA__12847__S _06917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12600_ _06789_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13580_ net73 decoded_imm\[15\] VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10792_ _03530_ _05320_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12531_ cpuregs.regs\[2\]\[0\] _06531_ _06752_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15250_ cpuregs.regs\[12\]\[10\] cpuregs.regs\[13\]\[10\] cpuregs.regs\[14\]\[10\]
+ cpuregs.regs\[15\]\[10\] _01970_ _01971_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__mux4_1
XFILLER_0_163_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12462_ _06078_ cpuregs.regs\[28\]\[0\] _06715_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_173_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10016__A1 _04053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14201_ _07901_ _07907_ VGND VGND VPWR VPWR _07908_ sky130_fd_sc_hd__nand2_1
X_11413_ _03845_ _03971_ _05991_ _06019_ _05960_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__o41a_1
XFILLER_0_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15181_ cpuregs.regs\[16\]\[6\] cpuregs.regs\[17\]\[6\] cpuregs.regs\[18\]\[6\] cpuregs.regs\[19\]\[6\]
+ _01985_ _01986_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12393_ cpuregs.regs\[27\]\[0\] _06531_ _06678_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11764__A1 _06116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10111__S1 _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14132_ count_instr\[43\] _07843_ _07848_ _07858_ VGND VGND VPWR VPWR _07859_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11344_ _05959_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_134_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15050__S1 _01909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14063_ _07810_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__clkbuf_1
X_11275_ _05896_ _05899_ _05902_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11516__B2 _06072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13014_ _07026_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__clkbuf_1
X_10226_ _04054_ _04934_ _04938_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__a21boi_1
XANTENNA__15906__B mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output249_A net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14810__B _01753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15194__A _03646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11926__S _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13707__A _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10157_ irq_mask\[21\] _04448_ timer\[21\] _04024_ _04027_ VGND VGND VPWR VPWR _04872_
+ sky130_fd_sc_hd__a221o_1
X_17822_ clknet_leaf_67_clk _00991_ VGND VGND VPWR VPWR reg_pc\[30\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_100_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15663__C1 _07775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09568__S0 _04275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17753_ clknet_leaf_85_clk _00922_ VGND VGND VPWR VPWR count_instr\[24\] sky130_fd_sc_hd__dfxtp_1
X_14965_ _01858_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__clkbuf_1
X_10088_ _04792_ _04796_ _04100_ _04804_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__a211o_4
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10178__S1 _04470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13916_ _07691_ _07708_ VGND VGND VPWR VPWR _07709_ sky130_fd_sc_hd__and2_1
X_16704_ _06970_ cpuregs.regs\[19\]\[13\] _03087_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17684_ clknet_leaf_100_clk _00853_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14896_ _05205_ _01812_ _01816_ _01820_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__o22a_1
X_16635_ _03054_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13847_ cpuregs.regs\[0\]\[20\] VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12757__S _06869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14538__A decoded_imm_j\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13442__A _07209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16566_ _06968_ cpuregs.regs\[18\]\[12\] _03015_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__mux2_1
XANTENNA__08448__A1 _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13778_ _07304_ _05107_ _07211_ reg_pc\[28\] _07221_ VGND VGND VPWR VPWR _07617_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__13441__A1 _03275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15517_ cpuregs.regs\[0\]\[25\] cpuregs.regs\[1\]\[25\] cpuregs.regs\[2\]\[25\] cpuregs.regs\[3\]\[25\]
+ _02030_ _02031_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__mux4_1
X_18305_ clknet_leaf_35_clk _01373_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dfxtp_1
XANTENNA__15718__B1 _02488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11452__B1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12729_ _06857_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__clkbuf_1
X_16497_ _02981_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_44_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18236_ clknet_leaf_8_clk _01307_ VGND VGND VPWR VPWR cpuregs.raddr1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15448_ cpuregs.regs\[12\]\[21\] cpuregs.regs\[13\]\[21\] cpuregs.regs\[14\]\[21\]
+ cpuregs.regs\[15\]\[21\] _01976_ _01977_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1013 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09948__A1 _03297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18167_ clknet_leaf_32_clk _01238_ VGND VGND VPWR VPWR decoded_imm_j\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15379_ _03659_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17118_ clknet_leaf_167_clk _00292_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09367__A _04051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18098_ clknet_leaf_92_clk _01202_ VGND VGND VPWR VPWR timer\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08620__A1 _03304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09940_ irq_mask\[15\] _04021_ timer\[15\] _04023_ _04188_ VGND VGND VPWR VPWR _04661_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17049_ clknet_leaf_13_clk _00223_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10306__A reg_pc\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09871_ irq_mask\[13\] _04448_ timer\[13\] _04024_ _04027_ VGND VGND VPWR VPWR _04594_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__11836__S _06359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08822_ net117 net85 VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__and2b_1
XANTENNA__09814__B decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08753_ net127 net95 VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10041__A _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08684_ net117 net85 VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__nor2_1
XANTENNA__10494__A1 _04289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11691__B1 _06066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14448__A decoded_imm_j\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09305_ net63 net49 _04040_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09976__S _04369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09236_ _03754_ _03759_ _03760_ _03753_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__a22o_2
XFILLER_0_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15280__S1 _02000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09167_ mem_rdata_q\[18\] _03918_ _03914_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11746__A1 _06252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09277__A _04013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09098_ _03834_ _03856_ _03857_ _03789_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13499__A1 _04419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11060_ _05720_ _05737_ _03454_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_112_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10011_ cpuregs.regs\[0\]\[17\] cpuregs.regs\[1\]\[17\] cpuregs.regs\[2\]\[17\] cpuregs.regs\[3\]\[17\]
+ _04477_ _04478_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__mux4_1
XANTENNA__10650__S _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10721__A2 _05301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12150__B _06081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13120__A0 _06941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14750_ count_cycle\[19\] count_cycle\[20\] _01715_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__and3_1
X_11962_ _06432_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13701_ _04913_ decoded_imm\[22\] _07527_ VGND VGND VPWR VPWR _07545_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09740__A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10913_ _05600_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11682__B1 _06066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09970__S0 _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12577__S _06774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14681_ _07971_ _08322_ _07986_ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_158_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _06395_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16420_ _02940_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__clkbuf_1
X_13632_ _07284_ _07471_ _07480_ VGND VGND VPWR VPWR _07481_ sky130_fd_sc_hd__o21a_1
X_10844_ _03499_ _05535_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_4_11_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16351_ _06957_ cpuregs.regs\[16\]\[7\] _02896_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__mux2_1
XANTENNA__11434__B1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13563_ _04602_ _07416_ _07374_ VGND VGND VPWR VPWR _07417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10775_ _05233_ _05234_ _05267_ _05270_ _05413_ _05414_ VGND VGND VPWR VPWR _05471_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15302_ net102 _02081_ _02148_ _02149_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__o22a_1
XANTENNA__10788__A2 _03518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12514_ _06297_ cpuregs.regs\[28\]\[25\] _06737_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16282_ _06957_ cpuregs.regs\[15\]\[7\] _02859_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__mux2_1
X_13494_ _07350_ _07351_ VGND VGND VPWR VPWR _07352_ sky130_fd_sc_hd__nor2_1
XANTENNA__11213__C _05851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output199_A net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18021_ clknet_leaf_104_clk _00028_ VGND VGND VPWR VPWR irq_pending\[5\] sky130_fd_sc_hd__dfxtp_1
X_15233_ cpuregs.regs\[4\]\[9\] cpuregs.regs\[5\]\[9\] cpuregs.regs\[6\]\[9\] cpuregs.regs\[7\]\[9\]
+ _01976_ _01977_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__mux4_1
XANTENNA__15271__S1 _01971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12445_ cpuregs.regs\[27\]\[25\] _06586_ _06700_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11737__A1 _06252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15164_ _02017_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__clkbuf_8
X_12376_ cpuregs.regs\[26\]\[25\] _06586_ _06663_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14115_ _07845_ _07846_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__nor2_1
X_11327_ _05945_ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16512__S _02979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15095_ _01941_ _01945_ _01949_ _01953_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__o22a_2
XANTENNA_output76_A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14046_ count_instr\[19\] count_instr\[15\] _07787_ _07795_ VGND VGND VPWR VPWR _07799_
+ sky130_fd_sc_hd__and4_1
XANTENNA__09789__S0 _04512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11258_ reg_next_pc\[16\] reg_out\[16\] _05876_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__mux2_1
XANTENNA__15636__B _03254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12162__A1 _06540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10209_ count_instr\[55\] _04015_ _04011_ count_instr\[23\] VGND VGND VPWR VPWR _04922_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11189_ _05831_ _05832_ _05829_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17805_ clknet_leaf_62_clk _00974_ VGND VGND VPWR VPWR reg_pc\[13\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__13337__S1 _04284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15997_ _03893_ _05990_ _05976_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14948_ _01849_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17736_ clknet_leaf_96_clk _00905_ VGND VGND VPWR VPWR count_instr\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11673__B1 _06066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14879_ count_cycle\[61\] _01804_ _01806_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12487__S _06726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17667_ clknet_leaf_8_clk _00836_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16618_ _03045_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_63_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17598_ clknet_leaf_129_clk _00767_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15798__S _08033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09713__S0 _04217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16549_ _06951_ cpuregs.regs\[18\]\[4\] _03004_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10323__S1 _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09021_ _03206_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__clkbuf_4
X_18219_ clknet_leaf_92_clk _01290_ VGND VGND VPWR VPWR instr_rdinstr sky130_fd_sc_hd__dfxtp_4
XFILLER_0_26_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15262__S1 _02014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11728__A1 _06252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16667__A1 _06319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10400__B2 instr_timer VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12950__S _06985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10036__A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10951__A2 _05215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09923_ cpuregs.regs\[16\]\[15\] cpuregs.regs\[17\]\[15\] cpuregs.regs\[18\]\[15\]
+ cpuregs.regs\[19\]\[15\] _04472_ _04473_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__mux4_1
XANTENNA__09149__A2 _03880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09854_ _04483_ _04576_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__nand2_1
X_08805_ _03478_ _03570_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__nand2_1
X_09785_ _04508_ _04509_ _04287_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__mux2_1
X_08736_ _03501_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__inv_2
XANTENNA_107 _06482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10467__A1 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09560__A _04290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10011__S0 _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11664__B1 _06066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_118 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08667_ net91 net123 VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__nand2_1
XANTENNA_129 net223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12397__S _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13405__A1 _03276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09609__B1 _04009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08598_ irq_state\[1\] irq_state\[0\] VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08607__C _00865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09704__S0 _04325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10560_ _05263_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__buf_4
XFILLER_0_146_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08904__A _00064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_130_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14625__B _07964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09219_ _03864_ _03958_ _03961_ _03927_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_20_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10491_ cpuregs.regs\[8\]\[31\] cpuregs.regs\[9\]\[31\] cpuregs.regs\[10\]\[31\]
+ cpuregs.regs\[11\]\[31\] _04329_ _04218_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_101_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13021__S _07021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12230_ cpuregs.regs\[24\]\[25\] _06586_ _06576_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12161_ _06113_ VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__buf_2
XANTENNA__12860__S _06928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_145_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10942__A2 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11112_ _03444_ _05785_ _05517_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__a21o_1
XANTENNA__15330__A1 _02012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12092_ _06501_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13341__B1 _04227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11043_ instr_sub _03457_ _05720_ _05721_ _03585_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__o32a_1
X_15920_ mem_rdata_q\[30\] _02654_ _02655_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__and3_1
XANTENNA__12161__A _06113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13892__A1 _03327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15851_ _02610_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_110_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13691__S _07224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15094__B1 _03674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_14802_ _01755_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__clkbuf_1
X_15782_ _02572_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__clkbuf_1
X_18570_ clknet_leaf_122_clk _01635_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09848__B1 _04012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12994_ cpuregs.regs\[3\]\[5\] _06544_ _07010_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14733_ _08364_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__clkbuf_1
X_17521_ clknet_leaf_136_clk _00690_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10002__S0 _04472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11655__B1 _06066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11945_ _06385_ _06422_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__nand2_4
XFILLER_0_99_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output114_A net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17452_ clknet_leaf_159_clk _00621_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _07968_ _08301_ VGND VGND VPWR VPWR _08313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11876_ _06383_ _06385_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__nand2_4
X_16403_ _06422_ _06713_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__nand2_4
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13615_ _03575_ _07236_ VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10827_ _05517_ _05518_ _05519_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__a21o_1
XANTENNA__11224__B _05860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17383_ clknet_leaf_180_clk _00552_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14595_ _03379_ _08248_ _08249_ VGND VGND VPWR VPWR _08250_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16334_ cpuregs.waddr\[2\] _06082_ _06083_ _06081_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__and4bb_4
X_13546_ _07394_ _07397_ _07400_ VGND VGND VPWR VPWR _07401_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10758_ _05380_ _05382_ _05395_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15244__S1 _02075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16265_ _02857_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__clkbuf_1
X_13477_ _03275_ _07329_ _07330_ _07334_ _07336_ VGND VGND VPWR VPWR _07337_ sky130_fd_sc_hd__a32o_1
XFILLER_0_152_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10689_ _03606_ _05388_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18004_ clknet_leaf_66_clk _01141_ VGND VGND VPWR VPWR irq_mask\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15216_ _02066_ _02067_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__or2_1
X_12428_ cpuregs.regs\[27\]\[17\] _06569_ _06689_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__mux2_1
X_16196_ _02814_ _02817_ _02818_ _02676_ net297 VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14372__A2 _07994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15147_ _03653_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__buf_8
XFILLER_0_168_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12359_ cpuregs.regs\[26\]\[17\] _06569_ _06652_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__mux2_1
XANTENNA__12770__S _06880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14551__A _07952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15321__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15078_ _03646_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_56_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13332__B1 _04225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14029_ count_instr\[14\] count_instr\[13\] count_instr\[12\] _07781_ VGND VGND VPWR
+ VPWR _07787_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_56_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09570_ _04299_ _04300_ _04287_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__mux2_1
XANTENNA__13635__A1 _04754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15180__S0 _02022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15813__C _03878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08521_ cpu_state\[2\] VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__buf_4
XFILLER_0_26_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17719_ clknet_leaf_83_clk _00888_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dfxtp_1
XANTENNA__11646__B1 _06066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09934__S0 _04487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16034__C1 _02634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13106__S _07068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08452_ _03196_ _03232_ _03235_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__or3b_1
XANTENNA__16585__A0 _06987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15483__S1 _02047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16417__S _02932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12071__A0 _06312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16337__A0 _06941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08724__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09004_ mem_16bit_buffer\[15\] _03727_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11177__A2 _04710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12374__A1 _06584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15557__A _01984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12680__S _06825_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10480__S0 _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14180__B _07815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09906_ _04626_ _04627_ _04369_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09837_ _04548_ _04552_ _04560_ net300 VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__a211o_4
XANTENNA__17922__D _08391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09768_ _04051_ _04493_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__nor2_1
XANTENNA__09290__A _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08719_ _03483_ _03484_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__and2_1
X_09699_ irq_pending\[8\] _04007_ _04418_ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_107_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11101__A2 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11730_ _06280_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_25_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ reg_pc\[16\] _06210_ _06101_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09058__A1 mem_rdata_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12855__S _06917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11391__C_N _03965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13400_ _07209_ _04186_ _07210_ reg_pc\[3\] VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__a22o_1
X_10612_ net88 net90 _05263_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14380_ decoded_imm_j\[6\] _07919_ VGND VGND VPWR VPWR _08052_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11592_ _06157_ cpuregs.regs\[10\]\[8\] _06086_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10612__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13331_ _07196_ _07197_ _04211_ VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__mux2_1
X_10543_ _04033_ _05230_ _05235_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16050_ _03402_ decoded_imm_j\[13\] _03403_ _02613_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13262_ _06949_ cpuregs.regs\[5\]\[3\] _07154_ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10474_ reg_pc\[31\] decoded_imm\[31\] VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11168__A2 _05277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15001_ _01881_ _01869_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12213_ _06256_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13193_ _07121_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09465__A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12144_ _06528_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16952_ clknet_leaf_53_clk _00080_ VGND VGND VPWR VPWR cpu_state\[6\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_21_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12075_ _06328_ cpuregs.regs\[22\]\[29\] _06482_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__mux2_1
X_11026_ _03458_ _05222_ _05597_ _05254_ _05705_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__a221o_1
X_15903_ instr_ori _02618_ _02626_ _02643_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__a22o_1
XANTENNA__10223__S0 _04280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15914__B is_alu_reg_reg VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output231_A net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16883_ _06598_ cpuregs.regs\[14\]\[31\] _03151_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15067__B1 _03675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11934__S _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18622_ clknet_leaf_10_clk _01682_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15834_ _05969_ _03634_ _03920_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__and3_1
XANTENNA__13617__A1 _04708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ clknet_leaf_1_clk _01618_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_15765_ timer\[28\] _03425_ _02560_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__or3_1
X_12977_ _07005_ cpuregs.regs\[31\]\[30\] _06942_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08528__B irq_active VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15930__A is_alu_reg_imm VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17504_ clknet_leaf_170_clk _00673_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14716_ count_cycle\[7\] count_cycle\[8\] count_cycle\[9\] _08346_ VGND VGND VPWR
+ VPWR _08353_ sky130_fd_sc_hd__and4_2
X_11928_ _06289_ cpuregs.regs\[20\]\[24\] _06409_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15696_ timer\[10\] _02508_ _02476_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__a21o_1
X_18484_ clknet_leaf_170_clk _01549_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16745__B _01955_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10851__A1 _04532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15465__S1 _02086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17435_ clknet_leaf_166_clk _00604_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_14647_ _08295_ _08296_ _08055_ VGND VGND VPWR VPWR _08297_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12765__S _06869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11859_ _06297_ cpuregs.regs\[11\]\[25\] _06370_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__mux2_1
XANTENNA__08792__A_N net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13450__A net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 _03600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15790__A1 _04156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17366_ clknet_leaf_114_clk _00535_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_14578_ _08231_ _08233_ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13529_ _07304_ _04526_ _07211_ reg_pc\[11\] _07221_ VGND VGND VPWR VPWR _07385_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16317_ _02885_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17297_ clknet_leaf_114_clk _00471_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16248_ _02848_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput103 net103 VGND VGND VPWR VPWR cpi_rs2[13] sky130_fd_sc_hd__buf_1
XFILLER_0_140_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput114 net114 VGND VGND VPWR VPWR cpi_rs2[23] sky130_fd_sc_hd__clkbuf_1
X_16179_ net283 net245 _02770_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput125 net125 VGND VGND VPWR VPWR cpi_rs2[4] sky130_fd_sc_hd__clkbuf_1
XANTENNA__09221__B2 _03737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput136 net136 VGND VGND VPWR VPWR eoi[14] sky130_fd_sc_hd__buf_1
Xoutput147 net147 VGND VGND VPWR VPWR eoi[24] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput158 net158 VGND VGND VPWR VPWR eoi[5] sky130_fd_sc_hd__clkbuf_1
XANTENNA__09772__A2 _04013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15096__B _01954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13609__B decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput169 net169 VGND VGND VPWR VPWR mem_addr[16] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12005__S _06446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16700__S _03087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10314__A _04052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09524__A2 _04250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11867__A0 _06328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08958__S1 _03662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11844__S _06359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09622_ reg_pc\[5\] decoded_imm\[5\] VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09553_ _04283_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__buf_6
XANTENNA__14281__A1 reg_next_pc\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08504_ _03196_ _03278_ cpu_state\[5\] _03286_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__and4bb_1
XANTENNA__15840__A _03215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09484_ _04055_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__buf_6
XFILLER_0_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08435_ _03218_ _03219_ _03220_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__o21ai_2
XANTENNA__15456__S1 _02075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08454__A mem_do_prefetch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12595__A1 _06598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13792__B1 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09269__B cpu_state\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10070__A2 _04104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09212__A1 _03954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10358__B1 _04237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14191__A _07898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09285__A _04021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16089__A2 _02711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10190_ cpuregs.regs\[8\]\[22\] cpuregs.regs\[9\]\[22\] cpuregs.regs\[10\]\[22\]
+ cpuregs.regs\[11\]\[22\] _04084_ _04086_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_148_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08971__A0 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15392__S0 _01995_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08949__S1 _03662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12900_ _06953_ cpuregs.regs\[31\]\[5\] _06943_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__mux2_1
X_13880_ _07675_ _07683_ VGND VGND VPWR VPWR _07684_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_161_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10530__A0 _04566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16797__A0 _06580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09224__S _03757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12831_ _06914_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__clkbuf_1
X_15550_ _02383_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12762_ _06877_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16013__A2 _02711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14501_ _08120_ _08162_ VGND VGND VPWR VPWR _08163_ sky130_fd_sc_hd__nor2_1
XANTENNA__15447__S1 _02031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11713_ _06265_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__buf_2
XFILLER_0_68_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15481_ _03719_ _02317_ _03674_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12693_ _06193_ cpuregs.regs\[12\]\[12\] _06836_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__mux2_1
XANTENNA__12585__S _06774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17220_ clknet_leaf_159_clk _00394_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_14432_ _08099_ VGND VGND VPWR VPWR _08100_ sky130_fd_sc_hd__inv_2
X_11644_ reg_pc\[14\] _06195_ _06203_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__o21a_1
XFILLER_0_166_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15772__A1 _05139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17151_ clknet_leaf_179_clk _00325_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14363_ _07915_ _07917_ _08016_ VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__and3_1
Xinput16 irq[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
X_11575_ _06142_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09451__A1 _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput27 irq[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
XANTENNA__08885__S0 _03649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16102_ _03783_ _03856_ _05961_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__o21ba_1
Xinput38 mem_rdata[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09894__S _04222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13314_ _07001_ cpuregs.regs\[5\]\[28\] _07176_ VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__mux2_1
Xinput49 mem_rdata[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
X_10526_ _05229_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__buf_4
XANTENNA__10061__A2 _04777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17082_ clknet_leaf_189_clk _00256_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15524__A1 _02012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16721__A0 _06987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14294_ reg_pc\[31\] _07953_ _07971_ _07960_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15909__B _02611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output181_A net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16033_ mem_rdata_q\[25\] _02711_ _02726_ _02728_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__a31o_1
X_13245_ _07148_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__clkbuf_1
X_10457_ _05161_ _05162_ _04121_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09195__A _03916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08411__C1 latched_branch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13176_ _06999_ cpuregs.regs\[4\]\[27\] _07104_ VGND VGND VPWR VPWR _07112_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10388_ _05094_ _05095_ _04320_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__mux2_1
X_12127_ _06266_ cpuregs.regs\[23\]\[21\] _06518_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__mux2_1
X_17984_ clknet_leaf_103_clk _01121_ VGND VGND VPWR VPWR irq_mask\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15383__S0 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11849__A0 _06257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12058_ _06483_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__clkbuf_1
X_16935_ clknet_leaf_101_clk _00116_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11009_ _05689_ _05644_ _05277_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__mux2_1
XANTENNA__09911__C1 _04188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16788__A0 _06571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16866_ _03177_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08539__A is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18605_ clknet_leaf_121_clk _01670_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_15817_ _03892_ _06016_ _02587_ _03994_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__a22o_1
XANTENNA__14263__A1 reg_next_pc\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16797_ _06580_ cpuregs.regs\[13\]\[22\] _03138_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__mux2_1
XANTENNA__15460__B1 _02197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18536_ clknet_leaf_152_clk _01601_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15748_ _04941_ _02506_ _02548_ _02545_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10285__C1 _04289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16004__A2 _03763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15438__S1 _02031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12495__S _06726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18467_ clknet_leaf_148_clk _01532_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09690__A1 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15679_ timer\[6\] _02495_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17418_ clknet_leaf_185_clk _00587_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15763__A1 _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14566__A2 _07952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18398_ clknet_leaf_179_clk _01463_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13774__A0 _05143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12577__A1 _06580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11412__B _03892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17349_ clknet_leaf_174_clk _00518_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15515__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09993__A2 _04708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14723__B _08350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15610__S1 _03639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08721__B net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15279__B1 _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10044__A _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16430__S _02943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08984_ _03744_ _03745_ _03230_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__mux2_1
XANTENNA__11574__S _06086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15126__S0 _01979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09605_ _04316_ _04323_ _04100_ _04334_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__a211o_4
XANTENNA__14254__A1 latched_branch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09536_ _03637_ _04262_ _04265_ _03225_ _04266_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__a221o_1
XANTENNA__09979__S _04320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09467_ _04036_ mem_wordsize\[1\] _04199_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08418_ _03201_ _03202_ _03203_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09398_ cpuregs.raddr1\[3\] cpuregs.raddr1\[2\] cpuregs.raddr1\[4\] _04098_ VGND
+ VGND VPWR VPWR _04132_ sky130_fd_sc_hd__or4_1
XFILLER_0_93_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12568__A1 _06571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16605__S _03003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09984__A2 _04022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11360_ _05973_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__buf_2
XFILLER_0_116_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11791__A2 reg_next_pc\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11749__S _06258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10311_ cpuregs.regs\[28\]\[26\] cpuregs.regs\[29\]\[26\] cpuregs.regs\[30\]\[26\]
+ cpuregs.regs\[31\]\[26\] _04084_ _04086_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__mux4_1
XANTENNA__15601__S1 _03684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11291_ _05913_ _05915_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12434__A _06677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13030_ cpuregs.regs\[3\]\[22\] _06580_ _07032_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__mux2_1
X_10242_ _04824_ _04949_ _04951_ _04953_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__o211a_1
XANTENNA__10426__S0 _04273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12740__A1 cpuregs.waddr\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12740__B2 _06861_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10173_ _04875_ _04878_ _04886_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__nand3_1
XANTENNA__15365__S0 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09743__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14981_ _04185_ _01869_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__nor2_1
X_16720_ _03099_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__clkbuf_1
X_13932_ _07714_ _07719_ VGND VGND VPWR VPWR _07720_ sky130_fd_sc_hd__and2_1
XANTENNA__15117__S0 _01970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13863_ cpuregs.regs\[0\]\[28\] VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__clkbuf_1
X_16651_ cpuregs.regs\[1\]\[20\] _06256_ _03062_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__mux2_1
XANTENNA__14245__A1 reg_next_pc\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15602_ cpuregs.regs\[8\]\[30\] cpuregs.regs\[9\]\[30\] cpuregs.regs\[10\]\[30\]
+ cpuregs.regs\[11\]\[30\] _03641_ _03684_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__mux4_1
X_12814_ _06080_ _06904_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__nand2_4
X_13794_ _05143_ _07631_ _07224_ VGND VGND VPWR VPWR _07632_ sky130_fd_sc_hd__mux2_1
X_16582_ _03003_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__buf_6
XFILLER_0_158_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18321_ clknet_leaf_38_clk _01389_ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dfxtp_1
XANTENNA__10267__C1 _04133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13712__B decoded_imm\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12745_ cpuregs.waddr\[2\] _06081_ _06082_ _06601_ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15533_ _03709_ _02366_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13204__S _07118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15464_ cpuregs.regs\[4\]\[22\] cpuregs.regs\[5\]\[22\] cpuregs.regs\[6\]\[22\] cpuregs.regs\[7\]\[22\]
+ _01973_ _01974_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__mux4_1
X_18252_ clknet_leaf_22_clk _01323_ VGND VGND VPWR VPWR decoded_imm\[10\] sky130_fd_sc_hd__dfxtp_4
X_12676_ _06125_ cpuregs.regs\[12\]\[4\] _06825_ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17203_ clknet_leaf_109_clk _00377_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_14415_ _08082_ _08083_ VGND VGND VPWR VPWR _08084_ sky130_fd_sc_hd__nand2_1
X_11627_ _06187_ _06118_ _06188_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__and3b_1
X_18183_ clknet_leaf_41_clk _01254_ VGND VGND VPWR VPWR instr_beq sky130_fd_sc_hd__dfxtp_1
X_15395_ _03709_ _02236_ _00068_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__o21a_1
XANTENNA__16515__S _02990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11231__A1 _05829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17134_ clknet_leaf_123_clk _00308_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_14346_ _08019_ _08020_ VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__xnor2_1
X_11558_ reg_pc\[5\] _06121_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08830__A_N net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10509_ instr_or instr_ori VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__or2_2
X_17065_ clknet_leaf_142_clk _00239_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14277_ _05909_ _06294_ _07945_ reg_next_pc\[25\] VGND VGND VPWR VPWR _07961_ sky130_fd_sc_hd__o22a_1
X_11489_ net65 net262 _03305_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__and3b_1
XANTENNA__12344__A _06640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16016_ is_beq_bne_blt_bge_bltu_bgeu is_sb_sh_sw VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__or2_1
X_13228_ _07139_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13159_ _06982_ cpuregs.regs\[4\]\[19\] _07093_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__mux2_1
XANTENNA__15356__S0 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09653__A _04100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17967_ clknet_leaf_0_clk _01104_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dfxtp_1
XANTENNA__14484__A1 reg_next_pc\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14484__B2 _07960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11298__A1 _03460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16918_ clknet_leaf_187_clk _00099_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_17898_ clknet_leaf_94_clk _01067_ VGND VGND VPWR VPWR count_cycle\[43\] sky130_fd_sc_hd__dfxtp_1
X_16849_ _03168_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13444__C1 _07283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09321_ _04055_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_66_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18519_ clknet_leaf_17_clk _01584_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13995__B1 _07759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11423__A _03412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13114__S _07045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09252_ _03957_ _03989_ _03991_ _03932_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__o31a_1
XANTENNA__15736__A1 _04842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15197__C1 _03639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13747__B1 _07210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09183_ _03790_ _03923_ _03931_ _03932_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12953__S _06985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08732__A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11773__A2 reg_next_pc\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16161__A1 net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12254__A _06603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15595__S0 _01968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09039__S _03730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15347__S0 _01999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08967_ _03200_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11289__A1 _03575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08898_ cpuregs.regs\[16\]\[2\] cpuregs.regs\[17\]\[2\] cpuregs.regs\[18\]\[2\] cpuregs.regs\[19\]\[2\]
+ _03661_ _03662_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10497__C1 _04188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10860_ _03497_ _05550_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14628__B _07964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12789__A1 _06575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09519_ net93 VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__clkbuf_4
X_10791_ _03514_ _05440_ _05399_ _05485_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_39_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12530_ _06751_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__buf_6
XFILLER_0_137_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12461_ _06714_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_173_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14200_ reg_next_pc\[2\] _06099_ _03189_ VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__mux2_1
X_11412_ _03783_ _03892_ _03923_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__and3_1
X_15180_ cpuregs.regs\[20\]\[6\] cpuregs.regs\[21\]\[6\] cpuregs.regs\[22\]\[6\] cpuregs.regs\[23\]\[6\]
+ _02022_ _02023_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__mux4_1
X_12392_ _06677_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14131_ count_instr\[45\] count_instr\[44\] VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__and2_1
XANTENNA__11764__A2 reg_next_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11343_ _05205_ _05958_ _03219_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16152__A1 net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12164__A _06124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15586__S0 _03641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14062_ _07808_ _07778_ _07809_ VGND VGND VPWR VPWR _07810_ sky130_fd_sc_hd__and3b_1
XFILLER_0_120_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11274_ reg_next_pc\[19\] reg_out\[19\] _05898_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__mux2_2
XANTENNA__11516__A2 reg_next_pc\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13013_ cpuregs.regs\[3\]\[14\] _06563_ _07021_ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__mux2_1
X_10225_ _04069_ _04937_ _04081_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15338__S0 _01979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15906__C mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17821_ clknet_leaf_67_clk _00990_ VGND VGND VPWR VPWR reg_pc\[29\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__13707__B decoded_imm\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10156_ _04858_ _04862_ _04870_ _04227_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_146_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17752_ clknet_leaf_85_clk _00921_ VGND VGND VPWR VPWR count_instr\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09568__S1 _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10412__A _03384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14964_ _07737_ _01857_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__and2_1
X_10087_ _04483_ _04799_ _04803_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__a21oi_1
X_16703_ _03090_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__clkbuf_1
X_13915_ _03335_ _07704_ _07705_ net133 VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__a22o_1
X_17683_ clknet_leaf_152_clk _00852_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_14895_ _01812_ _01819_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__nand2_1
XANTENNA__15415__B1 _00067_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16634_ cpuregs.regs\[1\]\[12\] _06192_ _03051_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__mux2_1
X_13846_ _07662_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15510__S0 _01985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08817__A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14538__B _07950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13777_ _07238_ _07613_ _07615_ _07232_ VGND VGND VPWR VPWR _07616_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16565_ _03017_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08448__A2 _03228_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10989_ _05281_ _05668_ _05670_ _05671_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__a211o_1
XANTENNA__15879__B_N decoder_trigger VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18304_ clknet_leaf_6_clk _01372_ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15516_ cpuregs.regs\[4\]\[25\] cpuregs.regs\[5\]\[25\] cpuregs.regs\[6\]\[25\] cpuregs.regs\[7\]\[25\]
+ _01979_ _01980_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__mux4_1
XFILLER_0_167_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12728_ _06328_ cpuregs.regs\[12\]\[29\] _06847_ VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16496_ cpuregs.regs\[17\]\[11\] _06557_ _02979_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18235_ clknet_leaf_9_clk _01306_ VGND VGND VPWR VPWR cpuregs.raddr1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12659_ _06328_ cpuregs.regs\[30\]\[29\] _06810_ VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__mux2_1
X_15447_ cpuregs.regs\[0\]\[21\] cpuregs.regs\[1\]\[21\] cpuregs.regs\[2\]\[21\] cpuregs.regs\[3\]\[21\]
+ _02030_ _02031_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_61_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18166_ clknet_leaf_24_clk _01237_ VGND VGND VPWR VPWR decoded_imm_j\[7\] sky130_fd_sc_hd__dfxtp_1
X_15378_ _03658_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__buf_6
XFILLER_0_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11755__A2 reg_next_pc\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17117_ clknet_leaf_13_clk _00291_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09367__B _04101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14329_ _07908_ _08003_ VGND VGND VPWR VPWR _08005_ sky130_fd_sc_hd__and2_1
X_18097_ clknet_leaf_92_clk _01201_ VGND VGND VPWR VPWR timer\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15577__S0 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17048_ clknet_leaf_176_clk _00222_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15351__C1 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10306__B decoded_imm\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08908__B1 _00067_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09870_ _04592_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__inv_2
XANTENNA__15329__S0 _02069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08821_ net116 _03584_ _03586_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__o21a_1
XANTENNA__09383__A _04040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15103__C1 _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_370 VGND VGND VPWR VPWR alphacore_370/HI trace_data[31] sky130_fd_sc_hd__conb_1
XANTENNA__12468__A0 _06114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11418__A _06003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08752_ net96 VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08683_ _03447_ _03448_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_136_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11140__B1 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15406__B1 _03657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15501__S0 _01990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09304_ _04039_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08446__B _03229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15709__A1 _04593_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09235_ _03786_ _03837_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10992__A _05255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14464__A decoded_imm_j\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09558__A _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09166_ _03850_ _03811_ _03812_ _03849_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10403__C1 _05110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15568__S0 _02030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09097_ _03743_ _03782_ _03853_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_165_Left_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13499__A2 _05260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10010_ cpuregs.regs\[4\]\[17\] cpuregs.regs\[5\]\[17\] cpuregs.regs\[6\]\[17\] cpuregs.regs\[7\]\[17\]
+ _04477_ _04478_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__mux4_1
X_09999_ _04716_ _04717_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__nand2_1
XANTENNA__13019__S _07021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10232__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12150__C _06082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11961_ _06150_ cpuregs.regs\[21\]\[7\] _06424_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__mux2_1
XANTENNA__12858__S _06928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11762__S _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13700_ _07542_ _07543_ VGND VGND VPWR VPWR _07544_ sky130_fd_sc_hd__nand2_1
XANTENNA__13543__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10912_ _05244_ _05250_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__nor2_2
XFILLER_0_86_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14680_ _07971_ _08322_ VGND VGND VPWR VPWR _08327_ sky130_fd_sc_hd__nand2_1
X_11892_ _06150_ cpuregs.regs\[20\]\[7\] _06387_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__mux2_1
XANTENNA__09970__S1 _04478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13631_ _03275_ _07476_ _07479_ _07232_ VGND VGND VPWR VPWR _07480_ sky130_fd_sc_hd__a211o_1
X_10843_ _03556_ _05534_ _05390_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13562_ _07284_ _07405_ _07415_ VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__o21a_1
X_16350_ _02903_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__clkbuf_1
X_10774_ _03512_ _05469_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__xor2_1
XFILLER_0_149_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15301_ decoded_imm\[12\] _02009_ _01963_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__a21o_1
XANTENNA__10788__A3 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12513_ _06742_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16281_ _02866_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__clkbuf_1
X_13493_ net98 decoded_imm\[9\] VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12593__S _06751_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_160_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_160_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_23_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18020_ clknet_leaf_105_clk _00027_ VGND VGND VPWR VPWR irq_pending\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15232_ cpuregs.regs\[8\]\[9\] cpuregs.regs\[9\]\[9\] cpuregs.regs\[10\]\[9\] cpuregs.regs\[11\]\[9\]
+ _01973_ _01974_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__mux4_1
X_12444_ _06705_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14384__B1 _08055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15163_ _03674_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__buf_6
XFILLER_0_152_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12375_ _06668_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16125__A1 _05413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09187__B _03916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10407__A reg_pc\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14114_ count_instr\[40\] _07843_ _07834_ VGND VGND VPWR VPWR _07846_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11326_ _05086_ _05944_ _03219_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15094_ _03656_ _01952_ _03674_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__a21o_1
XANTENNA_output261_A net261 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15409__S _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14045_ _07798_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__clkbuf_1
X_11257_ _05882_ _05885_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09789__S1 _04513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10208_ _04884_ _04888_ _04919_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__nand3_1
XANTENNA_output69_A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11188_ _03217_ _05825_ _05830_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17804_ clknet_leaf_56_clk _00973_ VGND VGND VPWR VPWR reg_pc\[12\] sky130_fd_sc_hd__dfxtp_1
X_10139_ _04018_ count_cycle\[53\] _04014_ count_cycle\[21\] _04853_ VGND VGND VPWR
+ VPWR _04854_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15996_ decoded_rd\[2\] _03636_ _02709_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__o21a_1
XFILLER_0_173_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17735_ clknet_leaf_96_clk _00904_ VGND VGND VPWR VPWR count_instr\[6\] sky130_fd_sc_hd__dfxtp_1
X_14947_ net208 net177 _01846_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__mux2_1
XANTENNA__12768__S _06880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17666_ clknet_leaf_16_clk _00835_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14878_ count_cycle\[60\] count_cycle\[61\] _01801_ _03240_ VGND VGND VPWR VPWR _01806_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16617_ cpuregs.regs\[1\]\[4\] _06124_ _03040_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13829_ cpuregs.regs\[0\]\[11\] VGND VGND VPWR VPWR _07654_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10288__S _04223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17597_ clknet_leaf_119_clk _00766_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12622__A0 _06184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09713__S1 _04219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16548_ _03008_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_151_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_151_clk sky130_fd_sc_hd__clkbuf_2
X_16479_ cpuregs.regs\[17\]\[3\] _06540_ _02968_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09020_ _03747_ _03781_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__nor2_1
X_18218_ clknet_leaf_92_clk _01289_ VGND VGND VPWR VPWR instr_rdcycleh sky130_fd_sc_hd__dfxtp_4
XFILLER_0_142_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11189__B1 _05829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09477__S0 _04207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18149_ clknet_leaf_70_clk alu_out\[23\] VGND VGND VPWR VPWR alu_out_q\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10400__A2 instr_maskirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09922_ cpuregs.regs\[20\]\[15\] cpuregs.regs\[21\]\[15\] cpuregs.regs\[22\]\[15\]
+ cpuregs.regs\[23\]\[15\] _04281_ _04470_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09853_ _04573_ _04574_ _04575_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__mux2_1
XANTENNA__15627__B1 _03657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08804_ _03482_ _03568_ _03569_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__o21ai_1
X_09784_ cpuregs.regs\[8\]\[11\] cpuregs.regs\[9\]\[11\] cpuregs.regs\[10\]\[11\]
+ cpuregs.regs\[11\]\[11\] _04282_ _04285_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__mux4_1
X_08735_ net101 net69 VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_1_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12678__S _06825_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13363__A _04036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_108 _07057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08666_ net91 net123 VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__or2_1
XANTENNA__10011__S1 _04478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_119 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08457__A reg_next_pc\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09609__A1 _04105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08597_ _03303_ _03254_ _03306_ _03375_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12613__A0 _06150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09704__S1 _04277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_142_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_142_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13302__S _07176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11611__A _06174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09218_ _03959_ _03955_ _03960_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__a21o_1
XANTENNA__09288__A instr_timer VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10490_ cpuregs.regs\[12\]\[31\] cpuregs.regs\[13\]\[31\] cpuregs.regs\[14\]\[31\]
+ cpuregs.regs\[15\]\[31\] _04329_ _04218_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__mux4_1
XANTENNA__15563__C1 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16107__A1 _03309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09149_ _03763_ _03880_ _03881_ _03904_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__a211o_1
XANTENNA__10927__B1 _05517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16613__S _03040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12160_ _06539_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08920__A _03662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11111_ _03441_ _05759_ _05784_ _03440_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_9_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11757__S _06258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09735__B decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12091_ _06125_ cpuregs.regs\[23\]\[4\] _06496_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ instr_sub _03582_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__nand2_1
XANTENNA__10155__A1 _04272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15850_ decoder_pseudo_trigger decoder_trigger VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _01752_ _01753_ _01754_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__and3b_1
XANTENNA__09751__A _04084_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15781_ _07778_ _07676_ _02571_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12993_ _07015_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14369__A _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17520_ clknet_leaf_130_clk _00689_ VGND VGND VPWR VPWR cpuregs.regs\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_14732_ _08362_ _08350_ _08363_ VGND VGND VPWR VPWR _08364_ sky130_fd_sc_hd__and3b_1
XANTENNA__10002__S1 _04473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11944_ cpuregs.waddr\[1\] cpuregs.waddr\[0\] VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_98_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08520__A1 _03297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17451_ clknet_leaf_131_clk _00620_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11505__B cpuregs.waddr\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11875_ _06082_ _06384_ _06081_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__and3b_4
X_14663_ _08308_ _08311_ VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__xnor2_1
XANTENNA_output107_A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16402_ _02930_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10826_ _03505_ _05502_ _03506_ _05390_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__o211a_1
X_13614_ _07462_ _07463_ VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__and2b_1
X_17382_ clknet_leaf_19_clk _00551_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14594_ _07958_ _07994_ _08248_ _07984_ VGND VGND VPWR VPWR _08249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16333_ _02893_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10836__S _05287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13545_ _07398_ _07399_ VGND VGND VPWR VPWR _07400_ sky130_fd_sc_hd__nand2_1
X_10757_ _03615_ _05452_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_41_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_133_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_133_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14357__B1 _07994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13476_ reg_pc\[7\] _07305_ _07335_ _07221_ VGND VGND VPWR VPWR _07336_ sky130_fd_sc_hd__a211o_1
X_16264_ reg_next_pc\[0\] _07778_ _02856_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10688_ _05300_ _03532_ _05338_ _05355_ _03607_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18003_ clknet_leaf_66_clk _01140_ VGND VGND VPWR VPWR irq_mask\[19\] sky130_fd_sc_hd__dfxtp_1
X_12427_ _06696_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15215_ cpuregs.regs\[8\]\[8\] cpuregs.regs\[9\]\[8\] cpuregs.regs\[10\]\[8\] cpuregs.regs\[11\]\[8\]
+ _01985_ _01986_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__mux4_2
XFILLER_0_125_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16195_ net257 net260 _01822_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_124_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16523__S _02990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15306__C1 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12358_ _06659_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15146_ cpuregs.regs\[8\]\[5\] cpuregs.regs\[9\]\[5\] cpuregs.regs\[10\]\[5\] cpuregs.regs\[11\]\[5\]
+ _01999_ _02000_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11667__S _06176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11309_ _05013_ _05930_ _03219_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__mux2_1
X_15077_ _03669_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__buf_6
X_12289_ _06622_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13332__A1 _04215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14028_ _07786_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09536__B1 _04265_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11343__A0 _05205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13096__A0 _06987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15979_ _04024_ _02635_ _02695_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__a21o_1
XANTENNA__15180__S1 _02023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13635__A2 _05261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09839__B2 instr_timer VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08520_ _03297_ _03299_ _03300_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__a21o_1
X_17718_ clknet_leaf_76_clk _00887_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dfxtp_1
XANTENNA__09934__S1 _04469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08451_ _03199_ mem_state\[0\] mem_state\[1\] _03234_ VGND VGND VPWR VPWR _03235_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17649_ clknet_leaf_47_clk _00818_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_77_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13911__A _07681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10746__S _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_124_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_124_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_98_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13122__S _07082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09003_ _03203_ _03752_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13571__A1 _04602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08740__A net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13358__A _07224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10481__S _04223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10480__S1 _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09905_ cpuregs.regs\[28\]\[14\] cpuregs.regs\[29\]\[14\] cpuregs.regs\[30\]\[14\]
+ cpuregs.regs\[31\]\[14\] _04290_ _04276_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10137__A1 _04391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09836_ _04328_ _04555_ _04559_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15076__A1 _05324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09767_ _04476_ _04482_ _04100_ _04492_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__a211o_2
XFILLER_0_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13093__A _07045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08718_ net106 net74 VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__nand2_1
XANTENNA__11637__A1 alu_out_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12834__A0 _06166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09698_ _04046_ _04419_ _04425_ _03225_ _04266_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__a221o_1
XANTENNA__11101__A3 _05044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11325__B _05943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08649_ timer\[4\] timer\[7\] timer\[3\] _03415_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__or4_1
XFILLER_0_84_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11660_ reg_pc\[16\] _06210_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__and2_1
XANTENNA__14636__B _07966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10611_ _05312_ _05313_ _05309_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11591_ _06156_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_115_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_115_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_153_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13032__S _07032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13330_ cpuregs.regs\[16\]\[0\] cpuregs.regs\[17\]\[0\] cpuregs.regs\[18\]\[0\] cpuregs.regs\[19\]\[0\]
+ _04207_ _04208_ VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__mux4_1
X_10542_ _05242_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13261_ _07157_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__clkbuf_1
X_10473_ _05113_ _05117_ _05118_ _05148_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__a31o_1
XANTENNA__16343__S _02896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12212_ _06574_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__clkbuf_1
X_15000_ _04227_ _04517_ _04525_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__or3_4
XFILLER_0_122_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09746__A _04280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13192_ _06947_ cpuregs.regs\[8\]\[2\] _07118_ VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12143_ _06328_ cpuregs.regs\[23\]\[29\] _06518_ VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16951_ clknet_leaf_53_clk _00079_ VGND VGND VPWR VPWR cpu_state\[5\] sky130_fd_sc_hd__dfxtp_2
X_12074_ _06491_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10128__A1 _04168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11025_ _03457_ _05221_ _05215_ _03459_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__a2bb2o_1
X_15902_ instr_xori _02618_ _02623_ _02643_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__a22o_1
X_16882_ _03185_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10223__S1 _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15067__A1 _03657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18621_ clknet_leaf_189_clk _01681_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09481__A _04206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15833_ decoded_imm_j\[18\] _05983_ _02596_ _02598_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__a211o_1
XANTENNA_output224_A net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13617__A2 _05260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11628__A1 alu_out_q\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18552_ clknet_leaf_3_clk _01617_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_15764_ _03423_ _02503_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__or2_2
X_12976_ _06335_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__buf_2
X_17503_ clknet_leaf_162_clk _00672_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14715_ _08352_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15930__B _02625_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18483_ clknet_leaf_155_clk _01548_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_11927_ _06413_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10300__A1 _04168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15695_ _04447_ _02506_ _02509_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_87_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17434_ clknet_leaf_112_clk _00603_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_14646_ _08232_ _07966_ _08290_ VGND VGND VPWR VPWR _08296_ sky130_fd_sc_hd__a21oi_1
X_11858_ _06375_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13450__B decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10809_ _05502_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17365_ clknet_leaf_164_clk _00534_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_106_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_106_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA_19 _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11789_ reg_out\[30\] alu_out_q\[30\] _06069_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14577_ _08232_ _07954_ _08226_ VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_172_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15790__A2 _03292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11251__A _04611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16316_ _06991_ cpuregs.regs\[15\]\[23\] _02881_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13528_ _07190_ _07381_ _07383_ VGND VGND VPWR VPWR _07384_ sky130_fd_sc_hd__or3_1
XFILLER_0_126_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17296_ clknet_leaf_165_clk _00470_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_191_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16247_ mem_rdata_q\[0\] _03783_ _03914_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13459_ _07190_ _07317_ _07319_ VGND VGND VPWR VPWR _07320_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_11_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput104 net104 VGND VGND VPWR VPWR cpi_rs2[14] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_93_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput115 net115 VGND VGND VPWR VPWR cpi_rs2[24] sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08560__A _03335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11564__A0 _06132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16178_ _02807_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__clkbuf_1
Xoutput126 net126 VGND VGND VPWR VPWR cpi_rs2[5] sky130_fd_sc_hd__buf_1
Xoutput137 net137 VGND VGND VPWR VPWR eoi[15] sky130_fd_sc_hd__buf_1
Xoutput148 net148 VGND VGND VPWR VPWR eoi[25] sky130_fd_sc_hd__buf_1
XFILLER_0_140_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15129_ _03719_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__buf_8
XANTENNA__16098__A3 _03916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput159 net159 VGND VGND VPWR VPWR eoi[6] sky130_fd_sc_hd__buf_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15393__A _03653_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09524__A3 _04255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09621_ _04258_ _04349_ _04350_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__or3b_2
XANTENNA__11426__A _03412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09552_ _04058_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12816__A0 _06078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12021__S _06460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08503_ mem_do_wdata VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__inv_2
XANTENNA__08496__B1 cpu_state\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12292__A1 _06571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09483_ _04214_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__buf_4
XANTENNA__15840__B _03979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12956__S _06985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16428__S _02943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13641__A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08434_ mem_state\[0\] mem_state\[1\] VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_144_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08735__A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08454__B _03237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13792__A1 _07304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13792__B2 reg_pc\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_159_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12691__S _06836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__14472__A _08035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08470__A _03252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10358__A1 _04231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08971__A1 mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15392__S1 _01937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09819_ count_instr\[12\] _04011_ _04017_ count_cycle\[44\] VGND VGND VPWR VPWR _04543_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_161_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10530__A1 _04602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_1010 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12830_ _06150_ cpuregs.regs\[6\]\[7\] _06906_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12761_ cpuregs.regs\[9\]\[7\] _06548_ _06869_ VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__mux2_1
XANTENNA__12866__S _06928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14500_ _08160_ _08156_ VGND VGND VPWR VPWR _08162_ sky130_fd_sc_hd__nor2_1
X_11712_ _06226_ reg_next_pc\[21\] _06262_ _06264_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__a211o_2
XFILLER_0_56_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10833__A2 _05440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12692_ _06838_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__clkbuf_1
X_15480_ cpuregs.regs\[4\]\[23\] cpuregs.regs\[5\]\[23\] cpuregs.regs\[6\]\[23\] cpuregs.regs\[7\]\[23\]
+ _01995_ _01937_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__mux4_1
XFILLER_0_83_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11643_ reg_pc\[14\] _06195_ _06093_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14431_ _08035_ _08092_ _08093_ _08095_ _08098_ VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__o32a_1
XANTENNA__13232__A0 _06987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15772__A2 _02486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12167__A _06131_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17150_ clknet_leaf_167_clk _00324_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11574_ _06141_ cpuregs.regs\[10\]\[6\] _06086_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__mux2_1
X_14362_ _03379_ _07984_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__nor2_4
Xinput17 irq[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10141__S0 _04282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 irq[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
XANTENNA__08885__S1 _03643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16101_ _03635_ _03799_ _03885_ _02755_ _02763_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__a41o_1
X_10525_ _03609_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__clkbuf_4
Xinput39 mem_rdata[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13313_ _07184_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__clkbuf_1
X_14293_ reg_next_pc\[31\] _05928_ _07944_ _07970_ VGND VGND VPWR VPWR _07971_ sky130_fd_sc_hd__o211a_2
X_17081_ clknet_leaf_13_clk _00255_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15909__C _02620_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13535__A1 _04419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15080__S0 _03669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09476__A _04074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16032_ decoded_imm\[5\] _02634_ _02727_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__a21o_1
X_13244_ _06999_ cpuregs.regs\[8\]\[27\] _07140_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__mux2_1
X_10456_ cpuregs.regs\[0\]\[30\] cpuregs.regs\[1\]\[30\] cpuregs.regs\[2\]\[30\] cpuregs.regs\[3\]\[30\]
+ _04477_ _04478_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11010__A2 _05213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08411__B1 _03195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13175_ _07111_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12106__S _06507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10387_ cpuregs.regs\[16\]\[28\] cpuregs.regs\[17\]\[28\] cpuregs.regs\[18\]\[28\]
+ cpuregs.regs\[19\]\[28\] _04273_ _04283_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__mux4_1
XANTENNA__16801__S _03138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08962__A1 _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12126_ _06519_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__clkbuf_1
X_17983_ clknet_leaf_63_clk _01120_ VGND VGND VPWR VPWR irq_active sky130_fd_sc_hd__dfxtp_4
XANTENNA__15383__S1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13726__A _05013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12057_ _06257_ cpuregs.regs\[22\]\[20\] _06482_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__mux2_1
X_16934_ clknet_leaf_101_clk _00115_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16237__A0 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11008_ _04945_ _04913_ _04880_ _04848_ _05264_ _05232_ VGND VGND VPWR VPWR _05689_
+ sky130_fd_sc_hd__mux4_1
X_16865_ _06580_ cpuregs.regs\[14\]\[22\] _03174_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__mux2_1
XANTENNA__11246__A _04602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18604_ clknet_leaf_99_clk _01669_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15941__A mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15816_ _03826_ _06016_ _02587_ _03987_ _02591_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__a221o_1
X_16796_ _03140_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15460__A1 decoded_imm\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18535_ clknet_leaf_156_clk _01600_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_15747_ _02476_ _02546_ _02547_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__or3b_1
XANTENNA__12776__S _06880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12959_ _06993_ cpuregs.regs\[31\]\[24\] _06985_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18466_ clknet_leaf_137_clk _01531_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08555__A _03330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15678_ _01872_ _02479_ _02495_ _02496_ _07775_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_173_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_54 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09690__A2 _04397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17417_ clknet_leaf_186_clk _00586_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10296__S _04321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14629_ _08269_ _08272_ _08280_ VGND VGND VPWR VPWR _08281_ sky130_fd_sc_hd__a21oi_1
X_18397_ clknet_leaf_183_clk _01462_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10037__B1 _04202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13774__A1 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17348_ clknet_leaf_180_clk _00517_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15515__A2 _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17279_ clknet_leaf_176_clk _00453_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09825__S0 _04216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15279__A1 _02012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08953__A1 _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08983_ mem_rdata_q\[13\] net37 _03208_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11855__S _06370_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15126__S1 _01980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09604_ _04289_ _04327_ _04333_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15851__A _02610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14254__A2 irq_state\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09535_ _04048_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_104_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12686__S _06825_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09466_ net35 net52 _04039_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10815__A2 _05440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08417_ _03193_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__clkbuf_4
X_09397_ _04052_ _04130_ _04080_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10028__B1 _04673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10579__A1 _04036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09433__A2 _04104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10674__S1 _05244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10310_ _05018_ _05019_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__xor2_1
XANTENNA__13310__S _07176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11290_ reg_next_pc\[22\] reg_out\[22\] _05898_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__mux2_2
XFILLER_0_104_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10241_ _04884_ _04952_ _04917_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__o21a_1
XANTENNA__16621__S _03040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10426__S1 _04469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12740__A2 _06862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10172_ _04884_ _04885_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_163_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15365__S1 _02014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14980_ _01862_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__16219__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15690__A1 _04415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13931_ _03330_ _07704_ _07705_ net138 VGND VGND VPWR VPWR _07719_ sky130_fd_sc_hd__a22o_1
XANTENNA__15117__S1 _01971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10503__B2 _05207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16650_ _03039_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__buf_6
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13862_ _07670_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15442__A1 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15601_ cpuregs.regs\[12\]\[30\] cpuregs.regs\[13\]\[30\] cpuregs.regs\[14\]\[30\]
+ cpuregs.regs\[15\]\[30\] _03641_ _03684_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__mux4_1
X_12813_ _06081_ _06082_ _06083_ cpuregs.waddr\[2\] VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_158_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16581_ _03025_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13793_ _07626_ _07629_ _07630_ _07284_ VGND VGND VPWR VPWR _07631_ sky130_fd_sc_hd__o22a_1
XANTENNA__13453__B1 _03631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18320_ clknet_leaf_37_clk _01388_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15532_ cpuregs.regs\[16\]\[26\] cpuregs.regs\[17\]\[26\] cpuregs.regs\[18\]\[26\]
+ cpuregs.regs\[19\]\[26\] _01995_ _01937_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__mux4_1
X_12744_ cpuregs.waddr\[2\] _06862_ _06867_ _06861_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ clknet_leaf_22_clk _01322_ VGND VGND VPWR VPWR decoded_imm\[9\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_155_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ cpuregs.regs\[16\]\[22\] cpuregs.regs\[17\]\[22\] cpuregs.regs\[18\]\[22\]
+ cpuregs.regs\[19\]\[22\] _02030_ _02031_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__mux4_1
XFILLER_0_166_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12675_ _06829_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17202_ clknet_leaf_111_clk _00376_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__14953__A0 net211 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14414_ decoded_imm_j\[9\] _07925_ VGND VGND VPWR VPWR _08083_ sky130_fd_sc_hd__or2_1
XFILLER_0_170_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13756__B2 reg_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ reg_pc\[11\] reg_pc\[10\] _06162_ reg_pc\[12\] VGND VGND VPWR VPWR _06188_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18182_ clknet_leaf_32_clk _01253_ VGND VGND VPWR VPWR instr_jal sky130_fd_sc_hd__dfxtp_4
X_15394_ cpuregs.regs\[16\]\[18\] cpuregs.regs\[17\]\[18\] cpuregs.regs\[18\]\[18\]
+ cpuregs.regs\[19\]\[18\] _01936_ _01937_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10114__S0 _04275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17133_ clknet_leaf_123_clk _00307_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14345_ _08007_ _08010_ VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09918__B decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11557_ _06126_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11510__A_N cpuregs.waddr\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08822__B net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15001__A _01881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10508_ instr_and instr_andi VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__or2_1
X_17064_ clknet_leaf_144_clk _00238_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_output99_A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11488_ _06054_ irq_pending\[31\] _06063_ net25 VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__a31o_1
X_14276_ reg_pc\[24\] _07953_ _07959_ _07960_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09188__A1 _03763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09188__B2 _03810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16015_ instr_jal VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__buf_2
X_10439_ _05119_ _05142_ _05145_ _04007_ irq_pending\[29\] VGND VGND VPWR VPWR _08390_
+ sky130_fd_sc_hd__o32a_1
X_13227_ _06982_ cpuregs.regs\[8\]\[19\] _07129_ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16531__S _02990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13158_ _07102_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15356__S1 _02014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12109_ _06510_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__clkbuf_1
X_13089_ _06980_ cpuregs.regs\[7\]\[18\] _07057_ VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__mux2_1
X_17966_ clknet_leaf_0_clk _01103_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15681__A1 _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14484__A2 _07948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16917_ clknet_leaf_10_clk _00098_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11298__A2 _05829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17897_ clknet_leaf_95_clk _01066_ VGND VGND VPWR VPWR count_cycle\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16848_ _06563_ cpuregs.regs\[14\]\[14\] _03163_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13444__B1 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16779_ _03131_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_1010 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09320_ _00069_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__clkbuf_8
X_18518_ clknet_leaf_188_clk _01583_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10258__B1 _04237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10353__S0 _04207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09251_ _03737_ _03844_ _03927_ _03990_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_173_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11423__B irq_mask\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18449_ clknet_leaf_115_clk _01514_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16706__S _03087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13747__A1 _07209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15292__S0 _01985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13747__B2 reg_pc\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09182_ _03739_ _03749_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__and2_2
XFILLER_0_133_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_78_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08732__B net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13130__S _07082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15595__S1 _02037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15932__A_N mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16449__A0 _06987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15347__S1 _02000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08966_ _03727_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_87_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15672__A1 _04185_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11289__A2 _05829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13683__B1 _03311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08897_ _00065_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_95_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_86_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_162_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14197__A _07904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10249__B1 _04017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09518_ _04248_ _04249_ _03384_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__and3b_1
XFILLER_0_67_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10790_ _05285_ _05484_ _05244_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10344__S0 _04758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09449_ _04180_ _04181_ _04063_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_96_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12460_ _06383_ _06713_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__nand2_4
XFILLER_0_35_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08923__A _03666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11411_ _03826_ _06016_ _05996_ _06018_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12391_ _06676_ _06532_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__nor2_4
XFILLER_0_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13040__S _07032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11342_ _05954_ _05957_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__xor2_1
X_14130_ count_instr\[45\] VGND VGND VPWR VPWR _07857_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15586__S1 _03684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10972__B2 _05440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14061_ count_instr\[23\] _07805_ count_instr\[24\] VGND VGND VPWR VPWR _07809_ sky130_fd_sc_hd__a21o_1
X_11273_ _05901_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16351__S _02896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14660__A _08232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08917__A1 _03638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13012_ _07025_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__clkbuf_1
X_10224_ _04935_ _04936_ _04064_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15338__S1 _01980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17820_ clknet_leaf_67_clk _00989_ VGND VGND VPWR VPWR reg_pc\[28\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__13276__A _07153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10155_ _04272_ _04865_ _04869_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15663__A1 _04101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17751_ clknet_leaf_85_clk _00920_ VGND VGND VPWR VPWR count_instr\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14963_ irq_delay irq_active _07755_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__mux2_1
X_10086_ _04328_ _04802_ _04237_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_86_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16702_ _06968_ cpuregs.regs\[19\]\[12\] _03087_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__mux2_1
X_13914_ _07707_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17682_ clknet_leaf_156_clk _00851_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_14894_ _01817_ _07277_ _07284_ _01818_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_18_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15415__A1 _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14819__B _01753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16633_ _03053_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__clkbuf_1
X_13845_ cpuregs.regs\[0\]\[19\] VGND VGND VPWR VPWR _07662_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15510__S1 _01986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13215__S _07129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16564_ _06966_ cpuregs.regs\[18\]\[11\] _03015_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__mux2_1
X_13776_ _04959_ _07236_ _07614_ VGND VGND VPWR VPWR _07615_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_69_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10988_ _05418_ _05622_ _05600_ _05562_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_58_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18303_ clknet_leaf_6_clk _01371_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15515_ net115 _01905_ _02349_ _02350_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__o22a_1
XANTENNA__15179__B1 _02017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12727_ _06856_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11452__A2 irq_pending\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16495_ _02980_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15274__S0 _02085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14926__A0 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18234_ clknet_leaf_9_clk _01305_ VGND VGND VPWR VPWR cpuregs.raddr1\[2\] sky130_fd_sc_hd__dfxtp_1
X_15446_ cpuregs.regs\[4\]\[21\] cpuregs.regs\[5\]\[21\] cpuregs.regs\[6\]\[21\] cpuregs.regs\[7\]\[21\]
+ _01979_ _01980_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__mux4_1
X_12658_ _06819_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11609_ _06171_ _06172_ _06075_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__o21a_1
X_18165_ clknet_leaf_32_clk _01236_ VGND VGND VPWR VPWR decoded_imm_j\[6\] sky130_fd_sc_hd__dfxtp_1
X_15377_ _02218_ _02219_ _01907_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12589_ cpuregs.regs\[2\]\[28\] _06592_ _06774_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17116_ clknet_leaf_12_clk _00290_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14328_ _07908_ _08003_ VGND VGND VPWR VPWR _08004_ sky130_fd_sc_hd__nor2_1
X_18096_ clknet_leaf_92_clk _01200_ VGND VGND VPWR VPWR timer\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15577__S1 _01997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17047_ clknet_leaf_169_clk _00221_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14259_ _05857_ _06245_ VGND VGND VPWR VPWR _07949_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08908__A1 _03664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13901__A1 _03349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09664__A reg_pc\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09030__A0 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15329__S1 _02070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08820_ _03454_ _03455_ _03585_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09581__A1 _03385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15103__B1 decoded_imm\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_360 VGND VGND VPWR VPWR alphacore_360/HI trace_data[21] sky130_fd_sc_hd__conb_1
Xalphacore_371 VGND VGND VPWR VPWR alphacore_371/HI trace_data[32] sky130_fd_sc_hd__conb_1
X_08751_ net128 VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__inv_2
X_17949_ clknet_leaf_77_clk _08390_ VGND VGND VPWR VPWR reg_out\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_77_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_68_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08682_ net118 net86 VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__nand2_1
XANTENNA__11140__A1 _03407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15406__A1 _03692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11140__B2 _04422_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09884__A2 _04008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11691__A2 _03358_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15501__S1 _01992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09303_ _03242_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08446__C _03191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14745__A _01714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16436__S _02943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14917__A0 net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15265__S0 _01985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09234_ _03837_ _03966_ _03975_ _03888_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08743__A net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14464__B _07934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09165_ _03908_ _03915_ _03917_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09096_ _03816_ _03770_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_151_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10954__A1 _05361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15568__S1 _02031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15893__B2 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11903__A0 _06193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10706__B2 _05404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10513__A _05211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09998_ reg_pc\[16\] decoded_imm\[16\] _04683_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__a21o_1
XANTENNA__11328__B _05943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08949_ cpuregs.regs\[0\]\[4\] cpuregs.regs\[1\]\[4\] cpuregs.regs\[2\]\[4\] cpuregs.regs\[3\]\[4\]
+ _03661_ _03662_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_4_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_68_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_4_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12150__D _06083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11960_ _06431_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16200__A _03730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13543__B decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10911_ _05598_ _05571_ _05543_ _05510_ _05286_ _05413_ VGND VGND VPWR VPWR _05599_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_168_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11682__A2 _03336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11891_ _06394_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16070__A1 decoded_imm\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13630_ _07254_ _07477_ _07478_ _07217_ VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__a22o_1
XANTENNA__16070__B2 mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10842_ _05500_ _05532_ _05533_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13561_ _03275_ _07410_ _07414_ VGND VGND VPWR VPWR _07415_ sky130_fd_sc_hd__a21o_1
XANTENNA__12874__S _06928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11434__A2 irq_pending\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10773_ _03549_ _05468_ _05363_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14655__A _07998_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15300_ _02020_ _02139_ _02147_ _01960_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__o211a_4
X_12512_ _06289_ cpuregs.regs\[28\]\[24\] _06737_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16280_ _06955_ cpuregs.regs\[15\]\[6\] _02859_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13492_ net98 decoded_imm\[9\] VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_136_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15231_ cpuregs.regs\[12\]\[9\] cpuregs.regs\[13\]\[9\] cpuregs.regs\[14\]\[9\] cpuregs.regs\[15\]\[9\]
+ _01970_ _01971_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12443_ cpuregs.regs\[27\]\[24\] _06584_ _06700_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__mux2_1
XANTENNA__15581__B1 _02197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15162_ _02012_ _02015_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__or2_1
XANTENNA__11510__C _06082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12374_ cpuregs.regs\[26\]\[24\] _06584_ _06663_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10407__B decoded_imm\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14113_ count_instr\[40\] _07843_ VGND VGND VPWR VPWR _07845_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11325_ _05938_ _05943_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__xor2_1
XFILLER_0_50_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15093_ _01950_ _01951_ _03713_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__mux2_1
XANTENNA__14390__A decoded_imm_j\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09484__A _04055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14044_ _07796_ _07778_ _07797_ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__and3b_1
X_11256_ _05887_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15884__B2 is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10207_ _04884_ _04888_ _04919_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__a21o_1
XANTENNA__11519__A _03195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11187_ _03217_ _05825_ _05830_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__and3_1
XANTENNA__12114__S _06507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10138_ count_instr\[53\] _04016_ _04012_ count_instr\[21\] VGND VGND VPWR VPWR _04853_
+ sky130_fd_sc_hd__a22o_1
X_17803_ clknet_leaf_56_clk _00972_ VGND VGND VPWR VPWR reg_pc\[11\] sky130_fd_sc_hd__dfxtp_2
X_15995_ _03885_ _03880_ _02702_ _03826_ _05973_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_59_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__11953__S _06424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09315__B2 _04050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_max_cap300_A net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17734_ clknet_leaf_96_clk _00903_ VGND VGND VPWR VPWR count_instr\[5\] sky130_fd_sc_hd__dfxtp_1
X_10069_ _04784_ _04785_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__xnor2_1
X_14946_ _01848_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11122__A1 _05361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17665_ clknet_leaf_188_clk _00834_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_14877_ _01804_ _01805_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__nor2_1
XANTENNA__11673__A2 _03348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16061__A1 decoded_imm\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10881__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16616_ _03044_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__clkbuf_1
X_13828_ _07653_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17596_ clknet_leaf_105_clk _00765_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16547_ _06949_ cpuregs.regs\[18\]\[3\] _03004_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__mux2_1
X_13759_ _07578_ _07581_ _07598_ VGND VGND VPWR VPWR _07599_ sky130_fd_sc_hd__and3_1
XANTENNA__12784__S _06880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08921__S0 _03641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16478_ _02971_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18217_ clknet_leaf_102_clk _01288_ VGND VGND VPWR VPWR instr_rdcycle sky130_fd_sc_hd__dfxtp_1
X_15429_ _02269_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14375__A1 _06863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09378__B decoded_imm\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09477__S1 _04208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18148_ clknet_leaf_70_clk alu_out\[22\] VGND VGND VPWR VPWR alu_out_q\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18079_ clknet_leaf_47_clk _01184_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09921_ net73 VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14623__A1_N _08012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09852_ _04320_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_111_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15627__A1 _00068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08803_ net108 net76 VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__or2b_1
X_09783_ cpuregs.regs\[12\]\[11\] cpuregs.regs\[13\]\[11\] cpuregs.regs\[14\]\[11\]
+ cpuregs.regs\[15\]\[11\] _04282_ _04285_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__mux4_1
XANTENNA__12959__S _06985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15843__B _03885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11863__S _06370_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08734_ net101 VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11113__A1 _05363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13363__B decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_109 decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08665_ instr_beq _03430_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__nor2_1
XANTENNA__11664__A2 _03330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08457__B _03199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15486__S0 _03645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16052__B2 _03940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08596_ _03248_ _03308_ _03374_ _03249_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14475__A decoded_imm_j\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15238__S0 _01982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09217_ _03818_ _03776_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__nor2_2
XFILLER_0_107_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09288__B instr_maskirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_588 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09148_ _03883_ _03884_ _03903_ _03878_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__o31a_1
XANTENNA__16107__A2 _03255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08596__A2 _03308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09079_ _03737_ _03751_ _03778_ _03840_ _03758_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__a32o_1
X_11110_ net120 _05143_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_15_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15866__B2 _02623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12090_ _06500_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__clkbuf_1
X_11041_ _03458_ _05709_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_168_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10243__A reg_pc\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16815__A0 _06598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13629__A0 _04611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14800_ count_cycle\[34\] _01748_ count_cycle\[35\] VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__a21o_1
XANTENNA__15245__S _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _06186_ _03298_ _03409_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__a21o_1
X_12992_ cpuregs.regs\[3\]\[4\] _06542_ _07010_ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__mux2_1
XANTENNA__09848__A2 _04016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14731_ count_cycle\[13\] _08359_ count_cycle\[14\] VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__a21o_1
X_11943_ _06421_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11655__A2 _03356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16043__A1 decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17450_ clknet_leaf_183_clk _00619_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14662_ _08309_ _08310_ VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11874_ cpuregs.waddr\[2\] _06083_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_28_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _07007_ cpuregs.regs\[16\]\[31\] _02895_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__mux2_1
X_13613_ _07445_ _07450_ _07461_ VGND VGND VPWR VPWR _07463_ sky130_fd_sc_hd__a21o_1
X_10825_ _03507_ _05499_ _03553_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__o21bai_1
X_17381_ clknet_leaf_187_clk _00550_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14593_ _08246_ _08247_ VGND VGND VPWR VPWR _08248_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16332_ _07007_ cpuregs.regs\[15\]\[31\] _02858_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__mux2_1
X_13544_ net70 decoded_imm\[12\] VGND VGND VPWR VPWR _07399_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09479__A _04078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10756_ _03615_ _05452_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_41_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10091__A1 _04271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14357__A1 _07986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16263_ _05941_ _07944_ _03292_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__a21o_1
X_13475_ _03387_ _04382_ VGND VGND VPWR VPWR _07335_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10687_ _05361_ _05365_ _05366_ _05387_ VGND VGND VPWR VPWR alu_out\[3\] sky130_fd_sc_hd__a31o_2
XANTENNA__10418__A _04054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18002_ clknet_leaf_66_clk _01139_ VGND VGND VPWR VPWR irq_mask\[18\] sky130_fd_sc_hd__dfxtp_1
X_15214_ _03709_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__buf_6
X_12426_ cpuregs.regs\[27\]\[16\] _06567_ _06689_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16194_ net297 _01822_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15145_ _03647_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__buf_8
XFILLER_0_23_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12357_ cpuregs.regs\[26\]\[16\] _06567_ _06652_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08830__B net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output81_A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15401__S0 _03645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11308_ _05925_ _05929_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_39_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15076_ _05324_ _01906_ _01930_ _01935_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__o22a_1
X_12288_ cpuregs.regs\[25\]\[16\] _06567_ _06615_ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09536__B2 _03225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14027_ _07784_ _07778_ _07785_ VGND VGND VPWR VPWR _07786_ sky130_fd_sc_hd__and3b_1
XANTENNA__15944__A mem_rdata_q\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11239_ _05872_ _05873_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_56_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15887__C_N _02613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15978_ _02645_ mem_rdata_q\[26\] mem_rdata_q\[27\] _02690_ VGND VGND VPWR VPWR _02695_
+ sky130_fd_sc_hd__and4bb_2
XFILLER_0_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10529__S0 _05230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14293__B1 _07944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09839__A2 _04308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17717_ clknet_leaf_76_clk _00886_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dfxtp_1
X_14929_ _01839_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09395__S0 _04071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11646__A2 _03353_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16034__B2 mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08450_ mem_do_wdata mem_do_rdata _03199_ _03227_ _03233_ VGND VGND VPWR VPWR _03234_
+ sky130_fd_sc_hd__o311a_1
X_17648_ clknet_leaf_49_clk _00817_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_19_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17579_ clknet_leaf_131_clk _00748_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14295__A _06863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09472__B1 _04145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14348__A1 reg_next_pc\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10328__A _04051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16714__S _03087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12019__S _06460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09002_ _03231_ _03755_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09224__A0 mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09775__A1 irq_pending\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09775__B2 _03385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08740__B net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16015__A instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15639__B1_N irq_state\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09904_ cpuregs.regs\[24\]\[14\] cpuregs.regs\[25\]\[14\] cpuregs.regs\[26\]\[14\]
+ cpuregs.regs\[27\]\[14\] _04290_ _04276_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__mux4_1
XANTENNA__15854__A _02612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09852__A _04320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09835_ _04068_ _04558_ _04081_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__a21o_1
XANTENNA__12689__S _06836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15076__A2 _01906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09766_ _04483_ _04486_ _04491_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14284__B1 _07944_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08468__A instr_timer VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08717_ net106 net74 VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__or2_1
X_09697_ _04420_ _04424_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16025__A1 decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08648_ timer\[5\] timer\[6\] timer\[1\] timer\[2\] VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14587__A1 _07954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08579_ irq_mask\[19\] irq_pending\[19\] VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__and2b_2
XFILLER_0_138_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10610_ net86 net87 _05263_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11590_ _06075_ _06152_ _06155_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_1007 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11270__A0 reg_next_pc\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10541_ _05233_ _05234_ _05238_ _05241_ _05243_ _05244_ VGND VGND VPWR VPWR _05245_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13260_ _06947_ cpuregs.regs\[5\]\[2\] _07154_ VGND VGND VPWR VPWR _07157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10472_ _04391_ _05150_ _05177_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11022__A0 _04959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12211_ cpuregs.regs\[24\]\[19\] _06573_ _06555_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__mux2_1
XANTENNA__09766__A1 _04483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13191_ _07120_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12142_ _06527_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__clkbuf_1
X_16950_ clknet_leaf_53_clk _00078_ VGND VGND VPWR VPWR cpu_state\[4\] sky130_fd_sc_hd__dfxtp_1
X_12073_ _06320_ cpuregs.regs\[22\]\[28\] _06482_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__mux2_1
XANTENNA__10128__A2 _04842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12522__A0 _06328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11024_ _05288_ _05399_ _05703_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__and3_1
X_15901_ instr_sltiu _02618_ _02643_ _02644_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__a22o_1
X_16881_ _06596_ cpuregs.regs\[14\]\[30\] _03151_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__mux2_1
XANTENNA__12599__S _06788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18620_ clknet_leaf_17_clk _01680_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15832_ _05969_ _03634_ _03918_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_144_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15763_ _02477_ _02558_ _02559_ _02545_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__o211a_1
X_18551_ clknet_leaf_11_clk _01616_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12975_ _07004_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output217_A net217 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14714_ _08349_ _08350_ _08351_ VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__and3b_1
X_17502_ clknet_leaf_118_clk _00671_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_18482_ clknet_leaf_128_clk _01547_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_11926_ _06281_ cpuregs.regs\[20\]\[23\] _06409_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__mux2_1
X_15694_ _02484_ _02507_ _02508_ _03240_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__a31o_1
XANTENNA__10300__A2 _05009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17433_ clknet_leaf_114_clk _00602_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_14645_ _08221_ _07967_ VGND VGND VPWR VPWR _08295_ sky130_fd_sc_hd__xnor2_1
X_11857_ _06289_ cpuregs.regs\[11\]\[24\] _06370_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13223__S _07129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10808_ _05500_ _05501_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__and2_1
X_17364_ clknet_leaf_122_clk _00533_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14576_ _08221_ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__buf_4
X_11788_ _06330_ _06331_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10064__A1 _04156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16315_ _02884_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13527_ _04360_ _07315_ _07382_ _07216_ VGND VGND VPWR VPWR _07383_ sky130_fd_sc_hd__o211a_1
XANTENNA__11251__B _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15939__A mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10739_ _05246_ _05335_ _05423_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__o21a_1
X_17295_ clknet_leaf_119_clk _00469_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15622__S0 _03645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16246_ _02847_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__clkbuf_1
X_13458_ _04360_ _05227_ _07318_ _07237_ VGND VGND VPWR VPWR _07319_ sky130_fd_sc_hd__o211a_1
XANTENNA__08841__A net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14562__B _07954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12409_ cpuregs.regs\[27\]\[8\] _06550_ _06678_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16177_ net282 net244 _02797_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__mux2_1
Xoutput105 net105 VGND VGND VPWR VPWR cpi_rs2[15] sky130_fd_sc_hd__clkbuf_1
X_13389_ _07237_ VGND VGND VPWR VPWR _07254_ sky130_fd_sc_hd__clkbuf_4
Xoutput116 net116 VGND VGND VPWR VPWR cpi_rs2[25] sky130_fd_sc_hd__buf_1
XANTENNA__08560__B _03336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput127 net127 VGND VGND VPWR VPWR cpi_rs2[6] sky130_fd_sc_hd__buf_1
Xoutput138 net138 VGND VGND VPWR VPWR eoi[16] sky130_fd_sc_hd__clkbuf_1
X_15128_ _01972_ _01975_ _01978_ _01981_ _01982_ _03639_ VGND VGND VPWR VPWR _01983_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput149 net149 VGND VGND VPWR VPWR eoi[26] sky130_fd_sc_hd__buf_1
X_15059_ _03671_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_71_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16255__A1 _03885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09620_ _04246_ _04247_ _04259_ _04256_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__a211o_1
XANTENNA__14266__B1 _07942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09551_ _04281_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__buf_6
XANTENNA__11619__A2 reg_next_pc\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08502_ _03239_ _03258_ _03282_ _03284_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08496__A1 _03218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09482_ _04068_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15840__C _03864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13641__B decoded_imm\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08433_ _03192_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__buf_4
XANTENNA__16471__A_N cpuregs.waddr\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08735__B net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13777__C1 _07232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13792__A2 _05139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16444__S _02943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13529__C1 _07221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15613__S0 _01995_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08751__A net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11004__B1 _05215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_975 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10492__S _04222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_148_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16494__A1 _06554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12504__A0 _06257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13308__S _07176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09818_ _04538_ _04540_ _04541_ _04537_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__a31o_1
XANTENNA__10521__A _05218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10530__A2 _04611_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09749_ _04471_ _04474_ _04430_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__mux2_1
XANTENNA__10240__B decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16619__S _03040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12760_ _06876_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09684__B1 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11711_ _06252_ _03346_ _06253_ _06263_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__a22o_1
XANTENNA__15757__B1 _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12691_ _06184_ cpuregs.regs\[12\]\[11\] _06836_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14430_ _08082_ _08087_ _08094_ _08096_ _08097_ VGND VGND VPWR VPWR _08098_ sky130_fd_sc_hd__a311o_1
X_11642_ _06202_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14361_ _07960_ _07915_ _07992_ _08034_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09987__B2 _04010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11573_ _06140_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__buf_2
XFILLER_0_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput18 irq[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16100_ _02762_ _05976_ _05973_ is_alu_reg_imm VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10141__S1 _04285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15604__S0 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13312_ _06999_ cpuregs.regs\[5\]\[27\] _07176_ VGND VGND VPWR VPWR _07184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10524_ _05226_ _05227_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__nor2_4
XFILLER_0_135_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 irq[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_2
X_17080_ clknet_leaf_176_clk _00254_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09757__A _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14292_ _05941_ _06340_ VGND VGND VPWR VPWR _07970_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08661__A _03412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16031_ instr_jal decoded_imm_j\[5\] _02610_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__and3_1
XANTENNA__15080__S1 _03646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13243_ _07147_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12183__A _06533_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10455_ cpuregs.regs\[4\]\[30\] cpuregs.regs\[5\]\[30\] cpuregs.regs\[6\]\[30\] cpuregs.regs\[7\]\[30\]
+ _04232_ _04233_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12743__A0 _06186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13174_ _06997_ cpuregs.regs\[4\]\[26\] _07104_ VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__mux2_1
X_10386_ cpuregs.regs\[20\]\[28\] cpuregs.regs\[21\]\[28\] cpuregs.regs\[22\]\[28\]
+ cpuregs.regs\[23\]\[28\] _04273_ _04283_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_107_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12125_ _06257_ cpuregs.regs\[23\]\[20\] _06518_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__mux2_1
X_17982_ clknet_leaf_63_clk _01119_ VGND VGND VPWR VPWR irq_delay sky130_fd_sc_hd__dfxtp_1
XANTENNA__12911__A _06165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13726__B decoded_imm\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16933_ clknet_leaf_179_clk _00114_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_12056_ _06459_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__buf_6
X_11007_ _05597_ _05674_ _05681_ _05688_ VGND VGND VPWR VPWR alu_out\[22\] sky130_fd_sc_hd__a211o_1
XANTENNA__09911__B2 _04187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12122__S _06507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16864_ _03176_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14407__A1_N _08035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18603_ clknet_leaf_99_clk _01668_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[20\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11246__B _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15941__B mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15815_ decoded_imm_j\[8\] _05973_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__and2_1
X_16795_ _06578_ cpuregs.regs\[13\]\[21\] _03138_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__mux2_1
XANTENNA__16529__S _02990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11961__S _06424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15460__A2 _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13742__A _05013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15746_ timer\[23\] timer\[22\] _02540_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__or3_2
X_18534_ clknet_leaf_144_clk _01599_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12958_ _06288_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_116_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10285__A1 _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11482__B1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11909_ _06216_ cpuregs.regs\[20\]\[15\] _06398_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18465_ clknet_leaf_157_clk _01530_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_15677_ timer\[5\] _02493_ _02488_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__a21oi_1
X_12889_ _06946_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09427__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17416_ clknet_leaf_173_clk _00585_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14628_ _08221_ _07964_ VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18396_ clknet_leaf_173_clk _01461_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10037__A1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11234__A0 _04532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10037__B2 irq_pending\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17347_ clknet_leaf_18_clk _00516_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14559_ _08121_ _08210_ _08211_ _08216_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17278_ clknet_leaf_17_clk _00452_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08571__A _03346_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16229_ net48 mem_16bit_buffer\[7\] _02831_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09825__S1 _04376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08982_ mem_rdata_q\[29\] net54 _03208_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09589__S0 _04274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13128__S _07082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10341__A reg_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09603_ _04328_ _04332_ _04237_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__a21o_1
XANTENNA__15987__B1 _03864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13652__A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09534_ net60 net258 _04035_ net46 _04264_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_104_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08746__A _03509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09465_ net92 VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08416_ net40 mem_rdata_q\[16\] _03200_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09396_ _04128_ _04129_ _00071_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10028__B2 _04746_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09577__A instr_maskirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10516__A _05215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10240_ reg_pc\[23\] decoded_imm\[23\] VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_991 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10200__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10171_ reg_pc\[22\] decoded_imm\[22\] VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_163_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16203__A _03218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15675__C1 _07775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13038__S _07032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13930_ _07718_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15690__A2 _02486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13861_ cpuregs.regs\[0\]\[27\] VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_141_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_190_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16349__S _02896_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15600_ _02428_ _02429_ _01907_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12812_ _06903_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__clkbuf_1
X_16580_ _06982_ cpuregs.regs\[18\]\[19\] _03015_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__mux2_1
X_13792_ _07304_ _05139_ _07305_ reg_pc\[29\] VGND VGND VPWR VPWR _07630_ sky130_fd_sc_hd__a22o_1
XANTENNA__09657__B1 _03252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14650__B1 _07967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15531_ net116 _01905_ _02364_ _02365_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11464__B1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12743_ _06186_ decoded_rd\[2\] _06863_ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18250_ clknet_leaf_22_clk _01321_ VGND VGND VPWR VPWR decoded_imm\[8\] sky130_fd_sc_hd__dfxtp_4
X_15462_ cpuregs.regs\[20\]\[22\] cpuregs.regs\[21\]\[22\] cpuregs.regs\[22\]\[22\]
+ cpuregs.regs\[23\]\[22\] _01979_ _01980_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_13_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12674_ _06114_ cpuregs.regs\[12\]\[3\] _06825_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11216__A0 _04419_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17201_ clknet_leaf_160_clk _00375_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14413_ decoded_imm_j\[9\] _07925_ VGND VGND VPWR VPWR _08082_ sky130_fd_sc_hd__nand2_1
XANTENNA__14953__A1 net180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ reg_pc\[12\] reg_pc\[11\] _06171_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18181_ clknet_leaf_31_clk _01252_ VGND VGND VPWR VPWR instr_auipc sky130_fd_sc_hd__dfxtp_1
X_15393_ _03653_ _02234_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_139_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10114__S1 _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17132_ clknet_leaf_149_clk _00306_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09487__A _04218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14344_ _08017_ _08018_ VGND VGND VPWR VPWR _08019_ sky130_fd_sc_hd__or2_1
X_11556_ _06125_ cpuregs.regs\[10\]\[4\] _06086_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10507_ _05209_ _05210_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__nand2_1
X_17063_ clknet_leaf_147_clk _00237_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15902__B1 _02623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14275_ _03294_ VGND VGND VPWR VPWR _07960_ sky130_fd_sc_hd__buf_4
X_11487_ irq_mask\[31\] _03428_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16014_ mem_rdata_q\[21\] _02712_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__and2_1
XANTENNA__08470__C_N _03253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13226_ _07138_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__clkbuf_1
X_10438_ _03680_ _05143_ _04752_ _05144_ _04202_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15428__S _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13737__A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13157_ _06980_ cpuregs.regs\[4\]\[18\] _07093_ VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__mux2_1
X_10369_ _04046_ _05076_ _04752_ _05077_ _04202_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_143_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12108_ _06193_ cpuregs.regs\[23\]\[12\] _06507_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__mux2_1
X_13088_ _07065_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__clkbuf_1
X_17965_ clknet_leaf_0_clk _01102_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15952__A net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12039_ _06473_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__clkbuf_1
X_16916_ clknet_leaf_15_clk _00097_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17896_ clknet_leaf_95_clk _01065_ VGND VGND VPWR VPWR count_cycle\[41\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15418__C1 _03692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10050__S0 _04057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16847_ _03167_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_158_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15969__B1 _06003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13472__A _04532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16630__A1 _06174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13444__A1 _07304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16778_ _06561_ cpuregs.regs\[13\]\[13\] _03127_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__mux2_1
XANTENNA__10258__A1 _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18517_ clknet_leaf_17_clk _01582_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15729_ _04777_ _02506_ _02534_ _02481_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_66_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10353__S1 _04208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15197__A1 _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09250_ _03959_ _03988_ _03960_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__a21o_1
X_18448_ clknet_leaf_113_clk _01513_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08871__B2 _03636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15292__S1 _01986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09181_ _03891_ _03747_ _03924_ _03930_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__a31o_1
XFILLER_0_173_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18379_ clknet_leaf_118_clk _01444_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08623__A1 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10430__A1 _04054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12027__S _06460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10981__A2 _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12551__A _06751_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16023__A mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08965_ _03205_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__buf_4
XANTENNA__15862__A _03309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15672__A2 _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09887__B1 _04156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08896_ _00064_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__buf_6
XFILLER_0_75_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10497__B2 _04023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12697__S _06836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16621__A1 _06140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09517_ _04245_ _04246_ _04247_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11446__B1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10344__S1 _04759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09448_ cpuregs.regs\[8\]\[3\] cpuregs.regs\[9\]\[3\] cpuregs.regs\[10\]\[3\] cpuregs.regs\[11\]\[3\]
+ _04055_ _04058_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__mux4_1
XANTENNA__16385__A0 _06991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09379_ reg_pc\[1\] decoded_imm\[1\] VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11410_ _06003_ _06017_ cpuregs.raddr1\[2\] _05973_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__15102__A _01959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12390_ cpuregs.waddr\[1\] cpuregs.waddr\[0\] VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__nand2_2
XFILLER_0_62_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11341_ reg_next_pc\[31\] reg_out\[31\] _05928_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__mux2_2
XFILLER_0_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16632__S _03051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14060_ count_instr\[24\] count_instr\[23\] _07805_ VGND VGND VPWR VPWR _07808_ sky130_fd_sc_hd__and3_1
X_11272_ _04754_ _05900_ _05827_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__mux2_1
XANTENNA__14660__B _07968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13011_ cpuregs.regs\[3\]\[13\] _06561_ _07021_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__mux2_1
X_10223_ cpuregs.regs\[16\]\[23\] cpuregs.regs\[17\]\[23\] cpuregs.regs\[18\]\[23\]
+ cpuregs.regs\[19\]\[23\] _04280_ _04059_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__mux4_1
XANTENNA__15112__A1 _05255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10154_ _04483_ _04868_ _04082_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__a21o_1
XANTENNA__11077__A _05323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15663__A2 _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17750_ clknet_leaf_86_clk _00919_ VGND VGND VPWR VPWR count_instr\[21\] sky130_fd_sc_hd__dfxtp_1
X_14962_ _01856_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13674__A1 _04913_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10085_ _04800_ _04801_ _04320_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__mux2_1
XANTENNA__11685__A0 _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16701_ _03089_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__clkbuf_1
X_13913_ _07691_ _07706_ VGND VGND VPWR VPWR _07707_ sky130_fd_sc_hd__and2_1
X_14893_ reg_pc\[31\] _07282_ _05200_ _03387_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__o2bb2a_1
X_17681_ clknet_leaf_142_clk _00850_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13844_ _07661_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16632_ cpuregs.regs\[1\]\[11\] _06183_ _03051_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13775_ _05227_ _05334_ _07216_ VGND VGND VPWR VPWR _07614_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16563_ _03016_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10987_ _03461_ _05301_ _05220_ _03463_ _05669_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__a221o_1
XFILLER_0_168_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16807__S _03138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18302_ clknet_leaf_6_clk _01370_ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15514_ decoded_imm\[24\] _02216_ _02197_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__a21o_1
XANTENNA__15179__A1 _01989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12726_ _06320_ cpuregs.regs\[12\]\[28\] _06847_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16494_ cpuregs.regs\[17\]\[10\] _06554_ _02979_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15445_ net111 _02081_ _02283_ _02284_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15274__S1 _02086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18233_ clknet_leaf_9_clk _01304_ VGND VGND VPWR VPWR cpuregs.raddr1\[1\] sky130_fd_sc_hd__dfxtp_1
X_12657_ _06320_ cpuregs.regs\[30\]\[28\] _06810_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_992 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15012__A _04702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11608_ reg_pc\[10\] _06162_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15376_ cpuregs.regs\[0\]\[17\] cpuregs.regs\[1\]\[17\] cpuregs.regs\[2\]\[17\] cpuregs.regs\[3\]\[17\]
+ _01908_ _01909_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__mux4_1
X_18164_ clknet_leaf_24_clk _01235_ VGND VGND VPWR VPWR decoded_imm_j\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11204__A3 _05840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12588_ _06782_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17115_ clknet_leaf_12_clk _00289_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14327_ compressed_instr _07989_ VGND VGND VPWR VPWR _08003_ sky130_fd_sc_hd__and2_1
XFILLER_0_170_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18095_ clknet_leaf_91_clk _01199_ VGND VGND VPWR VPWR timer\[10\] sky130_fd_sc_hd__dfxtp_1
X_11539_ reg_pc\[3\] reg_pc\[2\] _06090_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10963__A2 _05357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17046_ clknet_leaf_126_clk _00220_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15351__A1 _02020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14258_ _07899_ _07944_ _07946_ _07948_ reg_pc\[18\] VGND VGND VPWR VPWR _00979_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13209_ _06963_ cpuregs.regs\[8\]\[10\] _07129_ VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09664__B decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14189_ _07896_ _07897_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15103__B2 _01932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_350 VGND VGND VPWR VPWR alphacore_350/HI trace_data[11] sky130_fd_sc_hd__conb_1
Xalphacore_361 VGND VGND VPWR VPWR alphacore_361/HI trace_data[22] sky130_fd_sc_hd__conb_1
Xalphacore_372 VGND VGND VPWR VPWR alphacore_372/HI trace_data[33] sky130_fd_sc_hd__conb_1
X_08750_ _03504_ _03508_ _03512_ _03515_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__and4b_1
X_17948_ clknet_leaf_70_clk _08389_ VGND VGND VPWR VPWR reg_out\[28\] sky130_fd_sc_hd__dfxtp_1
X_08681_ net118 net86 VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17879_ clknet_leaf_88_clk _01048_ VGND VGND VPWR VPWR count_cycle\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11140__A2 _05324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13406__S _07225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13417__A1 _04262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09716__S0 _04072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11428__B1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09097__A1 _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09302_ mem_wordsize\[1\] VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_81_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15265__S1 _01986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09233_ _03970_ _03974_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13141__S _07093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09164_ _03916_ _03908_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10403__A1 _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10403__B2 _05087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09095_ _03738_ _03854_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_151_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12156__A1 _06536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15893__A2 _02635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10167__B1 _04673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10706__A2 _05398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09066__S _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10262__S0 _04071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09997_ _04714_ _04715_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__and2_1
X_08948_ cpuregs.regs\[4\]\[4\] cpuregs.regs\[5\]\[4\] cpuregs.regs\[6\]\[4\] cpuregs.regs\[7\]\[4\]
+ _03661_ _03662_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_4_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09590__A _04063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10014__S0 _04280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08879_ cpuregs.regs\[4\]\[2\] cpuregs.regs\[5\]\[2\] cpuregs.regs\[6\]\[2\] cpuregs.regs\[7\]\[2\]
+ _03641_ _03643_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13316__S _07176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10910_ _04708_ _04642_ _05230_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__mux2_1
X_11890_ _06141_ cpuregs.regs\[20\]\[6\] _06387_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__mux2_1
XANTENNA__14605__B1 _08035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16070__A2 _02650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10841_ _03501_ _03505_ _03503_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_158_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16627__S _03040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13560_ _07238_ _07411_ _07413_ _07190_ VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10772_ _03613_ _05467_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12511_ _06741_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13491_ _04419_ _07271_ _07343_ _07349_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15230_ _01905_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_136_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12442_ _06704_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15581__A1 decoded_imm\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13592__A0 _04642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12395__A1 _06536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15161_ cpuregs.regs\[12\]\[6\] cpuregs.regs\[13\]\[6\] cpuregs.regs\[14\]\[6\] cpuregs.regs\[15\]\[6\]
+ _02013_ _02014_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__mux4_1
XANTENNA__16362__S _02907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12373_ _06667_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09260__A1 _03892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11510__D _06083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14112_ _07843_ _07844_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__nor2_1
X_11324_ reg_out\[28\] _05941_ _05942_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15092_ cpuregs.regs\[16\]\[1\] cpuregs.regs\[17\]\[1\] cpuregs.regs\[18\]\[1\] cpuregs.regs\[19\]\[1\]
+ _03669_ _03646_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14043_ count_instr\[17\] _07792_ count_instr\[18\] VGND VGND VPWR VPWR _07797_ sky130_fd_sc_hd__a21o_1
XANTENNA__15884__A2 _02635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11255_ _04642_ _05886_ _05827_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__mux2_1
XANTENNA__13895__A1 _03322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10206_ _04917_ _04918_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__nand2_1
XANTENNA__11519__B _06065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11186_ reg_next_pc\[3\] reg_out\[3\] _03189_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__mux2_1
X_17802_ clknet_leaf_55_clk _00971_ VGND VGND VPWR VPWR reg_pc\[10\] sky130_fd_sc_hd__dfxtp_2
X_10137_ _04391_ _04824_ _04825_ _04852_ VGND VGND VPWR VPWR _08381_ sky130_fd_sc_hd__a31o_1
XANTENNA__13647__A1 _04810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15994_ _03867_ _02707_ _02708_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__a21o_1
XANTENNA__09315__A2 _04008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11658__A0 _06216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17733_ clknet_leaf_93_clk _00902_ VGND VGND VPWR VPWR count_instr\[4\] sky130_fd_sc_hd__dfxtp_1
X_10068_ reg_pc\[18\] decoded_imm\[18\] _04751_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__a21o_1
X_14945_ net207 net176 _01846_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16597__A0 _06999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17664_ clknet_leaf_17_clk _00833_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_14876_ count_cycle\[60\] _01801_ _07675_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10330__B1 instr_rdcycleh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10881__A1 _04602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11254__B _05885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16615_ cpuregs.regs\[1\]\[3\] _06113_ _03040_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__mux2_1
X_13827_ cpuregs.regs\[0\]\[10\] VGND VGND VPWR VPWR _07653_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09079__A1 _03737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08795__A_N net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16537__S _02967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17595_ clknet_leaf_166_clk _00764_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12083__A0 _06078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13758_ net86 decoded_imm\[27\] VGND VGND VPWR VPWR _07598_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16546_ _03007_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08844__A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10633__A1 _05334_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11830__A0 _06184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12709_ _06824_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08921__S1 _03684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13689_ _07304_ _04909_ _07305_ reg_pc\[22\] _07283_ VGND VGND VPWR VPWR _07534_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16477_ cpuregs.regs\[17\]\[2\] _06538_ _02968_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__mux2_1
XANTENNA__15021__B1 _01714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18216_ clknet_leaf_28_clk _01287_ VGND VGND VPWR VPWR instr_srai sky130_fd_sc_hd__dfxtp_2
XFILLER_0_54_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15428_ net109 _02268_ _01905_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18147_ clknet_leaf_46_clk alu_out\[21\] VGND VGND VPWR VPWR alu_out_q\[21\] sky130_fd_sc_hd__dfxtp_1
X_15359_ cpuregs.regs\[28\]\[16\] cpuregs.regs\[29\]\[16\] cpuregs.regs\[30\]\[16\]
+ cpuregs.regs\[31\]\[16\] _01990_ _01992_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__mux4_1
XFILLER_0_171_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16272__S _02859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09251__A1 _03737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18078_ clknet_leaf_73_clk _01183_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09920_ _04639_ _04640_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__xnor2_1
X_17029_ clknet_leaf_156_clk _00203_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12305__S _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09851_ cpuregs.regs\[16\]\[13\] cpuregs.regs\[17\]\[13\] cpuregs.regs\[18\]\[13\]
+ cpuregs.regs\[19\]\[13\] _04512_ _04513_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_111_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _03488_ _03565_ _03567_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__o21a_1
XANTENNA__11361__A2 _03874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09782_ _04420_ _04506_ _03225_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08733_ _03497_ _03498_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_147_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13136__S _07082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09711__C1 _04296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08664_ instr_bgeu instr_bge instr_bne VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__or3_1
XANTENNA__12040__S _06471_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08457__C net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16052__A2 decoded_imm_j\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15486__S1 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08595_ _03309_ cpu_state\[3\] _03310_ _01226_ _03373_ VGND VGND VPWR VPWR _03374_
+ sky130_fd_sc_hd__a311o_1
XANTENNA__16447__S _02954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08754__A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15238__S1 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11821__A0 _06150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_986 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08473__B instr_lui VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09216_ _03762_ _03892_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09288__C instr_retirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15563__B2 _02004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09147_ _03854_ _03902_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_954 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10483__S0 _04274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09078_ _03839_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_32_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12215__S _06576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11040_ _05485_ _05621_ _05717_ _05597_ _05718_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__a221o_1
XANTENNA__11888__A0 _06132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10243__B decoded_imm\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13629__A1 _04913_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15174__S0 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16211__A net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _07014_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11104__A2 _05398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_1015 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13046__S _07009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12301__A1 _06580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11355__A _03199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14730_ count_cycle\[13\] count_cycle\[14\] _08359_ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__and3_1
X_11942_ _06343_ cpuregs.regs\[20\]\[31\] _06386_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16043__A2 _02711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14661_ _08221_ _07968_ VGND VGND VPWR VPWR _08310_ sky130_fd_sc_hd__or2_1
X_11873_ cpuregs.waddr\[1\] cpuregs.waddr\[0\] VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__nor2_4
XANTENNA__12885__S _06943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _07445_ _07450_ _07461_ _03311_ VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16400_ _02929_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10824_ instr_sub VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__buf_4
X_17380_ clknet_leaf_16_clk _00549_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_14592_ _07958_ _08236_ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__or2_1
XANTENNA__13801__A1 _05143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13543_ net70 decoded_imm\[12\] VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16331_ _02892_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10755_ _05450_ _05451_ _05390_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12186__A _06183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10091__A2 _04806_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16262_ _02855_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__clkbuf_1
X_13474_ _07279_ _07273_ _07331_ _07333_ VGND VGND VPWR VPWR _07334_ sky130_fd_sc_hd__a31o_1
X_10686_ _05369_ _05378_ _05386_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__or3_1
XFILLER_0_125_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12368__A1 _06578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output197_A net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18001_ clknet_leaf_66_clk _01138_ VGND VGND VPWR VPWR irq_mask\[17\] sky130_fd_sc_hd__dfxtp_1
X_15213_ _02061_ _02062_ _02063_ _02064_ _01982_ _02004_ VGND VGND VPWR VPWR _02065_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09769__C1 _04188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12425_ _06695_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__clkbuf_1
X_16193_ _02814_ _02815_ _02816_ _02676_ net296 VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__a32o_1
XFILLER_0_124_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12914__A _06174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10918__A2 _05220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15306__A1 _01982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15144_ _01995_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__buf_8
XANTENNA__09495__A net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12356_ _06658_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11307_ reg_next_pc\[25\] reg_out\[25\] _05928_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__mux2_2
XFILLER_0_121_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15401__S1 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15075_ is_slli_srli_srai cpuregs.raddr2\[0\] decoded_imm\[0\] _01933_ _01934_ VGND
+ VGND VPWR VPWR _01935_ sky130_fd_sc_hd__a221o_1
X_12287_ _06621_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12125__S _06518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output74_A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14026_ count_instr\[12\] _07781_ count_instr\[13\] VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__a21o_1
XANTENNA__11249__B _05881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09536__A2 _04262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11238_ _05862_ _05864_ _05868_ _05871_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_56_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15944__B mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11169_ net117 _04710_ _05819_ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__a21o_2
XFILLER_0_93_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15977_ _02694_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17716_ clknet_leaf_76_clk _00885_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dfxtp_1
X_14928_ net199 net168 _01835_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__mux2_1
XANTENNA__09395__S1 _04073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16034__A2 decoded_imm_j\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10854__A1 _05414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17647_ clknet_leaf_47_clk _00816_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfxtp_4
XANTENNA__12795__S _06891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14859_ _01792_ _01793_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15242__B1 _03654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13480__A _04566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15171__S _01984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17578_ clknet_leaf_182_clk _00747_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14295__B _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16529_ cpuregs.regs\[17\]\[27\] _06590_ _02990_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14348__A2 _07948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10328__B _05037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12359__A1 _06569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09001_ _03762_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_171_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09224__A1 _03965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11567__C1 _06118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09775__A2 _04049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15848__A2 _03810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09903_ _04070_ _04624_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15854__B _02613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09834_ _04556_ _04557_ _04077_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16031__A instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09344__S _04078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09765_ _04053_ _04490_ _04095_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__a21o_1
XANTENNA__14284__A1 reg_next_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08468__B instr_maskirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15481__B1 _03674_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08716_ _03480_ _03481_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__and2_1
X_09696_ net49 _04030_ _04034_ net63 _04423_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__o221a_1
X_08647_ _03414_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14486__A decoded_imm_j\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08578_ irq_mask\[12\] irq_pending\[12\] VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__and2b_2
XANTENNA__14587__A2 _07956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10540_ _03531_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__buf_4
XFILLER_0_148_1019 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16733__A0 _06999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13547__B1 _03631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10471_ irq_pending\[30\] _04007_ _05173_ _05176_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__o22a_1
XFILLER_0_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12734__A _03298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16206__A net299 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12210_ _06247_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__buf_2
XANTENNA__11022__A1 _04945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13190_ _06945_ cpuregs.regs\[8\]\[1\] _07118_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__mux2_1
XANTENNA__10456__S0 _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12141_ _06320_ cpuregs.regs\[23\]\[28\] _06518_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16640__S _03051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12072_ _06490_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11784__S _06258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13565__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11023_ _05702_ _05682_ _05658_ _05633_ _05266_ _05395_ VGND VGND VPWR VPWR _05703_
+ sky130_fd_sc_hd__mux4_1
X_15900_ _03940_ _02613_ _02612_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__and3b_1
XANTENNA__15256__S _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16880_ _03184_ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__clkbuf_1
X_15831_ decoded_imm_j\[17\] _05983_ _02596_ _02597_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_144_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ clknet_leaf_189_clk _01615_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15762_ _05069_ _02479_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__nand2_1
X_12974_ _07003_ cpuregs.regs\[31\]\[29\] _06985_ VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__mux2_1
X_17501_ clknet_leaf_119_clk _00670_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10297__C1 _04296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14713_ count_cycle\[7\] _08346_ count_cycle\[8\] VGND VGND VPWR VPWR _08351_ sky130_fd_sc_hd__a21o_1
X_18481_ clknet_leaf_116_clk _01546_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_11925_ _06412_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output112_A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15693_ timer\[9\] timer\[8\] _02500_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__or3_2
XFILLER_0_87_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13504__S _07225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12038__A0 _06184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17432_ clknet_leaf_165_clk _00601_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15775__A1 _05170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11856_ _06374_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__clkbuf_1
X_14644_ reg_next_pc\[27\] _07948_ _08286_ _08294_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10807_ _03511_ _03514_ _03513_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17363_ clknet_leaf_98_clk _00532_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_14575_ _08212_ _07956_ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11787_ reg_pc\[30\] _06322_ _06101_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16314_ _06989_ cpuregs.regs\[15\]\[22\] _02881_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13526_ _04642_ _07276_ VGND VGND VPWR VPWR _07382_ sky130_fd_sc_hd__or2_1
X_10738_ _05277_ _05333_ _05435_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08662__C1 _03305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17294_ clknet_leaf_98_clk _00468_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15939__B mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11959__S _06424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13457_ _04262_ _05257_ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__or2_1
XANTENNA__15622__S1 _03647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16245_ net57 mem_16bit_buffer\[15\] _02830_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__mux2_1
X_10669_ _04532_ _04566_ _04602_ _04611_ _05230_ _05240_ VGND VGND VPWR VPWR _05370_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_113_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11549__C1 _06118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08841__B net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12408_ _06686_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11013__B2 _05281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10447__S0 _04472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13388_ _03399_ _07252_ VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16176_ _02806_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__clkbuf_1
Xoutput106 net106 VGND VGND VPWR VPWR cpi_rs2[16] sky130_fd_sc_hd__buf_1
XFILLER_0_23_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput117 net117 VGND VGND VPWR VPWR cpi_rs2[26] sky130_fd_sc_hd__clkbuf_1
Xoutput128 net128 VGND VGND VPWR VPWR cpi_rs2[7] sky130_fd_sc_hd__clkbuf_1
X_15127_ _01907_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__buf_8
XFILLER_0_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12339_ _06649_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__clkbuf_1
Xoutput139 net139 VGND VGND VPWR VPWR eoi[17] sky130_fd_sc_hd__buf_1
XFILLER_0_11_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15386__S0 _01908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15058_ _03670_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__buf_8
XANTENNA__11694__S _06176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14009_ count_instr\[8\] count_instr\[7\] count_instr\[6\] _07767_ VGND VGND VPWR
+ VPWR _07773_ sky130_fd_sc_hd__and4_2
XANTENNA__13475__A _03387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15138__S0 _01990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09550_ _04280_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__buf_6
X_08501_ instr_lw _03283_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__or2_1
XANTENNA__10827__A1 _05517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09481_ _04206_ _04212_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12029__A0 _06150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08432_ mem_do_rdata VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08879__S0 _03641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16725__S _03098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11252__A1 _05829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13529__B1 _07211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15613__S1 _01937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10773__S _05363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16026__A mem_rdata_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15865__A _02612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10763__A0 _03518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13385__A _04142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10802__A _05218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09817_ _04461_ _04501_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_126_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15454__B1 _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10530__A3 _04642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09748_ cpuregs.regs\[28\]\[10\] cpuregs.regs\[29\]\[10\] cpuregs.regs\[30\]\[10\]
+ cpuregs.regs\[31\]\[10\] _04472_ _04473_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__mux4_1
XANTENNA__09133__A0 mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09679_ cpuregs.regs\[24\]\[8\] cpuregs.regs\[25\]\[8\] cpuregs.regs\[26\]\[8\] cpuregs.regs\[27\]\[8\]
+ _04085_ _04087_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09684__A1 _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15206__B1 _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11710_ reg_out\[21\] alu_out_q\[21\] _06069_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12690_ _06837_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11641_ _06201_ cpuregs.regs\[10\]\[13\] _06176_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10765__A2_N _05221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14360_ reg_next_pc\[4\] _07947_ _08032_ _08033_ VGND VGND VPWR VPWR _08034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11572_ _06136_ _06139_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__nor2_2
XFILLER_0_25_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13311_ _07183_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__clkbuf_1
Xinput19 irq[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlymetal6s2s_1
X_10523_ _05209_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__buf_4
XANTENNA__15604__S1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14291_ reg_pc\[30\] _07953_ _07969_ _07960_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13242_ _06997_ cpuregs.regs\[8\]\[26\] _07140_ VGND VGND VPWR VPWR _07147_ sky130_fd_sc_hd__mux2_1
X_16030_ _02725_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__buf_2
X_10454_ _04231_ _05159_ _04082_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15390__C1 _02197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13173_ _07110_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15368__S0 _01985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16370__S _02907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10385_ _04328_ _05092_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_36_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12124_ _06495_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_36_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17981_ clknet_leaf_43_clk _01118_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_53_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14496__A1 reg_next_pc\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14496__B2 _08033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16932_ clknet_leaf_153_clk _00113_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_12055_ _06481_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12403__S _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11006_ _05281_ _05684_ _05687_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__a21o_1
XANTENNA__09372__B1 _04009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09911__A2 _04021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16863_ _06578_ cpuregs.regs\[14\]\[21\] _03174_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__mux2_1
XANTENNA__14248__A1 reg_next_pc\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15445__B1 _02283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08724__B_N net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18602_ clknet_leaf_151_clk _01667_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_15814_ decoded_imm_j\[7\] _05983_ _03977_ _02587_ _02590_ VGND VGND VPWR VPWR _01237_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15540__S0 _03645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16794_ _03139_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__clkbuf_1
X_18533_ clknet_leaf_135_clk _01598_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15745_ timer\[22\] _02540_ timer\[23\] VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12957_ _06992_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11543__A _06113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13234__S _07140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11482__A1 _06054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15748__A1 _04941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11908_ _06403_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__clkbuf_1
X_18464_ clknet_leaf_158_clk _01529_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_15676_ timer\[5\] _02493_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__or2_1
X_12888_ _06945_ cpuregs.regs\[31\]\[1\] _06943_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17415_ clknet_leaf_178_clk _00584_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14627_ _08050_ _08278_ VGND VGND VPWR VPWR _08279_ sky130_fd_sc_hd__or2_1
XANTENNA__09427__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18395_ clknet_leaf_181_clk _01460_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11839_ _06365_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16545__S _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10037__A2 _04754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17346_ clknet_leaf_187_clk _00515_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14558_ _08214_ _08215_ VGND VGND VPWR VPWR _08216_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08852__A net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13509_ _07363_ _07355_ _07364_ _03311_ VGND VGND VPWR VPWR _07366_ sky130_fd_sc_hd__a31o_1
XFILLER_0_130_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17277_ clknet_leaf_2_clk _00451_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16173__A1 net242 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14489_ _08131_ _08151_ VGND VGND VPWR VPWR _08152_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16228_ _02838_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15685__A _04382_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15359__S0 _01990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16280__S _02859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16159_ net272 net234 _02797_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08981_ mem_16bit_buffer\[14\] _03742_ _03205_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__mux2_4
XFILLER_0_54_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09589__S1 _04317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12313__S _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10622__A _05323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11170__B1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10341__B decoded_imm\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09602_ _04330_ _04331_ _04222_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__mux2_1
XANTENNA__15987__A1 _03767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15987__B2 _03880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09533_ _04036_ mem_wordsize\[1\] _04263_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13652__B decoded_imm\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13998__B1 _07759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09464_ _04195_ _04196_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_121_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08415_ net33 mem_rdata_q\[0\] _03200_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09395_ cpuregs.regs\[28\]\[2\] cpuregs.regs\[29\]\[2\] cpuregs.regs\[30\]\[2\] cpuregs.regs\[31\]\[2\]
+ _04071_ _04073_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__mux4_1
XFILLER_0_163_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16455__S _02954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10028__A2 _04744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08762__A net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10433__C1 _04188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10984__A0 _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15598__S0 _01908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08929__B1 _03692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10008__S _04078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10200__A2 _04745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10170_ reg_pc\[22\] decoded_imm\[22\] VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__nand2_1
XANTENNA__13686__C1 _07217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15427__B1 _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13860_ _07669_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_141_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09532__S _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12811_ cpuregs.regs\[9\]\[31\] _06598_ _06868_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__mux2_1
XANTENNA__13989__B1 _07759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10678__S _05239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13791_ _07238_ _07627_ _07628_ _07190_ VGND VGND VPWR VPWR _07629_ sky130_fd_sc_hd__a211o_1
XANTENNA__09657__A1 instr_rdcycleh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12459__A _06081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14650__A1 _07966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13054__S _07046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11363__A _03979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15530_ decoded_imm\[25\] _02216_ _02197_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__a21o_1
XANTENNA__12661__A0 _06336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12742_ cpuregs.waddr\[1\] _06862_ _06866_ _06861_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15461_ net112 _02081_ _02298_ _02299_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__o22a_1
X_12673_ _06828_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_13_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_190_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_190_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14674__A _07968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17200_ clknet_leaf_110_clk _00374_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11624_ _06071_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__buf_4
X_14412_ _03294_ _07925_ _07997_ _08080_ VGND VGND VPWR VPWR _08081_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09768__A _04051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18180_ clknet_leaf_32_clk _01251_ VGND VGND VPWR VPWR instr_lui sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_139_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ cpuregs.regs\[20\]\[18\] cpuregs.regs\[21\]\[18\] cpuregs.regs\[22\]\[18\]
+ cpuregs.regs\[23\]\[18\] _01995_ _01937_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17131_ clknet_leaf_149_clk _00305_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11555_ _06124_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__buf_2
X_14343_ decoded_imm_j\[3\] _07911_ VGND VGND VPWR VPWR _08018_ sky130_fd_sc_hd__nor2_1
XANTENNA__15589__S0 _02221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10506_ instr_sll instr_slli VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__nor2_2
X_14274_ _05909_ _06286_ _07942_ _05922_ VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__o211a_2
X_17062_ clknet_leaf_139_clk _00236_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11486_ _06054_ irq_pending\[30\] _06062_ net24 VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13225_ _06980_ cpuregs.regs\[8\]\[18\] _07129_ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__mux2_1
X_16013_ decoded_imm\[0\] _02711_ _02713_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__o21a_1
X_10437_ net54 _04811_ _04667_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09593__B1 _04225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13156_ _07101_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13737__B decoded_imm\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10368_ net52 _04811_ _04666_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__a21o_1
XANTENNA__14469__A1 _07998_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12107_ _06509_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__clkbuf_1
X_13087_ _06978_ cpuregs.regs\[7\]\[17\] _07057_ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__mux2_1
X_17964_ clknet_leaf_191_clk _01101_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dfxtp_1
XANTENNA__12133__S _06518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10299_ irq_mask\[25\] _04448_ timer\[25\] _04187_ _04188_ VGND VGND VPWR VPWR _05010_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16915_ clknet_leaf_190_clk _00096_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12038_ _06184_ cpuregs.regs\[22\]\[11\] _06471_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__mux2_1
XANTENNA__11152__A0 _05277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11257__B _05885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15952__B net299 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10161__B decoded_imm\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17895_ clknet_leaf_96_clk _01064_ VGND VGND VPWR VPWR count_cycle\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09440__S0 _04071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11972__S _06435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13753__A _05205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10050__S1 _04060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16846_ _06561_ cpuregs.regs\[14\]\[13\] _03163_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__mux2_1
XANTENNA__15969__A1 _04168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08847__A net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09442__S _04077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16777_ _03130_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13444__A2 _04307_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13989_ count_instr\[1\] _07756_ _07759_ VGND VGND VPWR VPWR _07760_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18516_ clknet_leaf_174_clk _01581_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_15728_ _02476_ _02532_ _02533_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__or3b_1
XFILLER_0_125_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18447_ clknet_leaf_165_clk _01512_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15659_ timer\[1\] VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_181_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_181_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09180_ _03895_ _03927_ _03928_ _03929_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18378_ clknet_leaf_98_clk _01443_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13601__C1 _07217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17329_ clknet_leaf_161_clk _00503_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16146__A1 net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09820__B2 _04013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15619__S _03653_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_1010 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10194__A1 _04296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_951 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11448__A _03412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08964_ _03400_ _03706_ _03726_ _03638_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__o22a_1
XANTENNA__15862__B _03304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15409__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08895_ cpuregs.regs\[20\]\[2\] cpuregs.regs\[21\]\[2\] cpuregs.regs\[22\]\[2\] cpuregs.regs\[23\]\[2\]
+ _03658_ _03659_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__mux4_1
XANTENNA__11143__B1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11882__S _06387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10497__A2 _04021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12891__A0 _06947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08757__A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16082__B1 _06016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14632__A1 reg_next_pc\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14632__B2 _08033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10249__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09516_ _04245_ _04246_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12643__A0 _06266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09447_ cpuregs.regs\[12\]\[3\] cpuregs.regs\[13\]\[3\] cpuregs.regs\[14\]\[3\] cpuregs.regs\[15\]\[3\]
+ _04055_ _04058_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__mux4_1
XFILLER_0_164_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16185__S _02770_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_172_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_172_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_148_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16334__A_N cpuregs.waddr\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09378_ reg_pc\[1\] decoded_imm\[1\] VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__nand2_1
XANTENNA__08492__A _03274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10527__A net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12218__S _06576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11340_ _05956_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__buf_2
XFILLER_0_22_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11271_ _05896_ _05899_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13010_ _07024_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10222_ cpuregs.regs\[20\]\[23\] cpuregs.regs\[21\]\[23\] cpuregs.regs\[22\]\[23\]
+ cpuregs.regs\[23\]\[23\] _04280_ _04059_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__mux4_1
XANTENNA__09670__S0 _04072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10153_ _04866_ _04867_ _04575_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__mux2_1
XANTENNA__15112__A2 _01906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14961_ net216 net185 _01846_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__mux2_1
X_10084_ cpuregs.regs\[8\]\[19\] cpuregs.regs\[9\]\[19\] cpuregs.regs\[10\]\[19\]
+ cpuregs.regs\[11\]\[19\] _04273_ _04283_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__mux4_1
XANTENNA__12888__S _06943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14669__A _08232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16700_ _06966_ cpuregs.regs\[19\]\[11\] _03087_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__mux2_1
X_13912_ _03333_ _07704_ _07705_ net132 VGND VGND VPWR VPWR _07706_ sky130_fd_sc_hd__a22o_1
X_17680_ clknet_leaf_134_clk _00849_ VGND VGND VPWR VPWR cpuregs.regs\[0\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08667__A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14892_ _05174_ _07279_ _07274_ _05076_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_18_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16631_ _03052_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__clkbuf_1
X_13843_ cpuregs.regs\[0\]\[18\] VGND VGND VPWR VPWR _07661_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12189__A _06192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16562_ _06963_ cpuregs.regs\[18\]\[10\] _03015_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__mux2_1
X_10986_ _03462_ _05398_ _05646_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__o21ai_1
X_13774_ _05143_ _05076_ _05227_ VGND VGND VPWR VPWR _07613_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18301_ clknet_leaf_5_clk _01369_ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15513_ _02336_ _02340_ _02027_ _02348_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__o211a_2
X_12725_ _06855_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16493_ _02967_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_163_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_163_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_167_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18232_ clknet_leaf_9_clk _01303_ VGND VGND VPWR VPWR cpuregs.raddr1\[0\] sky130_fd_sc_hd__dfxtp_1
X_15444_ decoded_imm\[20\] _02216_ _02197_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12656_ _06818_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09489__S0 _04217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15012__B _01885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18163_ clknet_leaf_23_clk _01234_ VGND VGND VPWR VPWR decoded_imm_j\[4\] sky130_fd_sc_hd__dfxtp_1
X_11607_ reg_pc\[10\] _06162_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__and2_1
X_15375_ cpuregs.regs\[4\]\[17\] cpuregs.regs\[5\]\[17\] cpuregs.regs\[6\]\[17\] cpuregs.regs\[7\]\[17\]
+ _01908_ _01909_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__mux4_1
X_12587_ cpuregs.regs\[2\]\[27\] _06590_ _06774_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__mux2_1
XANTENNA__16823__S _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09802__B2 instr_timer VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17114_ clknet_leaf_187_clk _00288_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14326_ _07909_ _07997_ VGND VGND VPWR VPWR _08002_ sky130_fd_sc_hd__or2_1
X_18094_ clknet_leaf_103_clk _01198_ VGND VGND VPWR VPWR timer\[9\] sky130_fd_sc_hd__dfxtp_1
X_11538_ irq_state\[0\] reg_next_pc\[3\] _03344_ _06072_ _06101_ VGND VGND VPWR VPWR
+ _06109_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17045_ clknet_leaf_116_clk _00219_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11469_ _03277_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__clkbuf_8
X_14257_ _07947_ VGND VGND VPWR VPWR _07948_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09566__B1 _04296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13208_ _07117_ VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__clkbuf_8
X_14188_ count_instr\[63\] count_instr\[62\] _07893_ _03240_ VGND VGND VPWR VPWR _07897_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10176__B2 _04013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13139_ _07092_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xalphacore_340 VGND VGND VPWR VPWR alphacore_340/HI trace_data[1] sky130_fd_sc_hd__conb_1
Xalphacore_351 VGND VGND VPWR VPWR alphacore_351/HI trace_data[12] sky130_fd_sc_hd__conb_1
Xalphacore_362 VGND VGND VPWR VPWR alphacore_362/HI trace_data[23] sky130_fd_sc_hd__conb_1
Xalphacore_373 VGND VGND VPWR VPWR alphacore_373/HI trace_data[34] sky130_fd_sc_hd__conb_1
X_17947_ clknet_leaf_74_clk _08388_ VGND VGND VPWR VPWR reg_out\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09869__A1 _04296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08680_ _03439_ _03442_ _03445_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__or3b_1
X_17878_ clknet_leaf_85_clk _01047_ VGND VGND VPWR VPWR count_cycle\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09172__S _03757_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16829_ _06544_ cpuregs.regs\[14\]\[5\] _03152_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09716__S1 _04074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09301_ _04036_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_165_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_154_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_154_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09232_ _03895_ _03971_ _03972_ _03822_ _03973_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09163_ _03818_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12038__S _06471_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10347__A _04272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16733__S _03098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10403__A2 _05086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09094_ _03750_ _03844_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__or2_2
XFILLER_0_32_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10066__B decoded_imm\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15349__S _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10167__B2 _04881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10262__S1 _04073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09996_ reg_pc\[17\] decoded_imm\[17\] VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_134_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11116__A0 _05174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08947_ _03707_ _03708_ _03709_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__mux2_1
XANTENNA__09404__S0 _04123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10014__S1 _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12501__S _06726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08878_ _03642_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14605__A1 _07754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10840_ _03503_ _03506_ _05501_ _03501_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09088__A2 _03737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10771_ _03519_ _05428_ _05429_ _05466_ _03520_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__o311a_1
XFILLER_0_165_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_145_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_145_clk sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_143_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_554 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12737__A _03364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_142_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15113__A _03654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12510_ _06281_ cpuregs.regs\[28\]\[23\] _06737_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__mux2_1
X_13490_ _07347_ _07348_ _07271_ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15030__A1 _03303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12441_ cpuregs.regs\[27\]\[23\] _06582_ _06700_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15581__A2 _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15318__C1 _01969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15160_ _03643_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12372_ cpuregs.regs\[26\]\[23\] _06582_ _06663_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_157_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11323_ reg_next_pc\[28\] _05928_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__or2_1
X_14111_ count_instr\[39\] _07840_ _07834_ VGND VGND VPWR VPWR _07844_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10691__S _05390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15091_ cpuregs.regs\[20\]\[1\] cpuregs.regs\[21\]\[1\] cpuregs.regs\[22\]\[1\] cpuregs.regs\[23\]\[1\]
+ _03669_ _03646_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__mux4_1
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14042_ count_instr\[15\] _07787_ _07795_ VGND VGND VPWR VPWR _07796_ sky130_fd_sc_hd__and3_1
X_11254_ _05882_ _05885_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10158__A1 _04168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_152_Left_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10205_ reg_pc\[23\] decoded_imm\[23\] VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11185_ _03219_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17801_ clknet_leaf_55_clk _00970_ VGND VGND VPWR VPWR reg_pc\[9\] sky130_fd_sc_hd__dfxtp_1
X_10136_ _03303_ _04844_ _04847_ _04851_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__a31o_1
X_15993_ decoded_rd\[1\] _05987_ _03880_ _05977_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__a22o_1
XANTENNA__13647__A2 _05260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17732_ clknet_leaf_101_clk _00901_ VGND VGND VPWR VPWR count_instr\[3\] sky130_fd_sc_hd__dfxtp_1
X_10067_ _04782_ _04783_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__nand2_1
X_14944_ _01847_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12411__S _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17663_ clknet_leaf_70_clk _00832_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfxtp_4
X_14875_ count_cycle\[60\] _01801_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__and2_1
X_16614_ _03043_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__clkbuf_1
X_13826_ _07652_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__clkbuf_1
X_17594_ clknet_leaf_111_clk _00763_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_161_Left_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14846__B _01753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16545_ _06947_ cpuregs.regs\[18\]\[2\] _03004_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13757_ _07191_ _07592_ _07594_ _07596_ VGND VGND VPWR VPWR _07597_ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_136_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_136_clk sky130_fd_sc_hd__clkbuf_2
X_10969_ _03572_ _05652_ _05363_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13242__S _07140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11551__A reg_pc\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12708_ _06846_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16476_ _02970_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__clkbuf_1
X_13688_ _04945_ _07277_ _07532_ _07238_ VGND VGND VPWR VPWR _07533_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18215_ clknet_leaf_39_clk _01286_ VGND VGND VPWR VPWR instr_and sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09021__A _03206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15958__A mem_do_wdata VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15427_ _01959_ _02259_ _02267_ _01933_ decoded_imm\[19\] VGND VGND VPWR VPWR _02268_
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_170_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12639_ _06809_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16553__S _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18146_ clknet_leaf_70_clk alu_out\[20\] VGND VGND VPWR VPWR alu_out_q\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14780__B1 _03240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15358_ _01982_ _02199_ _02201_ _02006_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__o211a_1
XANTENNA__10397__A1 _04214_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14309_ _07985_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__clkbuf_4
X_18077_ clknet_leaf_73_clk _01182_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_41_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16521__A1 _06582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15289_ cpuregs.regs\[12\]\[12\] cpuregs.regs\[13\]\[12\] cpuregs.regs\[14\]\[12\]
+ cpuregs.regs\[15\]\[12\] _01976_ _01977_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_170_Left_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12813__C _06083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17028_ clknet_leaf_157_clk _00202_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09850_ cpuregs.regs\[20\]\[13\] cpuregs.regs\[21\]\[13\] cpuregs.regs\[22\]\[13\]
+ cpuregs.regs\[23\]\[13\] _04512_ _04513_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_111_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ net107 _03566_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__or2_1
XANTENNA__09691__A _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09781_ net52 _04030_ _04034_ net35 _04423_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__o221a_1
XANTENNA__13638__A2 _04806_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08732_ net102 net70 VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__nand2_1
X_08663_ timer\[0\] _03427_ _03429_ net1 VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__a211o_1
X_08594_ _03196_ _03316_ _03318_ _03372_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__or4_1
XFILLER_0_163_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_127_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_127_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08754__B net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09215_ _03843_ _03902_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__or2b_1
XFILLER_0_161_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16463__S _02954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09146_ _03868_ _03866_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__or2_2
XFILLER_0_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09077_ _03786_ _03838_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_131_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08450__B1 _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10483__S1 _04317_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14523__B1 _07997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10524__B _05227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13877__A2 _07679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_168_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09979_ _04697_ _04698_ _04320_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__mux2_1
XANTENNA__15174__S1 _02014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16211__B net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13327__S _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14012__A _03239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12990_ cpuregs.regs\[3\]\[3\] _06540_ _07010_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11941_ _06420_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16638__S _03051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15542__S _03709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14660_ _08232_ _07968_ VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__nand2_1
XANTENNA__15787__C1 _03226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11872_ _06382_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_28_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _07459_ _07460_ VGND VGND VPWR VPWR _07461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10823_ _05219_ _05505_ _05516_ VGND VGND VPWR VPWR alu_out\[10\] sky130_fd_sc_hd__o21ai_2
XFILLER_0_138_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13262__A0 _06949_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_118_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_118_clk sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14591_ _07958_ _08236_ VGND VGND VPWR VPWR _08246_ sky130_fd_sc_hd__nand2_1
XANTENNA__13062__S _07046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16330_ _07005_ cpuregs.regs\[15\]\[30\] _02858_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__mux2_1
X_13542_ net69 decoded_imm\[11\] _07393_ _07395_ _07396_ VGND VGND VPWR VPWR _07397_
+ sky130_fd_sc_hd__a221oi_2
XANTENNA__15539__C1 _01968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10754_ _03519_ _05430_ _03520_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16261_ _07737_ _03216_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10685_ _05254_ _05260_ _05385_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__and3_1
X_13473_ _07217_ _07278_ _07332_ _07189_ VGND VGND VPWR VPWR _07333_ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18000_ clknet_leaf_79_clk _01137_ VGND VGND VPWR VPWR irq_mask\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15212_ cpuregs.regs\[0\]\[8\] cpuregs.regs\[1\]\[8\] cpuregs.regs\[2\]\[8\] cpuregs.regs\[3\]\[8\]
+ _01979_ _01980_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__mux4_1
X_12424_ cpuregs.regs\[27\]\[15\] _06565_ _06689_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__mux2_1
X_16192_ net257 net259 _01822_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10379__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09864__S0 _04280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15143_ cpuregs.regs\[12\]\[5\] cpuregs.regs\[13\]\[5\] cpuregs.regs\[14\]\[5\] cpuregs.regs\[15\]\[5\]
+ _01996_ _01997_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__mux4_1
X_12355_ cpuregs.regs\[26\]\[15\] _06565_ _06652_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__mux2_1
XANTENNA__10715__A _05292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11306_ _05898_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__buf_2
XFILLER_0_132_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15074_ _03277_ _03301_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__nand2_4
X_12286_ cpuregs.regs\[25\]\[15\] _06565_ _06615_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__mux2_1
X_14025_ count_instr\[13\] count_instr\[12\] _07781_ VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__and3_1
X_11237_ _05862_ _05864_ _05868_ _05871_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__and4_1
XANTENNA__12930__A _06215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15944__C mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09941__B1 _04017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output67_A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11168_ _04038_ _05277_ net100 _03297_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__a22o_1
X_10119_ cpuregs.regs\[28\]\[20\] cpuregs.regs\[29\]\[20\] cpuregs.regs\[30\]\[20\]
+ cpuregs.regs\[31\]\[20\] _04275_ _04278_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__mux4_1
XANTENNA__12141__S _06518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11099_ _03445_ _05773_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10450__A _04483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15976_ instr_waitirq _02693_ _03635_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__mux2_1
X_17715_ clknet_leaf_76_clk _00884_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11265__B _05894_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14927_ _01838_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10303__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11980__S _06435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17646_ clknet_leaf_47_clk _00815_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfxtp_4
XANTENNA__10854__A2 _05404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14858_ count_cycle\[54\] _01789_ _01723_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15242__A1 _01989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13809_ cpuregs.regs\[0\]\[1\] VGND VGND VPWR VPWR _07644_ sky130_fd_sc_hd__clkbuf_1
X_17577_ clknet_leaf_183_clk _00746_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_109_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_109_clk sky130_fd_sc_hd__clkbuf_2
X_14789_ count_cycle\[31\] _01741_ count_cycle\[32\] VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__a21o_1
XANTENNA__08574__B irq_pending\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16528_ _02997_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09472__A2 _04104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16459_ _06997_ cpuregs.regs\[29\]\[26\] _02954_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__mux2_1
XANTENNA__14592__A _07958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09000_ mem_16bit_buffer\[11\] _03761_ _03727_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__mux2_4
XFILLER_0_170_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09686__A _04099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11567__B1 _06098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09855__S0 _04512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18129_ clknet_leaf_26_clk alu_out\[3\] VGND VGND VPWR VPWR alu_out_q\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08983__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15848__A3 _03864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09902_ _04622_ _04623_ _04078_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15854__C _03940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09833_ cpuregs.regs\[16\]\[12\] cpuregs.regs\[17\]\[12\] cpuregs.regs\[18\]\[12\]
+ cpuregs.regs\[19\]\[12\] _04071_ _04073_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13147__S _07093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09764_ _04488_ _04489_ _04320_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__mux2_1
XANTENNA__15481__A1 _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08468__C instr_retirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08715_ net108 net76 VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__nand2_1
XANTENNA__15870__B _02613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12986__S _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09695_ _04421_ latched_is_lh _04422_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__o21a_2
XANTENNA__11890__S _06387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08646_ net23 _03394_ _03413_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__or3_1
XFILLER_0_96_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16430__A0 _06968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13244__A0 _06999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08577_ irq_mask\[15\] irq_pending\[15\] VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__and2b_2
XANTENNA__10058__B1 _04133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15092__S0 _03669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10470_ _04046_ _05174_ _04752_ _05175_ _04266_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12734__B _03277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14192__B_N irq_state\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09129_ _03878_ _03880_ _03881_ _03886_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10456__S1 _04478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12140_ _06526_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08785__A_N net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12071_ _06312_ cpuregs.regs\[22\]\[27\] _06482_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11022_ _04959_ _04945_ _05230_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__mux2_1
XANTENNA__13565__B decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11366__A _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15830_ _05987_ _06017_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__nor2_1
X_15761_ _03417_ _02547_ _02554_ _02557_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__o22ai_1
XANTENNA__12286__A1 _06565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16368__S _02907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12973_ _06327_ VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__buf_2
XANTENNA__09151__A1 _03781_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17500_ clknet_leaf_105_clk _00669_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13581__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14712_ _03304_ VGND VGND VPWR VPWR _08350_ sky130_fd_sc_hd__clkbuf_4
X_11924_ _06274_ cpuregs.regs\[20\]\[22\] _06409_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18480_ clknet_leaf_108_clk _01545_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15692_ timer\[8\] _02503_ timer\[9\] VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08675__A net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17431_ clknet_leaf_118_clk _00600_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14643_ _08012_ _08292_ _08293_ VGND VGND VPWR VPWR _08294_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_169_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11855_ _06281_ cpuregs.regs\[11\]\[23\] _06370_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output105_A net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15775__A2 _02486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10049__B1 _04082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10806_ _03512_ _03515_ _03613_ _05467_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__or4_1
XANTENNA__13330__S0 _04207_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17362_ clknet_leaf_99_clk _00531_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14574_ reg_next_pc\[21\] _07948_ _08218_ _08230_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__a22o_1
X_11786_ reg_pc\[30\] _06322_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__and2_1
XANTENNA__10144__S0 _04758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16313_ _02883_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__clkbuf_1
X_13525_ _04466_ _07315_ _07339_ _07254_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__o211a_1
X_10737_ _05243_ _05330_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__and2b_1
X_17293_ clknet_leaf_100_clk _00467_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15939__C mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15083__S0 _03669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14735__B1 _07877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16244_ _02846_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13456_ _04160_ _07315_ _07316_ _07216_ VGND VGND VPWR VPWR _07317_ sky130_fd_sc_hd__o211a_1
X_10668_ _03607_ _05222_ _05220_ _03608_ _05368_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__a221o_1
XFILLER_0_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11549__B1 _06098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12407_ cpuregs.regs\[27\]\[7\] _06548_ _06678_ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10447__S1 _04473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16175_ net281 net243 _02797_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__mux2_1
X_10599_ _05300_ _05301_ _05220_ _03535_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__a22o_1
X_13387_ _04039_ _04198_ _05257_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__mux2_1
XANTENNA__09611__C1 _04149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16831__S _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput107 net107 VGND VGND VPWR VPWR cpi_rs2[17] sky130_fd_sc_hd__buf_1
XFILLER_0_23_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput118 net118 VGND VGND VPWR VPWR cpi_rs2[27] sky130_fd_sc_hd__clkbuf_1
XANTENNA__08560__D _03338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15126_ cpuregs.regs\[16\]\[5\] cpuregs.regs\[17\]\[5\] cpuregs.regs\[18\]\[5\] cpuregs.regs\[19\]\[5\]
+ _01979_ _01980_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__mux4_1
Xoutput129 net129 VGND VGND VPWR VPWR cpi_rs2[8] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12338_ cpuregs.regs\[26\]\[7\] _06548_ _06641_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__mux2_1
XANTENNA__15386__S1 _01909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15057_ _03657_ _01916_ _03692_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__a21o_1
X_12269_ cpuregs.regs\[25\]\[7\] _06548_ _06604_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__mux2_1
X_14008_ _07771_ _07772_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__nor2_1
XANTENNA__13475__B _04382_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15138__S1 _01992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15971__A mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10180__A _04483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15959_ _03757_ _02678_ _02679_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__o21ai_1
XANTENNA__16278__S _02859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15182__S _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08500_ instr_lhu instr_lh VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09480_ _04209_ _04210_ _04211_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__mux2_1
XANTENNA__08585__A _03195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10383__S0 _04216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08431_ _03207_ _03216_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__and2_2
XFILLER_0_148_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17629_ clknet_leaf_113_clk _00798_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08879__S1 _03643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13529__A1 _07304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14726__B1 _07877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11004__A2 _05301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12046__S _06471_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16741__S _03075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15865__B _02613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10763__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13701__A1 _04913_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09355__S _04078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09816_ _04463_ _04501_ _04502_ _04464_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__or4b_1
XANTENNA__15454__A1 _02012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09747_ _04059_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08495__A mem_do_prefetch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09678_ cpuregs.regs\[28\]\[8\] cpuregs.regs\[29\]\[8\] cpuregs.regs\[30\]\[8\] cpuregs.regs\[31\]\[8\]
+ _04085_ _04087_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__mux4_1
XANTENNA__15206__A1 _01959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15206__B2 decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08629_ cpu_state\[5\] _03238_ _03251_ _03401_ is_sb_sh_sw VGND VGND VPWR VPWR _00079_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_96_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13768__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11640_ _06200_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__buf_2
XFILLER_0_37_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11571_ _06137_ _06138_ _06075_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__o21a_1
XANTENNA__09841__C1 _04149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_946 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15065__S0 _03670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13310_ _06997_ cpuregs.regs\[5\]\[26\] _07176_ VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15121__A _01918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10522_ net125 VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__14717__B1 _07877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14290_ _05941_ _06333_ _07944_ _05951_ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__o211a_2
XFILLER_0_135_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10453_ _05157_ _05158_ _04078_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__mux2_1
X_13241_ _07146_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16651__S _03062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15390__B1 _02027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13940__A1 _03358_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10384_ _05090_ _05091_ _04369_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__mux2_1
X_13172_ _06995_ cpuregs.regs\[4\]\[25\] _07104_ VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__mux2_1
XANTENNA__15368__S1 _01986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11951__A0 _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12123_ _06517_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_36_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17980_ clknet_leaf_44_clk _01117_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_36_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14496__A2 _07947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16931_ clknet_leaf_140_clk _00112_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12054_ _06248_ cpuregs.regs\[22\]\[19\] _06471_ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11005_ _05573_ _05601_ _05603_ _05570_ _05686_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__a221o_1
X_16862_ _03175_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15445__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18601_ clknet_leaf_177_clk _01666_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_15813_ _05960_ _03634_ _03878_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__and3_1
XANTENNA_output222_A net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16793_ _06575_ cpuregs.regs\[13\]\[20\] _03138_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__mux2_1
XANTENNA__15540__S1 _01991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15996__A2 _03636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18532_ clknet_leaf_116_clk _01597_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15744_ _04909_ _02506_ _02544_ _02545_ VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__o211a_1
X_12956_ _06991_ cpuregs.regs\[31\]\[23\] _06985_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11907_ _06208_ cpuregs.regs\[20\]\[14\] _06398_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__mux2_1
X_18463_ clknet_leaf_132_clk _01528_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_15675_ _04240_ _02477_ _02493_ _02494_ _07775_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__a221oi_1
X_12887_ _06095_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__buf_2
XANTENNA__11035__S _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17414_ clknet_leaf_18_clk _00583_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08555__D _03333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14626_ _08035_ _08277_ VGND VGND VPWR VPWR _08278_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _06216_ cpuregs.regs\[11\]\[15\] _06359_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__mux2_1
X_18394_ clknet_leaf_170_clk _01459_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17345_ clknet_leaf_10_clk _00514_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_14557_ _08196_ _08201_ _08213_ _08055_ VGND VGND VPWR VPWR _08215_ sky130_fd_sc_hd__a31o_1
X_11769_ reg_pc\[28\] _06306_ _06101_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08852__B net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13508_ _07363_ _07355_ _07364_ VGND VGND VPWR VPWR _07365_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17276_ clknet_leaf_7_clk _00450_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14488_ _08128_ _08139_ VGND VGND VPWR VPWR _08151_ sky130_fd_sc_hd__nor2_1
XANTENNA__08571__C _03348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16227_ net47 mem_16bit_buffer\[6\] _02831_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__mux2_1
X_13439_ _04456_ _07276_ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08938__A1 _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13931__A1 _03330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16158_ _02770_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15685__B _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15359__S1 _01992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15109_ _05288_ _01963_ _01965_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12390__A cpuregs.waddr\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16089_ is_jalr_addi_slti_sltiu_xori_ori_andi _02711_ _02754_ VGND VGND VPWR VPWR
+ _01348_ sky130_fd_sc_hd__o21a_1
X_08980_ _03740_ _03741_ _03203_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10622__B _05324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11170__A1 _04038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11170__B2 _03297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09601_ cpuregs.regs\[8\]\[6\] cpuregs.regs\[9\]\[6\] cpuregs.regs\[10\]\[6\] cpuregs.regs\[11\]\[6\]
+ _04329_ _04218_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__mux4_1
XANTENNA__16947__D _00075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09532_ net37 net54 _04039_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10356__S0 _04057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09463_ _04192_ _04193_ _04194_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_121_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14947__A0 net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08414_ net262 net65 _03198_ _03199_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09394_ cpuregs.regs\[24\]\[2\] cpuregs.regs\[25\]\[2\] cpuregs.regs\[26\]\[2\] cpuregs.regs\[27\]\[2\]
+ _04071_ _04073_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_35_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_31_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__08762__B net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15598__S1 _01909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10984__A1 _04848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08929__A1 _03657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13396__A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12504__S _06737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15675__A1 _04240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_98_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__15427__A1 _01959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15427__B2 decoded_imm\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13335__S _04211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12810_ _06902_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15116__A _01919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13790_ _07583_ _07614_ VGND VGND VPWR VPWR _07628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12459__B _06082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12741_ decoded_rd\[1\] _06863_ _06864_ VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11464__A2 irq_pending\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16646__S _03051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10672__A0 _04198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14938__A0 net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15460_ decoded_imm\[21\] _02216_ _02197_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__a21o_1
XFILLER_0_166_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12672_ _06105_ cpuregs.regs\[12\]\[2\] _06825_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14674__B _07969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14411_ _07998_ _08076_ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__or2_1
X_11623_ _06185_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__clkbuf_1
X_15391_ net107 _01906_ _02233_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__o21a_1
XANTENNA__09768__B _04493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13070__S _07046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_2
X_17130_ clknet_leaf_147_clk _00304_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14342_ decoded_imm_j\[3\] _07911_ VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__and2_1
X_11554_ _06120_ _06123_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__nor2_4
XFILLER_0_123_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15589__S1 _02222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10505_ instr_sra instr_srl instr_srai instr_srli VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__nor4_2
X_17061_ clknet_leaf_156_clk _00235_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14273_ reg_pc\[23\] _07953_ _07958_ _07935_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16381__S _02918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11485_ irq_mask\[30\] _03428_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_9 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14690__A _08335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16012_ is_sb_sh_sw mem_rdata_q\[7\] _02712_ mem_rdata_q\[20\] _02634_ VGND VGND
+ VPWR VPWR _02713_ sky130_fd_sc_hd__a221o_1
X_13224_ _07137_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__clkbuf_1
X_10436_ net88 VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09593__A1 _04206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13155_ _06978_ cpuregs.regs\[4\]\[17\] _07093_ VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__mux2_1
X_10367_ net86 VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12414__S _06689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15210__S0 _01973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16863__A0 _06578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12106_ _06184_ cpuregs.regs\[23\]\[11\] _06507_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13677__A0 _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13086_ _07064_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__clkbuf_1
X_17963_ clknet_leaf_191_clk _01100_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dfxtp_1
X_10298_ _04996_ _05000_ _04133_ _05008_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__o211a_4
XFILLER_0_97_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_89_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12037_ _06472_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__clkbuf_1
X_16914_ clknet_leaf_17_clk _00095_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11152__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17894_ clknet_leaf_93_clk _01063_ VGND VGND VPWR VPWR count_cycle\[39\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15418__A1 _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09440__S1 _04073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13753__B _05227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16845_ _03166_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15969__A2 _03636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08847__B net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16776_ _06559_ cpuregs.regs\[13\]\[12\] _03127_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__mux2_1
X_13988_ _06053_ VGND VGND VPWR VPWR _07759_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12101__A0 _06166_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15727_ timer\[17\] timer\[16\] timer\[18\] _02524_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__or4_2
XFILLER_0_34_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18515_ clknet_leaf_155_clk _01580_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_12939_ _06239_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_38_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15658_ _02477_ _02478_ _02480_ _02481_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18446_ clknet_leaf_112_clk _01511_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14584__B _07958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14609_ _08071_ _08256_ _08262_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18377_ clknet_leaf_99_clk _01442_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15589_ cpuregs.regs\[20\]\[29\] cpuregs.regs\[21\]\[29\] cpuregs.regs\[22\]\[29\]
+ cpuregs.regs\[23\]\[29\] _02221_ _02222_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_13_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17328_ clknet_leaf_164_clk _00502_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10966__A1 _05361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09820__A2 _04016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15354__B1 _02196_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17259_ clknet_leaf_150_clk _00433_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16291__S _02870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13904__A1 _03359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09033__A0 mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11915__A0 _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12324__S _06641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16854__A0 _06569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15201__S0 _03661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08963_ _03679_ _03716_ _03725_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__and3_2
XANTENNA__13668__B1 _03311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13944__A _07681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11143__A1 _03407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15862__C _02610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08894_ _00065_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__buf_4
XANTENNA__15409__A1 _02250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11143__B2 _04422_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08757__B net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13155__S _07093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_56_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14632__A2 _07947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09515_ _04193_ _04194_ _04192_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_151_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12994__S _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09446_ _04177_ _04178_ _04077_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09377_ net44 net258 _04035_ net41 _04111_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__a221o_1
XANTENNA__14396__B2 _08035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15440__S0 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11270_ reg_next_pc\[18\] reg_out\[18\] _05898_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__mux2_2
XANTENNA__10709__A1 _05361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_896 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09575__A1 _04272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10221_ _04932_ _04933_ _04430_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__mux2_1
XANTENNA__18132__D alu_out\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15648__A1 _03218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09670__S1 _04074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10152_ cpuregs.regs\[16\]\[21\] cpuregs.regs\[17\]\[21\] cpuregs.regs\[18\]\[21\]
+ cpuregs.regs\[19\]\[21\] _04579_ _04284_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__mux4_1
Xoutput290 net290 VGND VGND VPWR VPWR mem_wdata[5] sky130_fd_sc_hd__clkbuf_1
XANTENNA__15545__S _03713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14960_ _01855_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__clkbuf_1
X_10083_ cpuregs.regs\[12\]\[19\] cpuregs.regs\[13\]\[19\] cpuregs.regs\[14\]\[19\]
+ cpuregs.regs\[15\]\[19\] _04273_ _04283_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_7_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14669__B _07969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13911_ _07681_ VGND VGND VPWR VPWR _07705_ sky130_fd_sc_hd__buf_2
X_14891_ _03631_ _01814_ _01815_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__nor3_1
XANTENNA__08667__B net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16073__A1 decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16630_ cpuregs.regs\[1\]\[10\] _06174_ _03051_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__mux2_1
XANTENNA__16073__B2 mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13842_ _07660_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_18_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14084__B1 _07790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16561_ _03003_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__clkbuf_8
X_13773_ _07609_ _07610_ _07608_ VGND VGND VPWR VPWR _07612_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_48_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10985_ _05667_ _05617_ _05243_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__mux2_1
XANTENNA__16376__S _02907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10645__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15512_ _02342_ _02344_ _02347_ _02037_ _01969_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18300_ clknet_leaf_5_clk _01368_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dfxtp_1
X_12724_ _06312_ cpuregs.regs\[12\]\[27\] _06847_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__mux2_1
X_16492_ _02978_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__clkbuf_1
X_18231_ clknet_leaf_16_clk _01302_ VGND VGND VPWR VPWR decoded_rd\[4\] sky130_fd_sc_hd__dfxtp_1
X_15443_ _02020_ _02274_ _02282_ _01960_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__o211a_2
XFILLER_0_154_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12655_ _06312_ cpuregs.regs\[30\]\[27\] _06810_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10718__A _05416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12409__S _06678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09489__S1 _04219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11606_ _06116_ reg_next_pc\[10\] _06169_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18162_ clknet_leaf_24_clk _01233_ VGND VGND VPWR VPWR decoded_imm_j\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09263__A0 mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15374_ net106 _02081_ _02215_ _02217_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_61_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12586_ _06781_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09802__A2 _04308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17113_ clknet_leaf_171_clk _00287_ VGND VGND VPWR VPWR cpuregs.regs\[24\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14325_ _08001_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15336__B1 _01963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18093_ clknet_leaf_102_clk _01197_ VGND VGND VPWR VPWR timer\[8\] sky130_fd_sc_hd__dfxtp_1
X_11537_ _06098_ _06107_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12933__A _06223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15431__S0 _02030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17044_ clknet_leaf_112_clk _00218_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14256_ _07904_ VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__clkbuf_4
X_11468_ _06041_ irq_pending\[22\] _06052_ net15 VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13207_ _07128_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09566__A1 _04289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10419_ cpuregs.regs\[20\]\[29\] cpuregs.regs\[21\]\[29\] cpuregs.regs\[22\]\[29\]
+ cpuregs.regs\[23\]\[29\] _04477_ _04478_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__mux4_1
X_14187_ count_instr\[62\] _07893_ count_instr\[63\] VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10176__A2 _04145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11399_ _03767_ _03833_ _03947_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15639__A1 decoder_trigger VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13138_ _06961_ cpuregs.regs\[4\]\[9\] _07082_ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__mux2_1
Xalphacore_330 VGND VGND VPWR VPWR alphacore_330/HI cpi_insn[28] sky130_fd_sc_hd__conb_1
Xalphacore_341 VGND VGND VPWR VPWR alphacore_341/HI trace_data[2] sky130_fd_sc_hd__conb_1
Xalphacore_352 VGND VGND VPWR VPWR alphacore_352/HI trace_data[13] sky130_fd_sc_hd__conb_1
Xalphacore_363 VGND VGND VPWR VPWR alphacore_363/HI trace_data[24] sky130_fd_sc_hd__conb_1
X_17946_ clknet_leaf_78_clk _08387_ VGND VGND VPWR VPWR reg_out\[26\] sky130_fd_sc_hd__dfxtp_1
X_13069_ _07055_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__clkbuf_1
Xalphacore_374 VGND VGND VPWR VPWR alphacore_374/HI trace_data[35] sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_2_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10333__C1 _03302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17877_ clknet_leaf_88_clk _01046_ VGND VGND VPWR VPWR count_cycle\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08577__B irq_pending\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11284__A reg_next_pc\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15498__S0 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16828_ _03157_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14075__B1 _07790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16286__S _02859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16759_ _06542_ cpuregs.regs\[13\]\[4\] _03116_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09300_ net67 VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15190__S _03664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09231_ _03862_ _03864_ _03882_ _03966_ _03786_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__a32o_1
XFILLER_0_173_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18429_ clknet_leaf_184_clk _01494_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12319__S _06603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13004__A _07009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09162_ mem_rdata_q\[17\] _03913_ _03914_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10939__A1 _05281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09093_ _03767_ _03768_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__nor2_2
XFILLER_0_142_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15422__S0 _03661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12054__S _06471_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10167__A2 _04880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09995_ reg_pc\[17\] decoded_imm\[17\] VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__nand2_1
X_08946_ _03666_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11116__A1 _05143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09404__S1 _04124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _00065_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15489__S0 _03661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16055__A1 decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11419__A2 _03920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09599__A _04123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10770_ net128 net96 VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09429_ net55 net258 _04035_ net42 _04162_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15566__B1 _02397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__18127__D alu_out\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10538__A net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15030__A2 _04022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12440_ _06703_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_136_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09340__S0 _04072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12371_ _06666_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14110_ count_instr\[39\] count_instr\[35\] _07831_ _07839_ VGND VGND VPWR VPWR _07843_
+ sky130_fd_sc_hd__and4_2
XANTENNA__15869__B2 _02625_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11322_ _05909_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15090_ _03719_ _01946_ _01948_ _00067_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__o211a_1
X_14041_ count_instr\[18\] count_instr\[17\] count_instr\[16\] VGND VGND VPWR VPWR
+ _07795_ sky130_fd_sc_hd__and3_1
X_11253_ reg_next_pc\[15\] reg_out\[15\] _05876_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_1001 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10158__A2 _04871_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10204_ reg_pc\[23\] decoded_imm\[23\] VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__nand2_1
X_11184_ _05828_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__buf_4
X_17800_ clknet_leaf_57_clk _00969_ VGND VGND VPWR VPWR reg_pc\[8\] sky130_fd_sc_hd__dfxtp_2
X_10135_ _03637_ _04848_ _04048_ irq_pending\[20\] _04850_ VGND VGND VPWR VPWR _04851_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15992_ _06016_ _05991_ _02706_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__a21o_1
XANTENNA__08678__A net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10066_ reg_pc\[19\] decoded_imm\[19\] VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__or2_1
X_14943_ net206 net175 _01846_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__mux2_1
X_17731_ clknet_leaf_101_clk _00900_ VGND VGND VPWR VPWR count_instr\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16046__A1 decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17662_ clknet_leaf_72_clk _00831_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dfxtp_4
X_14874_ _01803_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10330__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_1011 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13825_ cpuregs.regs\[0\]\[9\] VGND VGND VPWR VPWR _07652_ sky130_fd_sc_hd__clkbuf_1
X_16613_ cpuregs.regs\[1\]\[2\] _06104_ _03040_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__mux2_1
X_17593_ clknet_leaf_161_clk _00762_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16544_ _03006_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_63_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13756_ _07281_ _07595_ _07282_ reg_pc\[27\] _07283_ VGND VGND VPWR VPWR _07596_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_63_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10968_ _05651_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12707_ _06248_ cpuregs.regs\[12\]\[19\] _06836_ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16475_ cpuregs.regs\[17\]\[1\] _06536_ _02968_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13687_ _03575_ _07277_ VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12139__S _06518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10899_ _05288_ _05455_ _05587_ _05298_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15021__A2 _01863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18214_ clknet_leaf_43_clk _01285_ VGND VGND VPWR VPWR instr_or sky130_fd_sc_hd__dfxtp_2
XFILLER_0_116_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15426_ _02005_ _02262_ _02266_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12638_ _06248_ cpuregs.regs\[30\]\[19\] _06799_ VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13032__A1 _06582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15958__B _03218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11978__S _06435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18145_ clknet_leaf_49_clk alu_out\[19\] VGND VGND VPWR VPWR alu_out_q\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15357_ _01989_ _02200_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__or2_1
X_12569_ _06772_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15404__S0 _03640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14308_ _03379_ _07984_ VGND VGND VPWR VPWR _07985_ sky130_fd_sc_hd__or2_1
X_18076_ clknet_leaf_75_clk _01181_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfxtp_4
X_15288_ cpuregs.regs\[0\]\[12\] cpuregs.regs\[1\]\[12\] cpuregs.regs\[2\]\[12\] cpuregs.regs\[3\]\[12\]
+ _01973_ _01974_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17027_ clknet_leaf_130_clk _00201_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14239_ _03294_ VGND VGND VPWR VPWR _07935_ sky130_fd_sc_hd__buf_2
XANTENNA__09539__B2 _04013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12813__D cpuregs.waddr\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15974__A _03965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ net75 VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_74_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _04501_ _04502_ _04503_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08588__A instr_waitirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08731_ net102 net70 VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__nor2_1
X_17929_ clknet_leaf_65_clk _08400_ VGND VGND VPWR VPWR reg_out\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16037__A1 decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08662_ irq_mask\[0\] _03428_ irq_pending\[0\] _03305_ VGND VGND VPWR VPWR _03429_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09711__B2 _04206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08593_ _03277_ _03247_ _03365_ _03371_ _03298_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__a32o_1
XANTENNA__10609__A0 _05013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11742__A reg_pc\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15214__A _03709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15548__B1 _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09214_ _03782_ _03869_ _03736_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_170_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11034__A0 _05013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11888__S _06387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09145_ mem_rdata_q\[24\] _03900_ _03846_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08770__B net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08450__A1 mem_do_wdata VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09076_ _03788_ _03837_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14523__A1 _07898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10093__A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13731__C1 _07217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09978_ cpuregs.regs\[0\]\[16\] cpuregs.regs\[1\]\[16\] cpuregs.regs\[2\]\[16\] cpuregs.regs\[3\]\[16\]
+ _04487_ _04469_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__mux4_1
XANTENNA__12512__S _06737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14287__B1 _07967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08498__A _03277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08929_ _03657_ _03691_ _03692_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_129_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16028__A1 decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15823__S _03635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09702__B2 _04014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11940_ _06336_ cpuregs.regs\[20\]\[30\] _06386_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14039__B1 _07675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11871_ _06343_ cpuregs.regs\[11\]\[31\] _06347_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13610_ net75 decoded_imm\[17\] VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ _05507_ _05509_ _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__and3_1
XANTENNA__09466__A0 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15124__A _01918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14590_ _08241_ _08243_ _08244_ VGND VGND VPWR VPWR _08245_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13541_ net68 decoded_imm\[10\] _07377_ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10753_ _03522_ _03546_ _03547_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16260_ _02854_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__clkbuf_1
X_13472_ _04532_ _07276_ VGND VGND VPWR VPWR _07332_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10684_ _05381_ _05384_ _03530_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__17696__D _00865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15211_ cpuregs.regs\[4\]\[8\] cpuregs.regs\[5\]\[8\] cpuregs.regs\[6\]\[8\] cpuregs.regs\[7\]\[8\]
+ _01976_ _01977_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__mux4_1
XANTENNA__11025__B1 _05215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12423_ _06694_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16191_ net296 _01822_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__or2_1
XANTENNA__09769__B2 _04023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09776__B decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11576__A1 alu_out_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15142_ _03647_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__buf_8
XANTENNA__09864__S1 _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12354_ _06657_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11305_ _05927_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14514__A1 decoded_imm_j\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15073_ _01932_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__buf_4
XFILLER_0_132_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12285_ _06620_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14024_ count_instr\[12\] _07781_ _07783_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11236_ reg_next_pc\[12\] reg_out\[12\] _05858_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08900__S _03664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13518__S _07374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11167_ net116 _04710_ _05818_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__a21o_2
XANTENNA__12422__S _06689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15475__C1 _02027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10118_ cpuregs.regs\[24\]\[20\] cpuregs.regs\[25\]\[20\] cpuregs.regs\[26\]\[20\]
+ cpuregs.regs\[27\]\[20\] _04275_ _04278_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__mux4_1
X_11098_ _05770_ _05771_ _05772_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__o21a_1
X_15975_ _05998_ _02692_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__nor2_1
XANTENNA__16829__S _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17714_ clknet_leaf_76_clk _00883_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10049_ _04231_ _04766_ _04082_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__a21o_1
X_14926_ net198 net167 _01835_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15227__C1 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17645_ clknet_leaf_47_clk _00814_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfxtp_4
X_14857_ count_cycle\[52\] count_cycle\[53\] count_cycle\[54\] _01786_ VGND VGND VPWR
+ VPWR _01792_ sky130_fd_sc_hd__and4_1
X_13808_ _07643_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__clkbuf_1
X_14788_ count_cycle\[32\] count_cycle\[31\] _01741_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__and3_1
X_17576_ clknet_leaf_172_clk _00745_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_11_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13739_ _07578_ _07579_ VGND VGND VPWR VPWR _07580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16527_ cpuregs.regs\[17\]\[26\] _06588_ _02990_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16564__S _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15625__S0 _03640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09209__A0 mem_rdata_q\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13005__A1 _06554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16458_ _02960_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15409_ net108 _02250_ _01905_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16389_ _06995_ cpuregs.regs\[16\]\[25\] _02918_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11567__A1 _06072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09855__S1 _04513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18128_ clknet_leaf_26_clk alu_out\[2\] VGND VGND VPWR VPWR alu_out_q\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18059_ clknet_leaf_73_clk _01164_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_123_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09901_ cpuregs.regs\[16\]\[14\] cpuregs.regs\[17\]\[14\] cpuregs.regs\[18\]\[14\]
+ cpuregs.regs\[19\]\[14\] _04329_ _04218_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__mux4_1
XANTENNA__09906__S _04369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09832_ cpuregs.regs\[20\]\[12\] cpuregs.regs\[21\]\[12\] cpuregs.regs\[22\]\[12\]
+ cpuregs.regs\[23\]\[12\] _04084_ _04086_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__mux4_1
XANTENNA__09393__C1 _04068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_171_Right_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12332__S _06641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14269__B1 _07942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_141_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16031__C _02610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09763_ cpuregs.regs\[8\]\[10\] cpuregs.regs\[9\]\[10\] cpuregs.regs\[10\]\[10\]
+ cpuregs.regs\[11\]\[10\] _04487_ _04469_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__mux4_1
XANTENNA__16739__S _03075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08714_ net108 net76 VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__or2_1
X_09694_ _04031_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15870__C _03940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09641__S _04369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13671__B _05257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08645_ irq_mask\[2\] _03412_ irq_pending\[2\] _03304_ VGND VGND VPWR VPWR _03413_
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_156_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08576_ _03351_ _03352_ _03353_ _03354_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_25_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11255__A0 _04642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15092__S1 _03646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09128_ _03883_ _03884_ _03885_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__o21a_1
XFILLER_0_162_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08423__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10230__A1 _04271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09059_ _03819_ _03820_ _03231_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12070_ _06489_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16249__A1 _03213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11021_ _05476_ _05700_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13338__S _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18140__D alu_out\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12242__S _06576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15119__A _01919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10551__A _05254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11366__B _03213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15760_ timer\[27\] VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _07002_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08956__A _03713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13483__B2 reg_pc\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13581__B decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14711_ count_cycle\[7\] count_cycle\[8\] _08346_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__and3_1
XANTENNA__10297__B2 _04206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11923_ _06411_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15691_ _02486_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08675__B net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13073__S _07057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17430_ clknet_leaf_97_clk _00599_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_14642_ _07966_ _07988_ _08277_ VGND VGND VPWR VPWR _08293_ sky130_fd_sc_hd__and3_1
X_11854_ _06373_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10049__A1 _04231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10805_ _03512_ _03515_ _03549_ _03552_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__a31oi_1
X_17361_ clknet_leaf_151_clk _00530_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13330__S1 _04208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14573_ _08012_ _08228_ _08229_ VGND VGND VPWR VPWR _08230_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11785_ _06329_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15607__S0 _01908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10144__S1 _04759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13524_ _07378_ _07379_ VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09787__A _04273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16312_ _06987_ cpuregs.regs\[15\]\[21\] _02881_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__mux2_1
X_10736_ _05226_ _05259_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17292_ clknet_leaf_152_clk _00466_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08691__A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15083__S1 _03646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16243_ net56 mem_16bit_buffer\[14\] _02830_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__mux2_1
X_13455_ _04466_ _05209_ VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__or2_1
X_10667_ _03606_ _05367_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11549__A1 _06072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12406_ _06685_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08414__A1 net262 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16174_ _02805_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__clkbuf_1
X_13386_ _07209_ _07250_ _07211_ reg_pc\[2\] VGND VGND VPWR VPWR _07251_ sky130_fd_sc_hd__a22o_1
XANTENNA__08414__B2 _03199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10598_ _05213_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15125_ _01919_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__buf_8
Xoutput108 net108 VGND VGND VPWR VPWR cpi_rs2[18] sky130_fd_sc_hd__buf_1
X_12337_ _06648_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__clkbuf_1
Xoutput119 net119 VGND VGND VPWR VPWR cpi_rs2[28] sky130_fd_sc_hd__buf_1
XFILLER_0_121_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15056_ _01914_ _01915_ _03664_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__mux2_1
X_12268_ _06611_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13248__S _07140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14007_ count_instr\[7\] _07769_ _07759_ VGND VGND VPWR VPWR _07772_ sky130_fd_sc_hd__o21ai_1
X_11219_ _05856_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_71_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12199_ cpuregs.regs\[24\]\[15\] _06565_ _06555_ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__mux2_1
Xoutput90 net90 VGND VGND VPWR VPWR cpi_rs1[30] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_71_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11276__B _05899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10080__S0 _04512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15971__B _02610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16559__S _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15999__B1 _03763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11991__S _06446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15958_ mem_do_wdata _03218_ _03219_ _03233_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__or4_1
XANTENNA__08866__A _03309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14909_ net220 net189 _01824_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__mux2_1
X_15889_ instr_lw _02635_ _02639_ is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR _01263_
+ sky130_fd_sc_hd__a22o_1
X_08430_ _03203_ mem_la_firstword_reg last_mem_valid VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__mux2_1
XANTENNA__10383__S1 _04376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17628_ clknet_leaf_106_clk _00797_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15620__C1 _03654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17559_ clknet_leaf_118_clk _00728_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13529__A2 _04526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16479__A1 _06540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10763__A2 _03524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13666__B decoded_imm\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13162__A0 _06984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09366__C1 _04100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13701__A2 decoded_imm\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13367__A2_N _04101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09815_ _04501_ _04503_ _04537_ _04538_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__o211ai_1
XANTENNA__16469__S _02931_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16651__A1 _06256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09746_ _04280_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09669__B1 _04013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11476__B1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09677_ _04070_ _04400_ _04404_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08495__B _03237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15206__A2 _02050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08628_ _03391_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__inv_2
XANTENNA__15611__C1 _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13768__A2 decoded_imm\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08559_ irq_mask\[0\] irq_pending\[0\] VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__and2b_2
XFILLER_0_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11570_ reg_pc\[5\] _06121_ reg_pc\[6\] VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10521_ _05218_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__inv_2
XANTENNA__15065__S1 _03671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12728__A0 _06328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13240_ _06995_ cpuregs.regs\[8\]\[25\] _07140_ VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10452_ cpuregs.regs\[24\]\[30\] cpuregs.regs\[25\]\[30\] cpuregs.regs\[26\]\[30\]
+ cpuregs.regs\[27\]\[30\] _04085_ _04087_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__mux4_1
XANTENNA__15390__A1 decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15390__B2 _02232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10203__A1 _04391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13171_ _07109_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__clkbuf_1
X_10383_ cpuregs.regs\[28\]\[28\] cpuregs.regs\[29\]\[28\] cpuregs.regs\[30\]\[28\]
+ cpuregs.regs\[31\]\[28\] _04216_ _04376_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_972 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15678__C1 _07775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12122_ _06248_ cpuregs.regs\[23\]\[19\] _06507_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13068__S _07046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16930_ clknet_leaf_142_clk _00111_ VGND VGND VPWR VPWR cpuregs.regs\[10\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_12053_ _06480_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11004_ _03470_ _05301_ _05215_ _03473_ _05685_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__a221o_1
XANTENNA__09372__A2 _04012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16861_ _06575_ cpuregs.regs\[14\]\[20\] _03174_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__mux2_1
XANTENNA__16379__S _02918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16642__A1 _06223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18600_ clknet_leaf_138_clk _01665_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_15812_ decoded_imm_j\[6\] _05983_ _03965_ _02587_ _02589_ VGND VGND VPWR VPWR _01236_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__13456__A1 _04160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16792_ _03115_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__buf_4
X_18531_ clknet_leaf_157_clk _01596_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_15743_ _07778_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__buf_2
X_12955_ _06280_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__buf_2
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output215_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11906_ _06402_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18462_ clknet_leaf_182_clk _01527_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12886_ _06944_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__clkbuf_1
X_15674_ timer\[4\] _02490_ _02488_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_169_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17413_ clknet_leaf_1_clk _00582_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11837_ _06364_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14625_ _07961_ _07964_ _08258_ VGND VGND VPWR VPWR _08277_ sky130_fd_sc_hd__and3_1
XFILLER_0_173_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18393_ clknet_leaf_1_clk _01458_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12936__A _06231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13531__S _07374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15312__A _02012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17344_ clknet_leaf_10_clk _00513_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14556_ _08196_ _08201_ _08213_ VGND VGND VPWR VPWR _08214_ sky130_fd_sc_hd__a21oi_1
X_11768_ reg_pc\[28\] _06306_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13507_ net68 decoded_imm\[10\] VGND VGND VPWR VPWR _07364_ sky130_fd_sc_hd__xnor2_1
X_10719_ _05417_ _05283_ _05295_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16842__S _03163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17275_ clknet_leaf_16_clk _00449_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14487_ _08148_ _08149_ VGND VGND VPWR VPWR _08150_ sky130_fd_sc_hd__nand2_1
X_11699_ _06065_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__buf_2
XFILLER_0_82_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11051__S _05230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08571__D _03349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13438_ _07297_ _07298_ _07296_ VGND VGND VPWR VPWR _07300_ sky130_fd_sc_hd__a21o_1
X_16226_ _02837_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11986__S _06435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16157_ _02796_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__clkbuf_1
X_13369_ _03399_ _07234_ VGND VGND VPWR VPWR _07235_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15108_ _03396_ _03703_ _01964_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__a21oi_2
X_16088_ is_alu_reg_imm _02619_ _02634_ instr_jalr VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__a211o_1
XANTENNA__12390__B cpuregs.waddr\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15039_ _05138_ _01863_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13695__A1 _07274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14892__B1 _07274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16289__S _02870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11170__A2 _05292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09600_ cpuregs.regs\[12\]\[6\] cpuregs.regs\[13\]\[6\] cpuregs.regs\[14\]\[6\] cpuregs.regs\[15\]\[6\]
+ _04329_ _04218_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_108_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_1008 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09531_ _03524_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_88_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18729_ net124 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11458__B1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10356__S1 _04060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09462_ _04192_ _04193_ _04194_ _04156_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__a31o_1
XANTENNA__10130__B1 _04009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08413_ mem_do_rinst VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__buf_4
XANTENNA__14947__A1 net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09393_ _04121_ _04122_ _04126_ _04068_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15222__A _01995_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10433__B2 _04187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12057__S _06482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10984__A2 _04810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11896__S _06387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09874__B decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13396__B decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10292__S0 _04217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15675__A2 _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13686__A1 _04754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15427__A2 _02259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12520__S _06737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14635__B1 _07997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09729_ net98 VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__buf_4
XFILLER_0_97_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12740_ cpuregs.waddr\[0\] _06862_ _06865_ _06861_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10672__A1 _04262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12671_ _06827_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _08071_ _08074_ _08075_ _08079_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__a31o_1
X_11622_ _06184_ cpuregs.regs\[10\]\[11\] _06176_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08617__A1 irq_mask\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15390_ decoded_imm\[17\] _02216_ _02027_ _02232_ _02197_ VGND VGND VPWR VPWR _02233_
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_64_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14341_ _07911_ _08004_ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11553_ _06121_ _06122_ _06075_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10504_ _05180_ _05181_ _05208_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__o21ai_1
X_17060_ clknet_leaf_157_clk _00234_ VGND VGND VPWR VPWR cpuregs.regs\[22\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14272_ reg_next_pc\[23\] _05898_ _07942_ _07957_ VGND VGND VPWR VPWR _07958_ sky130_fd_sc_hd__o211a_2
X_11484_ _06054_ irq_pending\[29\] _06061_ net22 VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16011_ instr_jalr is_lb_lh_lw_lbu_lhu is_alu_reg_imm VGND VGND VPWR VPWR _02712_
+ sky130_fd_sc_hd__or3_2
XFILLER_0_123_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09578__C1 _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13223_ _06978_ cpuregs.regs\[8\]\[17\] _07129_ VGND VGND VPWR VPWR _07137_ sky130_fd_sc_hd__mux2_1
X_10435_ _04010_ _05121_ _05141_ _04150_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10188__B1 _04068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13154_ _07100_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10283__S0 _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16312__A0 _06987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10366_ _05070_ _05071_ _05074_ _03302_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13126__A0 _06949_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12105_ _06508_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15210__S1 _01974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13085_ _06976_ cpuregs.regs\[7\]\[16\] _07057_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__mux2_1
X_17962_ clknet_leaf_191_clk _01099_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dfxtp_1
X_10297_ _05002_ _05004_ _05007_ _04206_ _04296_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__a221o_1
X_16913_ clknet_leaf_40_clk _00094_ VGND VGND VPWR VPWR last_mem_valid sky130_fd_sc_hd__dfxtp_1
X_12036_ _06175_ cpuregs.regs\[22\]\[10\] _06471_ VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__mux2_1
XANTENNA__11688__B1 _06101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17893_ clknet_leaf_93_clk _01062_ VGND VGND VPWR VPWR count_cycle\[38\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10586__S1 _05239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16615__A1 _06113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16844_ _06559_ cpuregs.regs\[14\]\[12\] _03163_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__mux2_1
XANTENNA__12430__S _06689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10360__B1 _04227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16775_ _03129_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16837__S _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13987_ count_instr\[1\] count_instr\[0\] _07755_ VGND VGND VPWR VPWR _07758_ sky130_fd_sc_hd__and3_1
X_18514_ clknet_leaf_128_clk _01579_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08566__D _03344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15726_ _02530_ timer\[18\] VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__and2b_1
XFILLER_0_125_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16379__A0 _06984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12938_ _06979_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18445_ clknet_leaf_160_clk _01510_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_66_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15657_ _07778_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_83_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _06934_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14608_ reg_next_pc\[24\] _07904_ _08260_ _03378_ _08261_ VGND VGND VPWR VPWR _08262_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__13601__A1 _04566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18376_ clknet_leaf_180_clk _01441_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09805__B1 _03252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15588_ _02417_ _02418_ _02110_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09900__S0 _04329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17327_ clknet_leaf_121_clk _00501_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16572__S _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10186__A _04369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14539_ _08196_ _08197_ VGND VGND VPWR VPWR _08198_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15354__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17258_ clknet_leaf_140_clk _00432_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_945 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16209_ _06081_ _06862_ _02826_ decoded_rd\[4\] VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09033__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17189_ clknet_leaf_148_clk _00363_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12605__S _06788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15201__S1 _03662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08962_ _03683_ _03720_ _03724_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__a21o_1
XANTENNA__11679__B1 reg_pc\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09967__S0 _04281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08893_ _00064_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11143__A2 _05414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12340__S _06641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15217__A _01936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10351__B1 _04225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09514_ reg_pc\[4\] decoded_imm\[4\] VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09445_ cpuregs.regs\[0\]\[3\] cpuregs.regs\[1\]\[3\] cpuregs.regs\[2\]\[3\] cpuregs.regs\[3\]\[3\]
+ _04084_ _04086_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__mux4_1
XANTENNA__11851__A0 _06266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08773__B net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09376_ _04037_ _04038_ _04110_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__and3_1
XFILLER_0_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15887__A _02612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15440__S1 _01997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10824__A instr_sub VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10220_ cpuregs.regs\[28\]\[23\] cpuregs.regs\[29\]\[23\] cpuregs.regs\[30\]\[23\]
+ cpuregs.regs\[31\]\[23\] _04281_ _04470_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__mux4_1
XANTENNA__10543__B _05230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13108__A0 _06999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11382__A2 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10151_ cpuregs.regs\[20\]\[21\] cpuregs.regs\[21\]\[21\] cpuregs.regs\[22\]\[21\]
+ cpuregs.regs\[23\]\[21\] _04579_ _04284_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__mux4_1
XANTENNA__10590__A0 _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput280 net280 VGND VGND VPWR VPWR mem_wdata[25] sky130_fd_sc_hd__clkbuf_1
Xoutput291 net291 VGND VGND VPWR VPWR mem_wdata[6] sky130_fd_sc_hd__clkbuf_1
X_10082_ _04797_ _04798_ _04575_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ _07677_ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__buf_2
XANTENNA__15127__A _01907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14890_ _07633_ _07636_ _01813_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__o21a_1
X_13841_ cpuregs.regs\[0\]\[17\] VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16657__S _03062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14966__A _06186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13772_ _07608_ _07609_ _07610_ VGND VGND VPWR VPWR _07611_ sky130_fd_sc_hd__or3_1
X_16560_ _03014_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__clkbuf_1
X_10984_ _04880_ _04848_ _04810_ _04754_ _05264_ _05235_ VGND VGND VPWR VPWR _05667_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_48_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10645__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15511_ _02345_ _02346_ _02002_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__mux2_1
X_12723_ _06854_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16491_ cpuregs.regs\[17\]\[9\] _06552_ _02968_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13081__S _07057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11390__A _03954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18230_ clknet_leaf_9_clk _01301_ VGND VGND VPWR VPWR decoded_rd\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12654_ _06817_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__clkbuf_1
X_15442_ _02088_ _02277_ _02279_ _02281_ _02018_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11605_ irq_state\[1\] _03333_ _06098_ _06168_ _06074_ VGND VGND VPWR VPWR _06169_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18161_ clknet_leaf_23_clk _01232_ VGND VGND VPWR VPWR decoded_imm_j\[2\] sky130_fd_sc_hd__dfxtp_1
X_15373_ decoded_imm\[16\] _02216_ _02197_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ cpuregs.regs\[2\]\[26\] _06588_ _06774_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__mux2_1
XANTENNA__09263__A1 _04000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17112_ clknet_leaf_176_clk _00286_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15336__A1 decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14324_ _07991_ _08000_ VGND VGND VPWR VPWR _08001_ sky130_fd_sc_hd__or2_1
X_11536_ reg_out\[3\] alu_out_q\[3\] latched_stalu VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18092_ clknet_leaf_100_clk _01196_ VGND VGND VPWR VPWR timer\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14255_ _05909_ _06237_ _07945_ reg_next_pc\[18\] VGND VGND VPWR VPWR _07946_ sky130_fd_sc_hd__o22a_2
X_17043_ clknet_leaf_20_clk _00217_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15431__S1 _02031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11467_ irq_mask\[22\] _06042_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13898__A1 _03321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_915 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14206__A _03294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13206_ _06961_ cpuregs.regs\[8\]\[9\] _07118_ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10418_ _04054_ _05124_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__nand2_1
XANTENNA__10256__S0 _04290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14186_ count_instr\[62\] _07893_ _07895_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__o21a_1
X_11398_ _03867_ _03923_ _03971_ _03880_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13137_ _07091_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15195__S0 _02046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10349_ cpuregs.regs\[16\]\[27\] cpuregs.regs\[17\]\[27\] cpuregs.regs\[18\]\[27\]
+ cpuregs.regs\[19\]\[27\] _04207_ _04208_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__mux4_1
Xalphacore_320 VGND VGND VPWR VPWR alphacore_320/HI cpi_insn[18] sky130_fd_sc_hd__conb_1
Xalphacore_331 VGND VGND VPWR VPWR alphacore_331/HI cpi_insn[29] sky130_fd_sc_hd__conb_1
Xalphacore_342 VGND VGND VPWR VPWR alphacore_342/HI trace_data[3] sky130_fd_sc_hd__conb_1
Xalphacore_353 VGND VGND VPWR VPWR alphacore_353/HI trace_data[14] sky130_fd_sc_hd__conb_1
X_17945_ clknet_leaf_78_clk _08386_ VGND VGND VPWR VPWR reg_out\[25\] sky130_fd_sc_hd__dfxtp_1
X_13068_ _06959_ cpuregs.regs\[7\]\[8\] _07046_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__mux2_1
Xalphacore_364 VGND VGND VPWR VPWR alphacore_364/HI trace_data[25] sky130_fd_sc_hd__conb_1
Xalphacore_375 VGND VGND VPWR VPWR alphacore_375/HI trace_valid sky130_fd_sc_hd__conb_1
XANTENNA__13256__S _07154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15037__A _05106_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12019_ _06105_ cpuregs.regs\[22\]\[2\] _06460_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__mux2_1
X_17876_ clknet_leaf_88_clk _01045_ VGND VGND VPWR VPWR count_cycle\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11530__C1 _06101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16827_ _06542_ cpuregs.regs\[14\]\[4\] _03152_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__mux2_1
XANTENNA__15498__S1 _02014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16758_ _03120_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08874__A _00068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10636__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15709_ _04593_ _02506_ _02519_ _02481_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__o211a_1
X_16689_ _06955_ cpuregs.regs\[19\]\[6\] _03076_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__mux2_1
X_09230_ _03894_ _03948_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18428_ clknet_leaf_175_clk _01493_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16772__A0 _06554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13586__A0 _04532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09161_ _03846_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_155_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18359_ clknet_leaf_10_clk _01424_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09254__B2 _03888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09092_ mem_rdata_q\[20\] _03851_ _03846_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15422__S1 _03662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09994_ _03385_ _04685_ _04707_ _03303_ _04713_ VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08945_ cpuregs.regs\[12\]\[4\] cpuregs.regs\[13\]\[4\] cpuregs.regs\[14\]\[4\] cpuregs.regs\[15\]\[4\]
+ _03649_ _03643_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__mux4_1
XANTENNA__13166__S _07104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08876_ _03640_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_4_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15489__S1 _03662_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16477__S _02968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15263__B1 _02017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12077__A0 _06336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14605__A3 _07984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08784__A net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09428_ _04037_ _04038_ _04161_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__and3_1
XANTENNA__15566__A1 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15030__A3 _04979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09359_ _04092_ _04093_ _04064_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12370_ cpuregs.regs\[26\]\[22\] _06580_ _06663_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__mux2_1
XANTENNA__15318__B2 _02004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09340__S1 _04074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11321_ _05940_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_133_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10554__A _05257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12245__S _06533_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14040_ count_instr\[17\] _07792_ _07794_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11252_ _05829_ _05882_ _05883_ _05884_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__a31o_4
XFILLER_0_30_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1013 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10203_ _04391_ _04887_ _04888_ _04916_ VGND VGND VPWR VPWR _08383_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12552__A1 _06554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11183_ _04160_ _05826_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__mux2_1
X_10134_ _04709_ _04849_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__nor2_2
X_15991_ _05970_ _02701_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__nor2_1
XANTENNA__08678__B net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13501__B1 _07232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17730_ clknet_leaf_101_clk _00899_ VGND VGND VPWR VPWR count_instr\[1\] sky130_fd_sc_hd__dfxtp_1
X_10065_ reg_pc\[19\] decoded_imm\[19\] VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__nand2_1
X_14942_ _01823_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17661_ clknet_leaf_72_clk _00830_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dfxtp_4
X_14873_ _01801_ _01753_ _01802_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__and3b_1
XANTENNA__16387__S _02918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output128_A net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16612_ _03042_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__clkbuf_1
X_13824_ _07651_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13804__A1 _07232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17592_ clknet_leaf_161_clk _00761_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08694__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16543_ _06945_ cpuregs.regs\[18\]\[1\] _03004_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__mux2_1
X_10967_ _03477_ _05640_ _03476_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__a21o_1
X_13755_ _05069_ VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12706_ _06845_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__clkbuf_1
X_16474_ _02969_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__clkbuf_1
X_10898_ _05292_ _05586_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__or2_1
X_13686_ _04754_ _07236_ _07530_ _07217_ VGND VGND VPWR VPWR _07531_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18213_ clknet_leaf_41_clk _01284_ VGND VGND VPWR VPWR instr_sra sky130_fd_sc_hd__dfxtp_2
XFILLER_0_127_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_75_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15425_ _03654_ _02265_ _03675_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12637_ _06808_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15958__C _03219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18144_ clknet_leaf_47_clk alu_out\[18\] VGND VGND VPWR VPWR alu_out_q\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11043__A1 instr_sub VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12568_ cpuregs.regs\[2\]\[18\] _06571_ _06763_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__mux2_1
X_15356_ cpuregs.regs\[16\]\[16\] cpuregs.regs\[17\]\[16\] cpuregs.regs\[18\]\[16\]
+ cpuregs.regs\[19\]\[16\] _02013_ _02014_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_306 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12791__A1 _06578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11519_ _03195_ _06065_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__or2_1
X_14307_ _03319_ _07983_ VGND VGND VPWR VPWR _07984_ sky130_fd_sc_hd__and2_2
XANTENNA__15404__S1 _03642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18075_ clknet_leaf_75_clk _01180_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dfxtp_4
XANTENNA__10464__A _05169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15287_ cpuregs.regs\[4\]\[12\] cpuregs.regs\[5\]\[12\] cpuregs.regs\[6\]\[12\] cpuregs.regs\[7\]\[12\]
+ _01970_ _01971_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__mux4_1
X_12499_ _06240_ cpuregs.regs\[28\]\[18\] _06726_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__mux2_1
XANTENNA__16850__S _03163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09539__A2 _04016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17026_ clknet_leaf_181_clk _00200_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14238_ reg_next_pc\[13\] _05876_ _07922_ _07933_ VGND VGND VPWR VPWR _07934_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_78_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14169_ count_instr\[57\] count_instr\[56\] _07881_ VGND VGND VPWR VPWR _07884_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_111_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_84_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08730_ _03494_ _03495_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__or2b_2
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17928_ clknet_leaf_55_clk _08399_ VGND VGND VPWR VPWR reg_out\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16037__A2 _02711_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10857__A1 _05361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08661_ _03412_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__buf_2
XFILLER_0_56_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17859_ clknet_leaf_93_clk _01028_ VGND VGND VPWR VPWR count_cycle\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16297__S _02870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12059__A0 _06266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08592_ _03368_ _03370_ _03364_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__or3b_1
XANTENNA__15340__S0 _01976_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10609__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15548__A1 _01959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15548__B2 decoded_imm\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09213_ _03935_ _03880_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09227__A1 _03895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15230__A _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11034__A1 _04959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09144_ _03850_ _03828_ _03830_ _03849_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12782__A1 _06569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09075_ _03836_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12065__S _06482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14523__A2 _07943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13685__A _05044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08779__A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14287__A1 reg_pc\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09977_ cpuregs.regs\[4\]\[16\] cpuregs.regs\[5\]\[16\] cpuregs.regs\[6\]\[16\] cpuregs.regs\[7\]\[16\]
+ _04487_ _04469_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__mux4_1
XANTENNA__14287__B2 _07960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10313__S _04077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08928_ _00068_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09702__A2 _04016_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08859_ is_sltiu_bltu_sltu _03431_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__and2_1
XANTENNA__15787__A1 _03384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11870_ _06381_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15331__S0 _01999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10821_ _05399_ _05513_ _05514_ _05478_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_28_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09466__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10752_ _05432_ _05433_ _05449_ VGND VGND VPWR VPWR alu_out\[6\] sky130_fd_sc_hd__o21ai_2
X_13540_ _03510_ decoded_imm\[8\] _07352_ _07350_ VGND VGND VPWR VPWR _07395_ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15539__B2 _02017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13471_ _04342_ _05259_ VGND VGND VPWR VPWR _07331_ sky130_fd_sc_hd__or2_1
X_10683_ _05382_ _05383_ _05242_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14211__A1 reg_pc\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15210_ cpuregs.regs\[16\]\[8\] cpuregs.regs\[17\]\[8\] cpuregs.regs\[18\]\[8\] cpuregs.regs\[19\]\[8\]
+ _01973_ _01974_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__mux4_1
X_12422_ cpuregs.regs\[27\]\[14\] _06563_ _06689_ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__mux2_1
XANTENNA__15140__A _03669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09769__A2 _04021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10459__S0 _04280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16190_ _02812_ _02813_ _02814_ _02676_ net295 VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12353_ cpuregs.regs\[26\]\[14\] _06563_ _06652_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__mux2_1
X_15141_ _01995_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__buf_8
XFILLER_0_121_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10284__A _04430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11304_ _04959_ _05838_ _05926_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_133_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15072_ _01931_ is_jalr_addi_slti_sltiu_xori_ori_andi _03387_ VGND VGND VPWR VPWR
+ _01932_ sky130_fd_sc_hd__a21o_2
XFILLER_0_121_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12284_ cpuregs.regs\[25\]\[14\] _06563_ _06615_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14023_ count_instr\[12\] _07781_ _07775_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13595__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11235_ _05870_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_4
XANTENNA__12703__S _06836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08689__A net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ _04038_ _05286_ net130 _03297_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__a22o_1
XANTENNA__09941__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output245_A net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10117_ _04215_ _04832_ _04296_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__a21oi_2
X_11097_ _03441_ _05759_ _05517_ _03440_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__a211o_1
XANTENNA__15570__S0 _01976_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15974_ _03965_ _05999_ _06000_ _03977_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__or4b_1
XANTENNA__10839__A1 _05219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17713_ clknet_leaf_76_clk _00882_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dfxtp_1
X_10048_ _04764_ _04765_ _04065_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__mux2_1
X_14925_ _01837_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12939__A _06239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17644_ clknet_leaf_47_clk _00813_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfxtp_4
X_14856_ _01791_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15322__S0 _01979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13789__A0 _05174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13807_ cpuregs.regs\[0\]\[0\] VGND VGND VPWR VPWR _07643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09457__A1 _04168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17575_ clknet_leaf_180_clk _00744_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14787_ count_cycle\[31\] _01741_ _01744_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11999_ _06297_ cpuregs.regs\[21\]\[25\] _06446_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16526_ _02996_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__clkbuf_1
X_13738_ net85 decoded_imm\[26\] VGND VGND VPWR VPWR _07579_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14873__B _01753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11989__S _06446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15625__S1 _03642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16457_ _06995_ cpuregs.regs\[29\]\[25\] _02954_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__mux2_1
XANTENNA__09209__A1 _03763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13669_ _07499_ _07508_ _07513_ VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11016__A1 _05363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15408_ _01959_ _02241_ _02249_ _01933_ decoded_imm\[18\] VGND VGND VPWR VPWR _02250_
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_115_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16388_ _02923_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11567__A2 _03321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15985__A _03228_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18127_ clknet_leaf_29_clk alu_out\[1\] VGND VGND VPWR VPWR alu_out_q\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15339_ cpuregs.regs\[8\]\[15\] cpuregs.regs\[9\]\[15\] cpuregs.regs\[10\]\[15\]
+ cpuregs.regs\[11\]\[15\] _02030_ _02031_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__mux4_1
XANTENNA__15389__S0 _01968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16580__S _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09983__A _04051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18058_ clknet_leaf_73_clk _01163_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dfxtp_4
XANTENNA__10870__S0 _05264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11319__A2 _05937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09900_ cpuregs.regs\[20\]\[14\] cpuregs.regs\[21\]\[14\] cpuregs.regs\[22\]\[14\]
+ cpuregs.regs\[23\]\[14\] _04329_ _04218_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__mux4_1
X_17009_ clknet_leaf_160_clk _00183_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12613__S _06788_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09831_ _04553_ _04554_ _04369_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__mux2_1
XANTENNA__14269__A1 reg_next_pc\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09762_ cpuregs.regs\[12\]\[10\] cpuregs.regs\[13\]\[10\] cpuregs.regs\[14\]\[10\]
+ cpuregs.regs\[15\]\[10\] _04487_ _04469_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__mux4_1
XANTENNA__15561__S0 _02074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09145__A0 mem_rdata_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08713_ _03478_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__inv_2
X_09693_ latched_is_lb VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__inv_2
XANTENNA__09696__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09696__B2 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08644_ _03317_ _03409_ _03411_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__nand3_2
XANTENNA__15313__S0 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08575_ irq_mask\[28\] irq_pending\[28\] VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__and2b_1
XANTENNA__14977__C1 _08335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16755__S _03116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11899__S _06398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08781__B net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_926 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09127_ _03804_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10766__B1 _05251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10230__A2 _04941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09058_ net62 mem_rdata_q\[7\] _03200_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11020_ _05244_ _05228_ _05334_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_130_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15552__S0 _02030_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12971_ _07001_ cpuregs.regs\[31\]\[28\] _06985_ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__mux2_1
XANTENNA__13483__A2 _04415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15135__A _01936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14710_ count_cycle\[7\] _08346_ _08348_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__o21a_1
XFILLER_0_169_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12691__A0 _06184_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11922_ _06266_ cpuregs.regs\[20\]\[21\] _06409_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__mux2_1
X_15690_ _04415_ _02486_ _02504_ _02505_ _06026_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__o221a_1
XANTENNA__15304__S0 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14641_ _08290_ _08291_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__or2_1
X_11853_ _06274_ cpuregs.regs\[11\]\[22\] _06370_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__mux2_1
XANTENNA__10279__A _03384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14974__A _07208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16665__S _03062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10804_ _05498_ VGND VGND VPWR VPWR alu_out\[9\] sky130_fd_sc_hd__buf_1
X_17360_ clknet_leaf_154_clk _00529_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11784_ _06328_ cpuregs.regs\[10\]\[29\] _06258_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__mux2_1
X_14572_ _07954_ _07988_ _08209_ VGND VGND VPWR VPWR _08229_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16311_ _02882_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__clkbuf_1
X_13523_ _04466_ decoded_imm\[10\] _07365_ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__a21o_1
XANTENNA__15607__S1 _01909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10735_ _03522_ _05431_ _05218_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__16185__A1 net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17291_ clknet_leaf_154_clk _00465_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08662__A2 _03428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08691__B net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11602__S _06086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16242_ _02845_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__clkbuf_1
X_10666_ _05221_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__buf_4
X_13454_ _05257_ VGND VGND VPWR VPWR _07315_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_output195_A net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_149_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11549__A2 _03327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12405_ cpuregs.regs\[27\]\[6\] _06546_ _06678_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__mux2_1
X_13385_ _04142_ VGND VGND VPWR VPWR _07250_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16173_ net280 net242 _02797_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__mux2_1
X_10597_ _03242_ _05231_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__or2_2
XANTENNA__08414__A2 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15124_ _01918_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__clkbuf_16
Xoutput109 net109 VGND VGND VPWR VPWR cpi_rs2[19] sky130_fd_sc_hd__clkbuf_1
X_12336_ cpuregs.regs\[26\]\[6\] _06546_ _06641_ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15696__B1 _02476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12267_ cpuregs.regs\[25\]\[6\] _06546_ _06604_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__mux2_1
X_15055_ cpuregs.regs\[0\]\[0\] cpuregs.regs\[1\]\[0\] cpuregs.regs\[2\]\[0\] cpuregs.regs\[3\]\[0\]
+ _03658_ _03659_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__mux4_1
XANTENNA__10742__A _05398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09375__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output72_A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14006_ count_instr\[7\] count_instr\[6\] _07767_ VGND VGND VPWR VPWR _07771_ sky130_fd_sc_hd__and3_1
X_11218_ _03188_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__buf_2
XANTENNA__09914__A2 _04165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09308__A reg_next_pc\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12198_ _06215_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__buf_2
Xoutput80 net80 VGND VGND VPWR VPWR cpi_rs1[21] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput91 net91 VGND VGND VPWR VPWR cpi_rs1[31] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_71_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11721__A2 reg_next_pc\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11149_ _05809_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__buf_2
XANTENNA__11276__C _05902_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10080__S1 _04513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15543__S0 _03661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09027__B _03213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_158_Left_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15957_ mem_state\[0\] _02677_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__nand2_1
XANTENNA__08866__B _03384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13264__S _07154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11573__A _06140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15045__A _03272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14908_ _01828_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12682__A0 _06150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15888_ _02634_ _02638_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17627_ clknet_leaf_166_clk _00796_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_14839_ count_cycle\[46\] count_cycle\[47\] count_cycle\[48\] _01774_ VGND VGND VPWR
+ VPWR _01780_ sky130_fd_sc_hd__and4_2
XFILLER_0_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17558_ clknet_leaf_97_clk _00727_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13631__C1 _07232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08882__A _03646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16509_ _02987_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__clkbuf_1
X_17489_ clknet_leaf_134_clk _00658_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_167_Left_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14108__B _07815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10763__A3 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11748__A _06296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_165_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15439__B1 _01968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11712__A2 reg_next_pc\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09814_ reg_pc\[11\] decoded_imm\[11\] VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__nand2_1
XANTENNA__16100__B2 is_alu_reg_imm VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15534__S0 _01995_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14111__B1 _07834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09745_ cpuregs.regs\[24\]\[10\] cpuregs.regs\[25\]\[10\] cpuregs.regs\[26\]\[10\]
+ cpuregs.regs\[27\]\[10\] _04281_ _04470_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_126_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09669__A1 _04105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13174__S _07104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11476__A1 _06054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _04053_ _04403_ _04095_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15206__A3 _02058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08627_ _03386_ _03400_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__nor2_1
XANTENNA__16485__S _02968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15611__B1 _01959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08558_ irq_mask\[29\] irq_pending\[29\] VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__and2b_1
XFILLER_0_65_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16167__A1 net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08489_ is_lb_lh_lw_lbu_lhu _03270_ _03272_ _03249_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__and4_1
XANTENNA__12518__S _06737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09841__A1 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10987__B1 _05220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10520_ _03612_ _05220_ _05223_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__a21o_1
XANTENNA__12745__C _06082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14018__B _07778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_162_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10451_ cpuregs.regs\[28\]\[30\] cpuregs.regs\[29\]\[30\] cpuregs.regs\[30\]\[30\]
+ cpuregs.regs\[31\]\[30\] _04085_ _04087_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__mux4_1
XANTENNA__15390__A2 _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16514__A _02967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09827__S _04222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13170_ _06993_ cpuregs.regs\[4\]\[24\] _07104_ VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10382_ cpuregs.regs\[24\]\[28\] cpuregs.regs\[25\]\[28\] cpuregs.regs\[26\]\[28\]
+ cpuregs.regs\[27\]\[28\] _04216_ _04376_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12121_ _06516_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_984 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13689__C1 _07283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10562__A _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12052_ _06240_ cpuregs.regs\[22\]\[18\] _06471_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11164__B1 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14969__A _08335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11003_ _03471_ _05398_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__nor2_1
XANTENNA__13873__A _03301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16860_ _03151_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15525__S0 _01999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15811_ _05960_ _03634_ _03822_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__and3_1
X_16791_ _03137_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18530_ clknet_leaf_135_clk _01595_ VGND VGND VPWR VPWR cpuregs.regs\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15742_ timer\[22\] _02540_ _02543_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__o21ai_1
X_12954_ _06990_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18461_ clknet_leaf_184_clk _01526_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11905_ _06201_ cpuregs.regs\[20\]\[13\] _06398_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output110_A net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16395__S _02918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15673_ timer\[4\] _02490_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__or2_1
X_12885_ _06941_ cpuregs.regs\[31\]\[0\] _06943_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__mux2_1
XANTENNA_output208_A net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17412_ clknet_leaf_7_clk _00581_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_14624_ reg_next_pc\[25\] _07948_ _08264_ _08276_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__a22o_1
X_11836_ _06208_ cpuregs.regs\[11\]\[14\] _06359_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__mux2_1
X_18392_ clknet_leaf_3_clk _01457_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17343_ clknet_leaf_189_clk _00512_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14555_ _08212_ _07952_ VGND VGND VPWR VPWR _08213_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12428__S _06689_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11767_ _06313_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11332__S _03219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14209__A irq_state\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13506_ _04456_ decoded_imm\[9\] VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_140_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10718_ _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__inv_2
X_17274_ clknet_leaf_188_clk _00448_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14486_ decoded_imm_j\[15\] _07939_ VGND VGND VPWR VPWR _08149_ sky130_fd_sc_hd__or2_1
XANTENNA__15905__B2 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11698_ irq_state\[1\] VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16225_ net46 mem_16bit_buffer\[5\] _02831_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__mux2_1
X_13437_ _07296_ _07297_ _07298_ VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__nand3_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10649_ _04342_ _04419_ _03518_ _04456_ _05239_ _05237_ VGND VGND VPWR VPWR _05351_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12952__A _06273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13392__A1 _03276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16156_ net271 net233 _02786_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__mux2_1
X_13368_ _04036_ _04160_ _05257_ VGND VGND VPWR VPWR _07234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_155_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15107_ is_slli_srli_srai cpuregs.raddr2\[3\] decoded_imm\[3\] _01933_ _01934_ VGND
+ VGND VPWR VPWR _01964_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12319_ cpuregs.regs\[25\]\[31\] _06598_ _06603_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__mux2_1
X_16087_ is_slli_srli_srai _02650_ _02648_ _02657_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13299_ _07177_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09348__B1 _04082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15038_ irq_mask\[28\] _01865_ _01901_ _01891_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__a211o_1
XANTENNA__11287__B _05906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14892__A1 _05174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13783__A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14892__B2 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10902__A0 _05461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15516__S0 _01979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08877__A _00065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16989_ clknet_leaf_1_clk _00163_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__14644__A1 reg_next_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09530_ _04257_ _04260_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12655__A0 _06312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18728_ net121 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09520__A0 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09461_ _04153_ _04155_ _04152_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_64_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_184_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_184_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_149_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08412_ prefetched_high_word _03193_ _03197_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__and3_2
XFILLER_0_148_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09392_ _00071_ _04125_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09501__A _04091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12338__S _06641_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10433__A2 _04448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11630__A1 _06186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10984__A3 _04754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11069__S0 _05237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10197__A1 _04271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09682__S0 _04056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12073__S _06482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10292__S1 _04219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11146__B1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12894__A0 _06949_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12801__S _06891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15507__S0 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16085__A0 is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15427__A3 _02267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14635__A1 _03294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09728_ _04452_ _04453_ _04392_ _04395_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__o211ai_1
XANTENNA__10321__S _00071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09659_ _04383_ _04384_ _04387_ _03301_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__o211a_2
Xclkbuf_leaf_175_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_175_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__10672__A2 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12670_ _06096_ cpuregs.regs\[12\]\[1\] _06825_ VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15596__C1 _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09411__A _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _06183_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__buf_2
XANTENNA__18146__D alu_out\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12248__S _06533_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10557__A _05260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08617__A2 irq_active VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11152__S _04745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14340_ _03294_ _07911_ _07997_ _08014_ VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__a22o_1
X_11552_ reg_pc\[4\] _06110_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10503_ irq_pending\[31\] _04007_ _05204_ _05207_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11483_ irq_mask\[29\] _03428_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__or2_1
X_14271_ _05857_ _06278_ VGND VGND VPWR VPWR _07957_ sky130_fd_sc_hd__or2_1
XFILLER_0_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13374__A1 _07232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16010_ _02611_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__clkbuf_4
X_10434_ _04168_ _05139_ _05140_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__a21o_1
X_13222_ _07136_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09557__S _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10188__A1 _04320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09673__S0 _04056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13079__S _07057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10365_ count_cycle\[27\] _04165_ _05073_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__a21o_1
X_13153_ _06976_ cpuregs.regs\[4\]\[16\] _07093_ VGND VGND VPWR VPWR _07100_ sky130_fd_sc_hd__mux2_1
XANTENNA__10283__S1 _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12104_ _06175_ cpuregs.regs\[23\]\[10\] _06507_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__mux2_1
XANTENNA__14323__B1 _07904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17961_ clknet_leaf_191_clk _01098_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dfxtp_1
X_13084_ _07063_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__clkbuf_1
X_10296_ _05005_ _05006_ _04321_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12035_ _06459_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__clkbuf_8
X_16912_ clknet_leaf_34_clk _00057_ VGND VGND VPWR VPWR mem_rdata_q\[31\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__12885__A0 _06941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17892_ clknet_leaf_92_clk _01061_ VGND VGND VPWR VPWR count_cycle\[37\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16843_ _03165_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15823__A0 decoded_imm_j\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16774_ _06557_ cpuregs.regs\[13\]\[11\] _03127_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__mux2_1
X_13986_ _07756_ _07757_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__nor2_1
X_18513_ clknet_leaf_116_clk _01578_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_15725_ _02477_ _02529_ _02530_ _02531_ _06026_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__o311a_1
XFILLER_0_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12937_ _06978_ cpuregs.regs\[31\]\[17\] _06964_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_166_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_166_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_103_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18444_ clknet_leaf_164_clk _01509_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15656_ _07208_ _02479_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _06297_ cpuregs.regs\[6\]\[25\] _06928_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09321__A _04055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _03195_ _03363_ _07959_ _07898_ VGND VGND VPWR VPWR _08261_ sky130_fd_sc_hd__o211a_1
X_18375_ clknet_leaf_154_clk _01440_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_11819_ _06141_ cpuregs.regs\[11\]\[6\] _06348_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15587_ cpuregs.regs\[8\]\[29\] cpuregs.regs\[9\]\[29\] cpuregs.regs\[10\]\[29\]
+ cpuregs.regs\[11\]\[29\] _03641_ _03684_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__mux4_1
XANTENNA__13601__A2 _05259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12799_ cpuregs.regs\[9\]\[25\] _06586_ _06891_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17326_ clknet_leaf_97_clk _00500_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14538_ decoded_imm_j\[19\] _07950_ VGND VGND VPWR VPWR _08197_ sky130_fd_sc_hd__or2_1
XANTENNA__09900__S1 _04218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11997__S _06446_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17257_ clknet_leaf_135_clk _00431_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_14469_ _07998_ _08119_ _07996_ VGND VGND VPWR VPWR _08134_ sky130_fd_sc_hd__o21a_1
XFILLER_0_141_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13365__A1 _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16208_ _06082_ _06862_ _02826_ decoded_rd\[3\] VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17188_ clknet_leaf_159_clk _00362_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16139_ _02787_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08961_ _03656_ _03723_ _03675_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12876__A0 _06328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09967__S1 _04470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08892_ _03656_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__buf_4
XANTENNA__14402__A decoded_imm_j\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10351__A1 _04215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14121__B _07815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15814__B1 _03977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09513_ reg_pc\[4\] decoded_imm\[4\] VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_157_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_157_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_148_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09444_ cpuregs.regs\[4\]\[3\] cpuregs.regs\[5\]\[3\] cpuregs.regs\[6\]\[3\] cpuregs.regs\[7\]\[3\]
+ _04084_ _04086_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__mux4_1
XFILLER_0_91_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_166_Right_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09375_ net64 net50 _04040_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__mux2_1
XANTENNA__16763__S _03116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09885__B decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14553__B1 _07904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_104_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10543__C _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09980__B1 _04095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10150_ _04863_ _04864_ _04287_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10590__A1 _04198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput270 net270 VGND VGND VPWR VPWR mem_wdata[16] sky130_fd_sc_hd__buf_1
Xoutput281 net281 VGND VGND VPWR VPWR mem_wdata[26] sky130_fd_sc_hd__clkbuf_1
Xoutput292 net292 VGND VGND VPWR VPWR mem_wdata[7] sky130_fd_sc_hd__clkbuf_1
X_10081_ cpuregs.regs\[0\]\[19\] cpuregs.regs\[1\]\[19\] cpuregs.regs\[2\]\[19\] cpuregs.regs\[3\]\[19\]
+ _04512_ _04513_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__mux4_1
XANTENNA__12531__S _06752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09732__B1 _04458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14608__B2 _03378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13840_ _07659_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_113_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14966__B _03298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13771_ net87 decoded_imm\[28\] VGND VGND VPWR VPWR _07610_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_148_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_148_clk sky130_fd_sc_hd__clkbuf_2
X_10983_ _03574_ _05665_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_48_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15510_ cpuregs.regs\[16\]\[24\] cpuregs.regs\[17\]\[24\] cpuregs.regs\[18\]\[24\]
+ cpuregs.regs\[19\]\[24\] _01985_ _01986_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12722_ _06304_ cpuregs.regs\[12\]\[26\] _06847_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__mux2_1
X_16490_ _02977_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15441_ _03687_ _02280_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11390__B _03987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12653_ _06304_ cpuregs.regs\[30\]\[26\] _06810_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__mux2_1
XANTENNA__16673__S _03039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11604_ reg_out\[10\] alu_out_q\[10\] _06067_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__mux2_1
XANTENNA__09799__B1 _04225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18160_ clknet_leaf_23_clk _01231_ VGND VGND VPWR VPWR decoded_imm_j\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15372_ _01932_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__buf_4
XFILLER_0_26_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12584_ _06780_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_61_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17111_ clknet_leaf_177_clk _00285_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14323_ _07989_ _07997_ _07999_ _07904_ reg_next_pc\[1\] VGND VGND VPWR VPWR _08000_
+ sky130_fd_sc_hd__a32o_1
X_11535_ _06106_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__clkbuf_1
X_18091_ clknet_leaf_102_clk _01195_ VGND VGND VPWR VPWR timer\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15336__A2 _02009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_122_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13347__A1 _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17042_ clknet_leaf_111_clk _00216_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_14254_ latched_branch irq_state\[0\] latched_store VGND VGND VPWR VPWR _07945_ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11466_ _06041_ irq_pending\[21\] _06051_ net14 VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__a31o_1
X_13205_ _07127_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_927 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10417_ _05122_ _05123_ _04575_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__mux2_1
X_14185_ count_instr\[62\] _07893_ _07826_ VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10256__S1 _04276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11397_ _03635_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13136_ _06959_ cpuregs.regs\[4\]\[8\] _07082_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10348_ cpuregs.regs\[20\]\[27\] cpuregs.regs\[21\]\[27\] cpuregs.regs\[22\]\[27\]
+ cpuregs.regs\[23\]\[27\] _04207_ _04208_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__mux4_1
Xalphacore_310 VGND VGND VPWR VPWR alphacore_310/HI cpi_insn[8] sky130_fd_sc_hd__conb_1
XANTENNA__15195__S1 _02047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_321 VGND VGND VPWR VPWR alphacore_321/HI cpi_insn[19] sky130_fd_sc_hd__conb_1
Xalphacore_332 VGND VGND VPWR VPWR alphacore_332/HI cpi_insn[30] sky130_fd_sc_hd__conb_1
XANTENNA__12858__A0 _06257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_343 VGND VGND VPWR VPWR alphacore_343/HI trace_data[4] sky130_fd_sc_hd__conb_1
X_10279_ _03384_ _04988_ _04989_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__and3_1
X_17944_ clknet_leaf_70_clk _08385_ VGND VGND VPWR VPWR reg_out\[24\] sky130_fd_sc_hd__dfxtp_1
X_13067_ _07054_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12441__S _06700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_354 VGND VGND VPWR VPWR alphacore_354/HI trace_data[15] sky130_fd_sc_hd__conb_1
Xalphacore_365 VGND VGND VPWR VPWR alphacore_365/HI trace_data[26] sky130_fd_sc_hd__conb_1
XANTENNA__08526__A1 _03305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09316__A instr_retirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12018_ _06462_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15037__B _01863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17875_ clknet_leaf_88_clk _01044_ VGND VGND VPWR VPWR count_cycle\[20\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16848__S _03163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11530__B1 _03326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16826_ _03156_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16757_ _06540_ cpuregs.regs\[13\]\[3\] _03116_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__mux2_1
X_13969_ _07745_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_139_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_139_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__13272__S _07154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15708_ timer\[13\] _02516_ _02518_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10636__A2 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_727 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16688_ _03082_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15024__A1 _03303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16221__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15639_ decoder_trigger do_waitirq irq_state\[0\] VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__o21ba_1
X_18427_ clknet_leaf_181_clk _01492_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[6\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16583__S _03026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13586__A1 _04810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09160_ _03849_ _03209_ _03210_ _03850_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18358_ clknet_leaf_189_clk _01423_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17309_ clknet_leaf_2_clk _00483_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09091_ _03849_ _03801_ _03802_ _03850_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18289_ clknet_leaf_37_clk _01357_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11364__A3 _03874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09993_ _03638_ _04708_ _04202_ irq_pending\[16\] _04712_ VGND VGND VPWR VPWR _04713_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__11756__A _06303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12351__S _06652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08944_ cpuregs.regs\[8\]\[4\] cpuregs.regs\[9\]\[4\] cpuregs.regs\[10\]\[4\] cpuregs.regs\[11\]\[4\]
+ _03649_ _03643_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__mux4_1
XANTENNA__10660__A _05225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11475__B _03428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08875_ _00064_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_4_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11521__B1 _06093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13971__A _07737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15263__A1 _02111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13182__S _07081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11491__A latched_branch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10088__B1 _04100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09427_ net34 net51 _04039_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__mux2_1
XANTENNA__15566__A2 _01905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09358_ cpuregs.regs\[8\]\[1\] cpuregs.regs\[9\]\[1\] cpuregs.regs\[10\]\[1\] cpuregs.regs\[11\]\[1\]
+ _04056_ _04091_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_43_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09245__A2 _03867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11588__B1 _06065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16515__A1 _06575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09289_ _04025_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11320_ _05076_ _05939_ _03219_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__mux2_1
XANTENNA__14526__B1 _07905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11251_ _04611_ _03841_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10202_ irq_pending\[22\] _04006_ _04912_ _04915_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__o22a_1
XANTENNA__09953__B1 _04673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11182_ _03219_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11760__B1 reg_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10133_ net45 _04745_ _04666_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11666__A _06223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12261__S _06604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15990_ _03636_ _03822_ _02702_ _02705_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__a31o_1
XANTENNA__13501__A1 _07274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10064_ _04156_ _04750_ _04751_ _04781_ VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__o31ai_1
X_14941_ _01845_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09181__A1 _03891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17660_ clknet_leaf_49_clk _00829_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dfxtp_4
X_14872_ count_cycle\[57\] count_cycle\[58\] _01795_ count_cycle\[59\] VGND VGND VPWR
+ VPWR _01802_ sky130_fd_sc_hd__a31o_1
XANTENNA__08975__A _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09570__S _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16611_ cpuregs.regs\[1\]\[1\] _06095_ _03040_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__mux2_1
X_13823_ cpuregs.regs\[0\]\[8\] VGND VGND VPWR VPWR _07651_ sky130_fd_sc_hd__clkbuf_1
X_17591_ clknet_leaf_121_clk _00760_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10079__B1 _04225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16542_ _03005_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__clkbuf_1
X_13754_ _04945_ _05261_ _07593_ _07274_ VGND VGND VPWR VPWR _07594_ sky130_fd_sc_hd__o211a_1
X_10966_ _05361_ _05643_ _05650_ VGND VGND VPWR VPWR alu_out\[19\] sky130_fd_sc_hd__a21o_1
XFILLER_0_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12705_ _06240_ cpuregs.regs\[12\]\[18\] _06836_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16473_ cpuregs.regs\[17\]\[0\] _06531_ _02968_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__mux2_1
X_13685_ _05044_ _07277_ VGND VGND VPWR VPWR _07530_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10897_ _05372_ _05379_ _05295_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__mux2_1
X_18212_ clknet_leaf_41_clk _01283_ VGND VGND VPWR VPWR instr_srl sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15424_ _02263_ _02264_ _03713_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__mux2_1
XANTENNA__14765__B1 _01723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12636_ _06240_ cpuregs.regs\[30\]\[18\] _06799_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_130_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18143_ clknet_leaf_46_clk alu_out\[17\] VGND VGND VPWR VPWR alu_out_q\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15355_ cpuregs.regs\[20\]\[16\] cpuregs.regs\[21\]\[16\] cpuregs.regs\[22\]\[16\]
+ cpuregs.regs\[23\]\[16\] _01970_ _01971_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12567_ _06771_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__clkbuf_1
X_14306_ _07977_ _07978_ _07982_ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__or3_2
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18074_ clknet_leaf_48_clk _01179_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11518_ latched_compr reg_pc\[1\] VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__or2b_1
X_15286_ net101 _02081_ _02133_ _02134_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__o22a_1
X_12498_ _06734_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17025_ clknet_leaf_183_clk _00199_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_150_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14237_ _05857_ _06198_ VGND VGND VPWR VPWR _07933_ sky130_fd_sc_hd__or2_1
X_11449_ irq_mask\[13\] _06042_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_78_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14168_ count_instr\[56\] _07881_ _07883_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__o21a_1
XANTENNA__11751__B1 _06093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15048__A _03670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13119_ _07081_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_111_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12171__S _06534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14099_ _07833_ _07835_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15493__A1 _03639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17927_ clknet_leaf_55_clk _08398_ VGND VGND VPWR VPWR reg_out\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16578__S _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09172__A1 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08660_ _03426_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__inv_2
X_17858_ clknet_leaf_93_clk _01027_ VGND VGND VPWR VPWR count_cycle\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16442__A0 _06980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09480__S _04211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16809_ _06592_ cpuregs.regs\[13\]\[28\] _03138_ VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__mux2_1
XANTENNA__13256__A0 _06941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08591_ _03248_ _03369_ _03367_ _03249_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__o211a_1
X_17789_ clknet_leaf_84_clk _00958_ VGND VGND VPWR VPWR count_instr\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15340__S1 _01977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13559__A1 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09212_ mem_rdata_q\[25\] _03954_ _03757_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__mux2_1
XANTENNA__14756__B1 _01723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14220__A2 _07906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11034__A2 _04945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09143_ _03861_ _03890_ _03899_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10655__A _05356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09074_ _03748_ _03789_ _03817_ _03834_ _03835_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__o221a_1
XANTENNA__14508__B1 _08050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08450__A3 _03199_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13731__A1 _05143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09976_ _04694_ _04695_ _04369_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__mux2_1
XANTENNA__16681__A0 _06947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08927_ _03689_ _03690_ _03664_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08858_ _03623_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08789_ _03504_ _03554_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__nor2_1
XANTENNA__15331__S1 _02000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10820_ _05292_ _05336_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__nor2_1
XANTENNA__14995__B1 _01714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10549__B _05225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10751_ _05434_ _05439_ _05446_ _05448_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__o211a_1
XANTENNA__09871__C1 _04027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13470_ _07325_ _07326_ _07328_ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__o21bai_1
X_10682_ _05232_ _05317_ _05316_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14211__A2 _07906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12421_ _06693_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__18154__D alu_out\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10459__S1 _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11160__S _04668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18732__A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15140_ _03669_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__buf_6
XFILLER_0_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12352_ _06656_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11303_ _03841_ _05924_ _05925_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15172__B1 _02006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15071_ is_slli_srli_srai VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12283_ _06619_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_95_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13722__A1 _03276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14022_ _07781_ _07782_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__nor2_1
XANTENNA__13595__B decoded_imm\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11234_ _04532_ _05869_ _05827_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08689__B net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13087__S _07057_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ net115 _04710_ _05817_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_56_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15475__A1 _01969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ _04830_ _04831_ _04287_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__mux2_1
X_11096_ _03592_ _05086_ _05390_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__a21o_1
X_15973_ mem_rdata_q\[26\] _02690_ _02691_ _02650_ _04022_ VGND VGND VPWR VPWR _01295_
+ sky130_fd_sc_hd__a32o_2
XANTENNA_output238_A net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15570__S1 _01977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09154__A1 _03895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17712_ clknet_leaf_83_clk _00881_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10047_ cpuregs.regs\[24\]\[18\] cpuregs.regs\[25\]\[18\] cpuregs.regs\[26\]\[18\]
+ cpuregs.regs\[27\]\[18\] _04472_ _04473_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__mux4_1
X_14924_ net197 net166 _01835_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__mux2_1
XANTENNA__15227__A1 _01969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17643_ clknet_leaf_47_clk _00812_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfxtp_4
X_14855_ _01789_ _01753_ _01790_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__and3b_1
XFILLER_0_89_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15778__A2 _02486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15322__S1 _01980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13789__A1 _05086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13806_ _07642_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13333__S0 _04758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17574_ clknet_leaf_19_clk _00743_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_14786_ count_cycle\[31\] _01741_ _01717_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09457__A2 _04186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11998_ _06451_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__clkbuf_1
X_16525_ cpuregs.regs\[17\]\[25\] _06586_ _02990_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__mux2_1
X_13737_ net85 decoded_imm\[26\] VGND VGND VPWR VPWR _07578_ sky130_fd_sc_hd__nand2_1
X_10949_ _05634_ _05572_ _05331_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12955__A _06280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_128_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16456_ _02959_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__clkbuf_1
X_13668_ _07499_ _07508_ _07513_ _03311_ VGND VGND VPWR VPWR _07514_ sky130_fd_sc_hd__a31o_1
XFILLER_0_156_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15407_ _02004_ _02244_ _02248_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__a21o_1
X_12619_ _06787_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__buf_6
X_16387_ _06993_ cpuregs.regs\[16\]\[24\] _02918_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__mux2_1
XANTENNA__16861__S _03174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13599_ _07433_ _07448_ _07447_ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18126_ clknet_leaf_42_clk alu_out\[0\] VGND VGND VPWR VPWR alu_out_q\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15338_ cpuregs.regs\[12\]\[15\] cpuregs.regs\[13\]\[15\] cpuregs.regs\[14\]\[15\]
+ cpuregs.regs\[15\]\[15\] _01979_ _01980_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__mux4_1
XANTENNA__13961__B2 net148 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15389__S1 _02037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11972__A0 _06193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18057_ clknet_leaf_71_clk _01162_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dfxtp_4
XANTENNA__13786__A _05086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15269_ decoded_imm\[10\] _02009_ _01963_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__a21o_1
XANTENNA__09983__B _04702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10870__S1 _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17008_ clknet_leaf_164_clk _00182_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08599__B _03293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09393__A1 _04121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09830_ cpuregs.regs\[28\]\[12\] cpuregs.regs\[29\]\[12\] cpuregs.regs\[30\]\[12\]
+ cpuregs.regs\[31\]\[12\] _04329_ _04376_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__mux4_1
X_09761_ _04055_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__buf_6
XFILLER_0_77_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15561__S1 _02075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08712_ _03476_ _03477_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__or2b_1
XANTENNA__15506__A _01984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09692_ latched_is_lb _04363_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__and2_1
XANTENNA__10386__S0 _04273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08643_ cpu_state\[0\] _03274_ _03410_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__nor3_2
XANTENNA__15313__S1 _02014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08574_ irq_mask\[14\] irq_pending\[14\] VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__and2b_2
XFILLER_0_95_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_61_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10463__B1 net300 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13401__A0 _04160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10385__A _04328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09126_ _03854_ _03863_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__and2b_1
XFILLER_0_150_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_802 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10766__B2 _05461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09057_ mem_rdata_q\[23\] net48 _03208_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13704__A1 _04945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14901__A0 net214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09384__A1 _03384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10324__S _04063_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09959_ reg_pc\[15\] decoded_imm\[15\] decoded_imm\[14\] reg_pc\[14\] VGND VGND VPWR
+ VPWR _04679_ sky130_fd_sc_hd__o211a_1
XANTENNA__15552__S1 _02031_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11944__A cpuregs.waddr\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12970_ _06319_ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_51_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11921_ _06410_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__18149__D alu_out\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15304__S1 _02014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__18727__A net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14640_ _08287_ _08289_ VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__and2_1
X_11852_ _06372_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15090__C1 _00067_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14974__B _01865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10803_ _05486_ _05491_ _05497_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__or3_2
XFILLER_0_95_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12443__A1 _06584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14571_ _08226_ _08227_ VGND VGND VPWR VPWR _08228_ sky130_fd_sc_hd__nand2_1
X_11783_ _06327_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__buf_2
XFILLER_0_68_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_52_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16310_ _06984_ cpuregs.regs\[15\]\[20\] _02881_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__mux2_1
X_13522_ _07376_ _07377_ VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__nand2_1
XANTENNA__10454__B1 _04082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15151__A _02005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10734_ _03522_ _05431_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__nor2_1
X_17290_ clknet_leaf_144_clk _00464_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16241_ net54 mem_16bit_buffer\[13\] _02830_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13453_ _07297_ _07312_ _07309_ _03631_ VGND VGND VPWR VPWR _07314_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_97_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10665_ _03608_ _05364_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__nand2_1
XANTENNA__16681__S _03076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14990__A _04382_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12404_ _06684_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__clkbuf_1
X_16172_ _02804_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__clkbuf_1
X_13384_ _07243_ _07244_ _07246_ VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10596_ _05288_ _05291_ _05297_ _05298_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15123_ cpuregs.regs\[20\]\[5\] cpuregs.regs\[21\]\[5\] cpuregs.regs\[22\]\[5\] cpuregs.regs\[23\]\[5\]
+ _01976_ _01977_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_58_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12335_ _06647_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12714__S _06847_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15054_ cpuregs.regs\[4\]\[0\] cpuregs.regs\[5\]\[0\] cpuregs.regs\[6\]\[0\] cpuregs.regs\[7\]\[0\]
+ _03658_ _03659_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__mux4_1
X_12266_ _06610_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09375__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14005_ _07769_ _07770_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__nor2_1
X_11217_ _05855_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09308__B decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput70 net70 VGND VGND VPWR VPWR cpi_rs1[12] sky130_fd_sc_hd__buf_1
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12197_ _06564_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__clkbuf_1
Xoutput81 net81 VGND VGND VPWR VPWR cpi_rs1[22] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_71_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput92 net92 VGND VGND VPWR VPWR cpi_rs1[3] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11148_ _05324_ net106 _04745_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__mux2_1
XANTENNA__15543__S1 _03642_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11079_ _03449_ _05755_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__xnor2_1
X_15956_ mem_state\[1\] VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__inv_2
XANTENNA__08866__C _03305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09324__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14907_ net219 net188 _01824_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__mux2_1
X_15887_ _02612_ mem_rdata_q\[14\] _02613_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__or3b_1
XANTENNA__16856__S _03163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14959__A0 net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17626_ clknet_leaf_106_clk _00795_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_14838_ _01779_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14423__A2 _07948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15620__B2 _03675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14769_ count_cycle\[25\] count_cycle\[26\] _01729_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__and3_1
X_17557_ clknet_leaf_100_clk _00726_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_43_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_85_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10445__B1 _04017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16508_ cpuregs.regs\[17\]\[17\] _06569_ _02979_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17488_ clknet_leaf_116_clk _00657_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16439_ _02950_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__16591__S _03026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15923__A2 _02617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13934__A1 _03348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18109_ clknet_leaf_81_clk _01213_ VGND VGND VPWR VPWR timer\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10933__A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12624__S _06799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15231__S0 _01970_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08403__A latched_branch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11173__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15439__A1 _02111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09813_ _04535_ _04536_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__nand2_1
XANTENNA__15534__S1 _01937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09744_ _04469_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11483__B _03428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09675_ _04401_ _04402_ _00071_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08626_ _03399_ _03315_ _03312_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_96_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14794__B _08350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15611__A1 decoded_imm\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15611__B2 _02440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08557_ irq_mask\[18\] irq_pending\[18\] VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__and2b_2
XANTENNA__08792__B net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13190__S _07118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__16067__A _02610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_611 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08488_ _03239_ _03271_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__nor2_4
XANTENNA__09841__A2 _04544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13925__A1 _03353_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10450_ _04483_ _05155_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10739__A1 _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11936__A0 _06320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09109_ _03866_ _03868_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__and2b_2
XFILLER_0_161_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10381_ _04105_ count_cycle\[60\] _03253_ count_cycle\[28\] _05088_ VGND VGND VPWR
+ VPWR _05089_ sky130_fd_sc_hd__a221o_1
XANTENNA__11400__A2 _03916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16875__A0 _06590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15678__A1 _01872_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12120_ _06240_ cpuregs.regs\[23\]\[18\] _06507_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__mux2_1
XANTENNA__09409__A _04051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13689__B1 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12051_ _06479_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11164__A1 _03407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11164__B2 _03297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11002_ _05683_ _05634_ _05395_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__mux2_1
XANTENNA__15525__S1 _02000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15810_ decoded_imm_j\[5\] _05983_ _03954_ _02587_ _02588_ VGND VGND VPWR VPWR _01235_
+ sky130_fd_sc_hd__a221o_1
X_16790_ _06573_ cpuregs.regs\[13\]\[19\] _03127_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__mux2_1
X_15741_ timer\[22\] _02540_ _02488_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12953_ _06989_ cpuregs.regs\[31\]\[22\] _06985_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14985__A _04227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10675__A0 _04198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15289__S0 _01976_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11904_ _06401_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__clkbuf_1
X_18460_ clknet_leaf_173_clk _01525_ VGND VGND VPWR VPWR cpuregs.regs\[17\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15672_ _04185_ _02477_ _02492_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__a21oi_1
X_12884_ _06942_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__buf_6
XANTENNA__15063__C1 _03654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17411_ clknet_leaf_11_clk _00580_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14623_ _08012_ _08274_ _08275_ _07962_ VGND VGND VPWR VPWR _08276_ sky130_fd_sc_hd__o2bb2a_1
X_11835_ _06363_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__clkbuf_1
X_18391_ clknet_leaf_12_clk _01456_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output103_A net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_25 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_16_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11613__S _06176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17342_ clknet_leaf_18_clk _00511_ VGND VGND VPWR VPWR cpuregs.regs\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ decoded_imm_j\[20\] VGND VGND VPWR VPWR _08212_ sky130_fd_sc_hd__buf_2
XFILLER_0_138_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11766_ _06312_ cpuregs.regs\[10\]\[27\] _06258_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__mux2_1
XANTENNA__10978__A1 _05225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13505_ _07362_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10717_ _03524_ net93 net92 net89 _03609_ _05231_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__mux4_2
XFILLER_0_125_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15366__B1 _01968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17273_ clknet_leaf_17_clk _00447_ VGND VGND VPWR VPWR cpuregs.regs\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14485_ decoded_imm_j\[15\] _07939_ VGND VGND VPWR VPWR _08148_ sky130_fd_sc_hd__nand2_1
X_11697_ reg_pc\[20\] _06242_ _06250_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__o21a_1
XANTENNA__15905__A2 _02635_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16224_ _02836_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__clkbuf_1
X_13436_ _04262_ decoded_imm\[5\] VGND VGND VPWR VPWR _07298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09045__A0 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10648_ _04160_ _04251_ _04198_ _03524_ _05239_ _05237_ VGND VGND VPWR VPWR _05350_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16155_ _02795_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__clkbuf_1
X_13367_ _03387_ _04101_ _07210_ reg_pc\[1\] VGND VGND VPWR VPWR _07233_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_3_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10579_ _03242_ _04036_ _03609_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15213__S0 _01982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15106_ _01934_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__buf_6
XANTENNA__09319__A _04053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12318_ _06637_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__clkbuf_1
X_16086_ _02753_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13298_ _06984_ cpuregs.regs\[5\]\[20\] _07176_ VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09348__A1 _04070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15037_ _05106_ _01863_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__nor2_1
X_12249_ _06599_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11287__C _05911_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13783__B decoded_imm\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15516__S1 _01980_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16988_ clknet_leaf_3_clk _00162_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[3\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14644__A2 _07948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18727_ net110 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_160_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15939_ mem_rdata_q\[21\] mem_rdata_q\[22\] mem_rdata_q\[23\] _02664_ VGND VGND VPWR
+ VPWR _02665_ sky130_fd_sc_hd__nor4_4
XFILLER_0_64_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09520__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09989__A _03225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09460_ reg_pc\[3\] decoded_imm\[3\] VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__or2_1
XANTENNA__08954__S0 _03649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10130__A2 _04012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08893__A _00064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08411_ prefetched_high_word clear_prefetched_high_word_q _03195_ latched_branch
+ _03196_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_121_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17609_ clknet_leaf_186_clk _00778_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_09391_ cpuregs.regs\[16\]\[2\] cpuregs.regs\[17\]\[2\] cpuregs.regs\[18\]\[2\] cpuregs.regs\[19\]\[2\]
+ _04123_ _04124_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__mux4_1
XFILLER_0_171_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13604__B1 _07210_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18589_ clknet_leaf_180_clk _01654_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_814 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11091__B1 _05251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13907__A1 _03323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09928__S _04121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15109__B1 _01965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11759__A reg_pc\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10197__A2 _04909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09682__S1 _04091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09027__A_N _03206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13974__A _07737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14332__A1 _07901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11146__A1 _03407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11146__B2 _04422_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15507__S1 _02014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08787__B net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14301__C irq_pending\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14635__A2 _07966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09727_ _04392_ _04395_ _04452_ _04453_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__a211o_1
XANTENNA__16496__S _02979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09511__A1 _04168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10657__B1 _05301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09899__A _04328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08945__S0 _03649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09658_ count_cycle\[7\] _04013_ _04386_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08609_ cpu_state\[3\] VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14399__A1 _07899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15596__B1 _01959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10672__A3 _04342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09589_ cpuregs.regs\[24\]\[6\] cpuregs.regs\[25\]\[6\] cpuregs.regs\[26\]\[6\] cpuregs.regs\[27\]\[6\]
+ _04274_ _04317_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11620_ _06075_ _06178_ _06179_ _06182_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__a31o_2
XFILLER_0_38_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ reg_pc\[4\] _06110_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10502_ _03680_ _05205_ _04752_ _05206_ _04202_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__a221o_1
X_14270_ reg_pc\[22\] _07953_ _07956_ _07935_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11482_ _06054_ irq_pending\[28\] _06060_ net21 VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11909__A0 _06216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13221_ _06976_ cpuregs.regs\[8\]\[16\] _07129_ VGND VGND VPWR VPWR _07136_ sky130_fd_sc_hd__mux2_1
X_10433_ irq_mask\[29\] _04448_ timer\[29\] _04187_ _04188_ VGND VGND VPWR VPWR _05140_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__09578__B2 _04023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09673__S1 _04091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13152_ _07099_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10364_ count_instr\[27\] _04011_ _04009_ _05072_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12103_ _06495_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17960_ clknet_leaf_191_clk _01097_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dfxtp_1
X_13083_ _06974_ cpuregs.regs\[7\]\[15\] _07057_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__mux2_1
XANTENNA__14323__B2 reg_next_pc\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10295_ cpuregs.regs\[8\]\[25\] cpuregs.regs\[9\]\[25\] cpuregs.regs\[10\]\[25\]
+ cpuregs.regs\[11\]\[25\] _04325_ _04277_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__mux4_1
XANTENNA__09573__S _04223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12034_ _06470_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__clkbuf_1
X_16911_ clknet_leaf_34_clk _00056_ VGND VGND VPWR VPWR mem_rdata_q\[30\] sky130_fd_sc_hd__dfxtp_2
X_17891_ clknet_leaf_92_clk _01060_ VGND VGND VPWR VPWR count_cycle\[36\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16076__A1 decoded_imm\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16076__B2 mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16842_ _06557_ cpuregs.regs\[14\]\[11\] _03163_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__mux2_1
XANTENNA__14087__B1 _07826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15284__C1 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15823__A1 _03737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output220_A net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16773_ _03128_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__clkbuf_1
X_13985_ count_instr\[0\] _07755_ _06054_ VGND VGND VPWR VPWR _07757_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10648__A0 _04160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18512_ clknet_leaf_108_clk _01577_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_15724_ _04737_ _02479_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__nand2_1
X_12936_ _06231_ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__buf_2
XFILLER_0_88_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18443_ clknet_leaf_122_clk _01508_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_15655_ _02475_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__clkbuf_4
X_12867_ _06933_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12439__S _06700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11343__S _03219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _06354_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_83_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _08257_ _08246_ _08259_ VGND VGND VPWR VPWR _08260_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18374_ clknet_leaf_139_clk _01439_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_15586_ cpuregs.regs\[12\]\[29\] cpuregs.regs\[13\]\[29\] cpuregs.regs\[14\]\[29\]
+ cpuregs.regs\[15\]\[29\] _03641_ _03684_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__mux4_1
X_12798_ _06896_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09805__A2 _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ clknet_leaf_98_clk _00499_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14537_ decoded_imm_j\[19\] _07950_ VGND VGND VPWR VPWR _08196_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11749_ _06297_ cpuregs.regs\[10\]\[25\] _06258_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15434__S0 _02111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17256_ clknet_leaf_132_clk _00430_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14468_ _08131_ _08132_ _08012_ VGND VGND VPWR VPWR _08133_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13419_ _07211_ VGND VGND VPWR VPWR _07282_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13365__A2 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16207_ _04156_ _07898_ _06863_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__and3_1
X_17187_ clknet_leaf_133_clk _00361_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12174__S _06534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14399_ _07899_ _07921_ _07992_ _08069_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__a31o_1
XFILLER_0_113_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16138_ net293 net255 _02786_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08960_ _03721_ _03722_ _03713_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__mux2_1
X_16069_ decoded_imm\[20\] _02650_ _02746_ mem_rdata_q\[20\] _02749_ VGND VGND VPWR
+ VPWR _01333_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_5_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__10336__C1 _04202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08891_ _00067_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__inv_2
XANTENNA__09741__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09741__B2 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15814__A1 decoded_imm_j\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09512_ _04010_ _04205_ _04243_ _04150_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__o211a_1
XANTENNA__10103__A2 decoded_imm\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11761__B _06118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09443_ _04069_ _04175_ _04081_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12349__S _06652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15042__A2 _01865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09374_ _04102_ _04103_ _04108_ _03303_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09009__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16064__B _02610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14553__A1 _07898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14553__B2 reg_next_pc\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08783__A2 _03518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09980__A1 _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput260 net260 VGND VGND VPWR VPWR mem_la_wstrb[2] sky130_fd_sc_hd__clkbuf_1
XANTENNA__11119__B2 _05254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10590__A2 _04160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput271 net271 VGND VGND VPWR VPWR mem_wdata[17] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput282 net282 VGND VGND VPWR VPWR mem_wdata[27] sky130_fd_sc_hd__clkbuf_1
X_10080_ cpuregs.regs\[4\]\[19\] cpuregs.regs\[5\]\[19\] cpuregs.regs\[6\]\[19\] cpuregs.regs\[7\]\[19\]
+ _04512_ _04513_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__mux4_1
Xoutput293 net293 VGND VGND VPWR VPWR mem_wdata[8] sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09732__B2 _03225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14608__A2 _07904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13770_ net87 decoded_imm\[28\] VGND VGND VPWR VPWR _07609_ sky130_fd_sc_hd__and2_1
X_10982_ _05517_ _03464_ _05662_ _05664_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__o31a_1
XFILLER_0_69_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12721_ _06853_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_154_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__18157__D alu_out\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12259__S _06604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15440_ cpuregs.regs\[24\]\[20\] cpuregs.regs\[25\]\[20\] cpuregs.regs\[26\]\[20\]
+ cpuregs.regs\[27\]\[20\] _01996_ _01997_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__mux4_1
X_12652_ _06816_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09248__A0 mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11055__B1 _05221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11603_ _06167_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09799__A1 _04289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15371_ _02202_ _02206_ _02027_ _02214_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__o211a_4
XFILLER_0_38_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12583_ cpuregs.regs\[2\]\[25\] _06586_ _06774_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15416__S0 _02046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_169_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17110_ clknet_leaf_127_clk _00284_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14322_ compressed_instr decoded_imm_j\[1\] _07998_ VGND VGND VPWR VPWR _07999_ sky130_fd_sc_hd__mux2_1
X_11534_ _06105_ cpuregs.regs\[10\]\[2\] _06086_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__mux2_1
X_18090_ clknet_leaf_100_clk _01194_ VGND VGND VPWR VPWR timer\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17041_ clknet_leaf_160_clk _00215_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13347__A2 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14253_ _07942_ VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__buf_4
XFILLER_0_162_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15741__B1 _02488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11465_ irq_mask\[21\] _06042_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13204_ _06959_ cpuregs.regs\[8\]\[8\] _07118_ VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10416_ cpuregs.regs\[24\]\[29\] cpuregs.regs\[25\]\[29\] cpuregs.regs\[26\]\[29\]
+ cpuregs.regs\[27\]\[29\] _04579_ _04284_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__mux4_1
X_14184_ _07893_ _07894_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11396_ cpuregs.raddr1\[0\] _03636_ _06005_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13135_ _07090_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12722__S _06847_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10347_ _04272_ _05055_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14503__A decoded_imm_j\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_311 VGND VGND VPWR VPWR alphacore_311/HI cpi_insn[9] sky130_fd_sc_hd__conb_1
Xalphacore_322 VGND VGND VPWR VPWR alphacore_322/HI cpi_insn[20] sky130_fd_sc_hd__conb_1
XFILLER_0_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xalphacore_333 VGND VGND VPWR VPWR alphacore_333/HI cpi_insn[31] sky130_fd_sc_hd__conb_1
X_17943_ clknet_leaf_67_clk _08384_ VGND VGND VPWR VPWR reg_out\[23\] sky130_fd_sc_hd__dfxtp_1
X_13066_ _06957_ cpuregs.regs\[7\]\[7\] _07046_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__mux2_1
Xalphacore_344 VGND VGND VPWR VPWR alphacore_344/HI trace_data[5] sky130_fd_sc_hd__conb_1
X_10278_ _04984_ _04987_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__nand2_1
Xalphacore_355 VGND VGND VPWR VPWR alphacore_355/HI trace_data[16] sky130_fd_sc_hd__conb_1
XANTENNA__16049__A1 decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_366 VGND VGND VPWR VPWR alphacore_366/HI trace_data[27] sky130_fd_sc_hd__conb_1
XANTENNA__09723__A1 _04168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12017_ _06096_ cpuregs.regs\[22\]\[1\] _06460_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__mux2_1
XANTENNA__13119__A _07081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17874_ clknet_leaf_88_clk _01043_ VGND VGND VPWR VPWR count_cycle\[19\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11530__B2 _06072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16825_ _06540_ cpuregs.regs\[14\]\[3\] _03152_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12958__A _06288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16756_ _03119_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13968_ _07737_ _07744_ VGND VGND VPWR VPWR _07745_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10716__S0 _05413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14480__B1 _07994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09332__A _04054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10097__B2 _04813_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15707_ timer\[13\] _02516_ _02488_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12919_ _06966_ cpuregs.regs\[31\]\[11\] _06964_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__mux2_1
X_13899_ _07691_ _07696_ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__and2_1
X_16687_ _06953_ cpuregs.regs\[19\]\[5\] _03076_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__mux2_1
XANTENNA__15024__A2 _04022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18426_ clknet_leaf_166_clk _01491_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15638_ _02463_ _03307_ _02464_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14232__B1 _07901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11046__B1 _05218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18357_ clknet_leaf_17_clk _01422_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15569_ cpuregs.regs\[4\]\[28\] cpuregs.regs\[5\]\[28\] cpuregs.regs\[6\]\[28\] cpuregs.regs\[7\]\[28\]
+ _01973_ _01974_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_155_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17308_ clknet_leaf_12_clk _00482_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09090_ _03754_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08462__A1 irq_mask\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18288_ clknet_leaf_39_clk _01356_ VGND VGND VPWR VPWR mem_state\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14535__A1 reg_next_pc\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17239_ clknet_leaf_155_clk _00413_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_116_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10417__S _04575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11349__A1 _03891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11349__B2 _03736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_6_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10021__A1 _04168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09992_ _04709_ _04711_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__nor2_2
XANTENNA__12632__S _06799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08943_ reg_sh\[3\] reg_sh\[2\] reg_sh\[4\] VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__15867__A_N _02613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08874_ _00068_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_4_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13463__S _07225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16774__S _03127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09426_ net89 VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13026__A1 _06575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13699__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09357_ cpuregs.regs\[12\]\[1\] cpuregs.regs\[13\]\[1\] cpuregs.regs\[14\]\[1\] cpuregs.regs\[15\]\[1\]
+ _04056_ _04091_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_986 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12807__S _06891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09288_ instr_timer instr_maskirq instr_retirq VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__nor3_2
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14307__B _07983_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11250_ _05872_ _05877_ _05881_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10201_ _03637_ _04913_ _04673_ _04914_ _04266_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11181_ _03217_ _05825_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11760__A1 reg_pc\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10132_ net79 VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11158__S _04668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10063_ _04752_ _04753_ _04755_ _04780_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__a211oi_1
X_14940_ net205 net174 _01835_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__mux2_1
XANTENNA__09181__A2 _03747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14871_ count_cycle\[58\] count_cycle\[59\] _01798_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__and3_1
X_16610_ _03041_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15154__A _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13822_ _07650_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__clkbuf_1
X_17590_ clknet_leaf_98_clk _00759_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10079__A1 _04054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13753_ _05205_ _05227_ VGND VGND VPWR VPWR _07593_ sky130_fd_sc_hd__or2_1
X_16541_ _06941_ cpuregs.regs\[18\]\[0\] _03004_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10965_ _05385_ _05597_ _05601_ _05528_ _05649_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__a221o_1
XANTENNA__14993__A _04414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12704_ _06844_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__clkbuf_1
X_13684_ _07527_ _07528_ VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__nor2_1
X_16472_ _02967_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_80_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10896_ _03619_ _05583_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18211_ clknet_leaf_42_clk _01282_ VGND VGND VPWR VPWR instr_xor sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12635_ _06807_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__clkbuf_1
X_15423_ cpuregs.regs\[24\]\[19\] cpuregs.regs\[25\]\[19\] cpuregs.regs\[26\]\[19\]
+ cpuregs.regs\[27\]\[19\] _03640_ _03642_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15354_ net105 _02081_ _02196_ _02198_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__o22a_1
X_18142_ clknet_leaf_45_clk alu_out\[16\] VGND VGND VPWR VPWR alu_out_q\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12566_ cpuregs.regs\[2\]\[17\] _06569_ _06763_ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14305_ _07979_ _07980_ _07981_ VGND VGND VPWR VPWR _07982_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11517_ reg_pc\[1\] latched_compr VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__nand2b_1
X_18073_ clknet_leaf_74_clk _01178_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dfxtp_4
X_15285_ decoded_imm\[11\] _02009_ _01963_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__a21o_1
X_12497_ _06232_ cpuregs.regs\[28\]\[17\] _06726_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__mux2_1
XANTENNA_output95_A net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14236_ reg_pc\[12\] _07926_ _07932_ _07912_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__a22o_1
X_17024_ clknet_leaf_186_clk _00198_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11448_ _03412_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_150_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11200__A0 _04262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14167_ count_instr\[56\] _07881_ _07826_ VGND VGND VPWR VPWR _07883_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11379_ _03916_ _03777_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__nor2_1
XANTENNA__11751__A1 reg_pc\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13118_ _06383_ _06904_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_111_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ count_instr\[35\] _07831_ _07834_ VGND VGND VPWR VPWR _07835_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17926_ clknet_leaf_54_clk _08397_ VGND VGND VPWR VPWR reg_out\[6\] sky130_fd_sc_hd__dfxtp_1
X_13049_ _07044_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11503__A1 _06066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17857_ clknet_leaf_101_clk _01026_ VGND VGND VPWR VPWR count_cycle\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13283__S _07165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16808_ _03146_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__clkbuf_1
X_08590_ decoder_trigger do_waitirq instr_waitirq VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__o21ai_1
X_17788_ clknet_leaf_84_clk _00957_ VGND VGND VPWR VPWR count_instr\[59\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09555__S0 _04282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16739_ _07005_ cpuregs.regs\[19\]\[30\] _03075_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10001__A _03384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16607__B cpuregs.waddr\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09211_ _03753_ _03823_ _03824_ _03754_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__a22o_2
XFILLER_0_173_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18409_ clknet_leaf_99_clk _01474_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09142_ _03835_ _03897_ _03898_ _03855_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__a22o_1
XANTENNA__08435__A1 _03218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11034__A3 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14508__A1 _07972_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09073_ _03215_ _03738_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__nor2_2
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13192__A0 _06947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09975_ cpuregs.regs\[12\]\[16\] cpuregs.regs\[13\]\[16\] cpuregs.regs\[14\]\[16\]
+ cpuregs.regs\[15\]\[16\] _04232_ _04233_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_168_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16769__S _03116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08926_ cpuregs.regs\[0\]\[3\] cpuregs.regs\[1\]\[3\] cpuregs.regs\[2\]\[3\] cpuregs.regs\[3\]\[3\]
+ _03658_ _03659_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__mux4_1
XANTENNA__13495__A1 _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08857_ _03604_ _03516_ _03605_ _03622_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__and4b_1
XANTENNA__09794__S0 _04282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08795__B net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ _03508_ _03552_ _03553_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11258__A0 reg_next_pc\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10750_ _05298_ _05447_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__nand2_1
XANTENNA__08499__C_N cpu_state\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09409_ _04051_ _04142_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10681_ _05313_ _05315_ _05239_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12537__S _06752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14318__A _07992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12420_ cpuregs.regs\[27\]\[13\] _06561_ _06689_ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10233__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12351_ cpuregs.regs\[26\]\[13\] _06561_ _06652_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__mux2_1
XANTENNA__11430__B1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11302_ _05920_ _05923_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__and2_1
XANTENNA__15172__A1 _02020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15070_ _03388_ _01929_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__nor2_1
XANTENNA__13876__B instr_retirq VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12282_ cpuregs.regs\[25\]\[13\] _06561_ _06615_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13368__S _05257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14021_ count_instr\[11\] _07777_ _07759_ VGND VGND VPWR VPWR _07782_ sky130_fd_sc_hd__o21ai_1
X_11233_ _05865_ _05868_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15149__A _03675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16121__A0 net263 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11164_ _03407_ _05324_ net129 _03297_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16679__S _03076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14988__A _04335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ cpuregs.regs\[0\]\[20\] cpuregs.regs\[1\]\[20\] cpuregs.regs\[2\]\[20\] cpuregs.regs\[3\]\[20\]
+ _04275_ _04278_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_73_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11095_ _03442_ _03591_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__nor2_1
X_15972_ mem_rdata_q\[27\] _02645_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__nor2_1
XANTENNA__08986__A _03747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17711_ clknet_leaf_76_clk _00880_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dfxtp_1
X_10046_ cpuregs.regs\[28\]\[18\] cpuregs.regs\[29\]\[18\] cpuregs.regs\[30\]\[18\]
+ cpuregs.regs\[31\]\[18\] _04472_ _04473_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__mux4_1
X_14923_ _01836_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__clkbuf_1
X_17642_ clknet_leaf_46_clk _00811_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dfxtp_4
X_14854_ count_cycle\[52\] _01786_ count_cycle\[53\] VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13805_ _05174_ _07641_ _07224_ VGND VGND VPWR VPWR _07642_ sky130_fd_sc_hd__mux2_1
X_17573_ clknet_leaf_187_clk _00742_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13333__S1 _04759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14785_ _01743_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__clkbuf_1
X_11997_ _06289_ cpuregs.regs\[21\]\[24\] _06446_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16524_ _02995_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__clkbuf_1
X_13736_ _07577_ VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__clkbuf_1
X_10948_ _05633_ _05598_ _05240_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10472__A1 _04391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16455_ _06993_ cpuregs.regs\[29\]\[24\] _02954_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__mux2_1
X_10879_ _03493_ _05568_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__xor2_1
X_13667_ _07511_ _07512_ VGND VGND VPWR VPWR _07513_ sky130_fd_sc_hd__nand2_1
XANTENNA__12447__S _06700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15406_ _03692_ _02247_ _03657_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12618_ _06798_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__clkbuf_1
X_13598_ _07433_ _07447_ _07448_ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__nand3_1
XFILLER_0_143_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16386_ _02922_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__clkbuf_1
X_18125_ clknet_leaf_21_clk _01229_ VGND VGND VPWR VPWR latched_compr sky130_fd_sc_hd__dfxtp_2
X_15337_ net104 _02081_ _02181_ _02182_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__o22a_1
X_12549_ cpuregs.regs\[2\]\[9\] _06552_ _06752_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_959 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18056_ clknet_leaf_47_clk _01161_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dfxtp_4
XANTENNA__13786__B decoded_imm\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15268_ _02103_ _02107_ _02027_ _02117_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__o211a_4
XANTENNA__09917__A1 irq_pending\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17007_ clknet_leaf_124_clk _00181_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_14219_ reg_next_pc\[7\] _05834_ _07901_ _07920_ VGND VGND VPWR VPWR _07921_ sky130_fd_sc_hd__o211a_2
XFILLER_0_50_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15059__A _03671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15199_ cpuregs.regs\[16\]\[7\] cpuregs.regs\[17\]\[7\] cpuregs.regs\[18\]\[7\] cpuregs.regs\[19\]\[7\]
+ _03645_ _01991_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10083__S0 _04273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14898__A net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16589__S _03026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16663__A1 _06303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09760_ _04484_ _04485_ _04121_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__mux2_1
XANTENNA__13477__A1 _03275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08896__A _00064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08711_ net109 net77 VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__nand2_1
X_17909_ clknet_leaf_85_clk _01078_ VGND VGND VPWR VPWR count_cycle\[54\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11488__B1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09691_ _03510_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10386__S1 _04283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08642_ cpu_state\[2\] cpu_state\[4\] VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__or2_4
XFILLER_0_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08573_ irq_mask\[13\] irq_pending\[13\] VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__and2b_2
XANTENNA__14977__A1 irq_mask\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15522__A _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10666__A _05221_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12357__S _06652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13401__A1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09605__B1 _04100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09125_ _03862_ _03739_ _03882_ _03767_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__a22o_1
XANTENNA__13977__A _07737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10766__A2 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09056_ _03728_ _03732_ _03734_ _03735_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11497__A irq_state\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09908__A1 _04082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13188__S _07118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13704__A2 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12820__S _06906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09958_ _04597_ _04677_ _04676_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__a21o_1
X_08909_ _00068_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__clkinv_4
X_09889_ net72 VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_51_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _06257_ cpuregs.regs\[20\]\[20\] _06409_ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11851_ _06266_ cpuregs.regs\[11\]\[21\] _06370_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__mux2_1
XANTENNA__14968__B2 _04150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10802_ _05218_ _05496_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14570_ _08219_ _08225_ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__nand2_1
X_11782_ _06116_ reg_next_pc\[29\] _06324_ _06326_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__a211o_2
XFILLER_0_95_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10454__A1 _04231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10733_ _03546_ _05430_ _05363_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__mux2_1
X_13521_ net69 decoded_imm\[11\] VGND VGND VPWR VPWR _07377_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12267__S _06604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13452_ _07297_ _07309_ _07312_ VGND VGND VPWR VPWR _07313_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16240_ _02844_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10664_ _03608_ _05364_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_14_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12403_ cpuregs.regs\[27\]\[5\] _06544_ _06678_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13383_ _07247_ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16171_ net279 net241 _02797_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__mux2_1
X_10595_ _05228_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12334_ cpuregs.regs\[26\]\[5\] _06544_ _06641_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__mux2_1
X_15122_ _01919_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__buf_6
XFILLER_0_50_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13098__S _07068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15053_ _01907_ _01910_ _01912_ _03654_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12265_ cpuregs.regs\[25\]\[5\] _06544_ _06604_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14004_ count_instr\[6\] _07767_ _07759_ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__o21ai_1
X_11216_ _04419_ _05854_ _05827_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12196_ cpuregs.regs\[24\]\[14\] _06563_ _06555_ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__mux2_1
Xoutput71 net71 VGND VGND VPWR VPWR cpi_rs1[13] sky130_fd_sc_hd__clkbuf_1
Xoutput82 net82 VGND VGND VPWR VPWR cpi_rs1[23] sky130_fd_sc_hd__buf_1
Xoutput93 net93 VGND VGND VPWR VPWR cpi_rs1[4] sky130_fd_sc_hd__buf_1
X_11147_ _03407_ net128 net105 _04422_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__a22o_2
XFILLER_0_128_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14656__B1 _07997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09758__S0 _04232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11078_ _05323_ _03451_ _05752_ _05754_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__a31o_1
X_15955_ _02675_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__buf_2
X_10029_ _04150_ _04740_ _04743_ _04747_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__a31o_1
X_14906_ _01827_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08866__D _03631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15886_ instr_lh _02635_ _02637_ is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR _01262_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14959__A1 net184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17625_ clknet_leaf_114_clk _00794_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_14837_ _01777_ _01753_ _01778_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__and3b_1
XFILLER_0_53_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17556_ clknet_leaf_152_clk _00725_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13631__A1 _03275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14768_ count_cycle\[25\] _01729_ _01731_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__o21a_1
XANTENNA__09835__B1 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16507_ _02986_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__clkbuf_1
X_13719_ _07217_ _07519_ _07560_ _07561_ VGND VGND VPWR VPWR _07562_ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09930__S0 _04232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17487_ clknet_leaf_144_clk _00656_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12177__S _06534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14699_ _08340_ _08341_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16438_ _06976_ cpuregs.regs\[29\]\[16\] _02943_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13797__A _05174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15488__S _03653_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16369_ _02913_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10748__A2 _05440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18108_ clknet_leaf_81_clk _01212_ VGND VGND VPWR VPWR timer\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10933__B net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18039_ clknet_leaf_67_clk _00016_ VGND VGND VPWR VPWR irq_pending\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15231__S1 _01971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10425__S _04430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_986 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08403__B latched_store VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11110__A net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11173__A2 _04710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16636__A1 _06200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12370__A1 _06580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09812_ reg_pc\[12\] decoded_imm\[12\] VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10381__B1 _03253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14647__B1 _08055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09743_ _04058_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09523__C1 _04202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09674_ cpuregs.regs\[12\]\[8\] cpuregs.regs\[13\]\[8\] cpuregs.regs\[14\]\[8\] cpuregs.regs\[15\]\[8\]
+ _04056_ _04091_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_143_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08625_ reg_sh\[4\] reg_sh\[3\] reg_sh\[2\] VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__or3_4
XANTENNA__15072__B1 _03387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15252__A _01989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15611__A2 _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08556_ irq_mask\[11\] irq_pending\[11\] VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__and2b_2
XFILLER_0_76_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08629__B2 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13622__B2 reg_pc\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08487_ cpu_state\[2\] VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16782__S _03127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12087__S _06496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10987__A2 _05301_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16572__A0 _06974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13386__B1 _07211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15398__S _03653_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16083__A _03213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13500__A _04602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09396__S _00071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09108_ _03827_ _03867_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__or2b_1
XANTENNA__10295__S0 _04325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16324__A0 _06999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10380_ count_instr\[60\] _04015_ instr_rdinstr count_instr\[28\] VGND VGND VPWR
+ VPWR _05088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09039_ net59 mem_rdata_q\[4\] _03730_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__mux2_1
XANTENNA__15678__A2 _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13689__A1 _07304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09409__B _04142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10047__S0 _04472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12050_ _06232_ cpuregs.regs\[22\]\[17\] _06471_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11164__A2 _05324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11001_ _05682_ _05658_ _05232_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__mux2_1
XANTENNA__12361__A1 _06571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16627__A1 _06165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16088__C1 instr_jalr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15740_ _04871_ _02506_ _02542_ _02481_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__o211a_1
X_12952_ _06273_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__buf_2
XANTENNA__10124__B1 _04225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10675__A1 _04160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15289__S1 _01977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11903_ _06193_ cpuregs.regs\[20\]\[12\] _06398_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__mux2_1
X_15671_ _02484_ _02490_ _02491_ _03240_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__a31o_1
X_12883_ _06346_ _06713_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__nand2_4
X_17410_ clknet_leaf_188_clk _00579_ VGND VGND VPWR VPWR cpuregs.regs\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15162__A _02012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14622_ _07998_ _08258_ _07997_ VGND VGND VPWR VPWR _08275_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18390_ clknet_leaf_189_clk _01455_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11834_ _06201_ cpuregs.regs\[11\]\[13\] _06359_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17341_ clknet_leaf_16_clk _00088_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_83_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11765_ _06311_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__buf_2
X_14553_ _07898_ _07952_ _08050_ _07904_ reg_next_pc\[20\] VGND VGND VPWR VPWR _08211_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_166_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16012__C1 _02634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10716_ _05294_ _05289_ _05290_ _05306_ _05413_ _05414_ VGND VGND VPWR VPWR _05415_
+ sky130_fd_sc_hd__mux4_1
X_13504_ _04456_ _07361_ _07225_ VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__mux2_1
XANTENNA__15366__A1 _02012_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17272_ clknet_leaf_177_clk _00446_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_101_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11696_ reg_pc\[20\] _06242_ _06093_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__a21oi_1
X_14484_ reg_next_pc\[14\] _07948_ _08147_ _07960_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16223_ net45 mem_16bit_buffer\[4\] _02831_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__mux2_1
X_10647_ _05346_ _05348_ _05246_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__mux2_1
X_13435_ _03524_ decoded_imm\[5\] VGND VGND VPWR VPWR _07297_ sky130_fd_sc_hd__or2_2
XFILLER_0_67_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13366_ _07189_ VGND VGND VPWR VPWR _07232_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10286__S0 _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16154_ net270 net232 _02786_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10578_ _05251_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10060__C1 _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15105_ _05413_ _01906_ _01962_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__o21a_1
XANTENNA__15213__S1 _02004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12317_ cpuregs.regs\[25\]\[30\] _06596_ _06603_ VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__mux2_1
X_13297_ _07153_ VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__buf_6
X_16085_ is_lb_lh_lw_lbu_lhu _02752_ _03635_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09348__A2 _04079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15036_ irq_mask\[27\] _01865_ _01900_ _01891_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__a211o_1
X_12248_ cpuregs.regs\[24\]\[31\] _06598_ _06533_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12179_ _06165_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__buf_2
XANTENNA__10363__B1 instr_rdcycleh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09335__A _04069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16987_ clknet_leaf_12_clk _00161_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16867__S _03174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18726_ net99 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_160_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15938_ mem_rdata_q\[15\] _02638_ _02662_ _02663_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_88_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11863__A0 _06312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08954__S1 _03643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15869_ instr_bge _02618_ _02622_ _02625_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__a22o_1
X_08410_ net66 VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__clkinv_4
XANTENNA__13291__S _07165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17608_ clknet_leaf_173_clk _00777_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09390_ _00070_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09808__B1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18588_ clknet_leaf_166_clk _01653_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17539_ clknet_leaf_11_clk _00708_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15800__A _08033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13368__A0 _04036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14416__A decoded_imm_j\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12040__A0 _06193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16334__C _06083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15109__A1 _05288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11759__B reg_pc\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08890__S0 _03653_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11146__A2 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16609__A1 _06077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12370__S _06663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09726_ reg_pc\[9\] decoded_imm\[9\] VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__and2_1
XANTENNA__09511__A2 _04241_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09657_ instr_rdcycleh count_cycle\[39\] _03252_ _04385_ VGND VGND VPWR VPWR _04386_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08945__S1 _03643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11714__S _06258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08608_ _03383_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__clkbuf_1
X_09588_ cpuregs.regs\[28\]\[6\] cpuregs.regs\[29\]\[6\] cpuregs.regs\[30\]\[6\] cpuregs.regs\[31\]\[6\]
+ _04274_ _04317_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__mux4_1
XANTENNA__16793__A0 _06575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15596__A1 decoded_imm\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15596__B2 _02426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10409__A1 reg_pc\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08539_ is_beq_bne_blt_bge_bltu_bgeu _03317_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16545__A0 _06947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11550_ _06116_ reg_next_pc\[4\] _06119_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13359__A0 _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10501_ net57 _04811_ _04667_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11481_ irq_mask\[28\] _03428_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__or2_1
XANTENNA__12545__S _06752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13220_ _07135_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__clkbuf_1
X_10432_ _05138_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__inv_2
XANTENNA__09578__A2 _04308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13151_ _06974_ cpuregs.regs\[4\]\[15\] _07093_ VGND VGND VPWR VPWR _07099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10363_ count_instr\[59\] _04015_ instr_rdcycleh count_cycle\[59\] VGND VGND VPWR
+ VPWR _05072_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12102_ _06506_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13082_ _07062_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14323__A2 _07997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10294_ cpuregs.regs\[12\]\[25\] cpuregs.regs\[13\]\[25\] cpuregs.regs\[14\]\[25\]
+ cpuregs.regs\[15\]\[25\] _04325_ _04277_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__mux4_1
XANTENNA__13531__A0 _04532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13376__S _07225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12033_ _06166_ cpuregs.regs\[22\]\[9\] _06460_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__mux2_1
X_16910_ clknet_leaf_35_clk _00055_ VGND VGND VPWR VPWR mem_rdata_q\[29\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__12280__S _06615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17890_ clknet_leaf_92_clk _01059_ VGND VGND VPWR VPWR count_cycle\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16841_ _03164_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16687__S _03076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15591__S _02110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16772_ _06554_ cpuregs.regs\[13\]\[10\] _03127_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__mux2_1
X_13984_ count_instr\[0\] _07755_ VGND VGND VPWR VPWR _07756_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18511_ clknet_leaf_20_clk _01576_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10648__A1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15723_ timer\[17\] _02527_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__and2b_1
XFILLER_0_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12935_ _06977_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output213_A net213 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18442_ clknet_leaf_97_clk _01507_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ timer\[0\] _03427_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12866_ _06289_ cpuregs.regs\[6\]\[24\] _06928_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14605_ _07754_ _08257_ _07984_ _08035_ _08258_ VGND VGND VPWR VPWR _08259_ sky130_fd_sc_hd__o32a_1
X_18373_ clknet_leaf_141_clk _01438_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_11817_ _06132_ cpuregs.regs\[11\]\[5\] _06348_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15585_ _02414_ _02415_ _01907_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09266__A1 _03892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12797_ cpuregs.regs\[9\]\[24\] _06584_ _06891_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17324_ clknet_leaf_151_clk _00498_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _08071_ _08190_ _08191_ _08195_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08933__S _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11748_ _06296_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__buf_2
XFILLER_0_138_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16000__A2 _03636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17255_ clknet_leaf_142_clk _00429_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15434__S1 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12455__S _06677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14467_ _08130_ _08126_ _08127_ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__and3_1
X_11679_ reg_pc\[17\] reg_pc\[16\] _06210_ reg_pc\[18\] VGND VGND VPWR VPWR _06235_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16206_ net299 _02824_ _02825_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__nor3_1
XANTENNA__13140__A _07081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13418_ _07209_ VGND VGND VPWR VPWR _07281_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10259__S0 _04329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17186_ clknet_leaf_185_clk _00360_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14398_ reg_next_pc\[7\] _07947_ _08068_ _08033_ VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12573__A1 _06575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16137_ _02770_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__clkbuf_4
X_13349_ _07215_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15198__S0 _03649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09764__S _04320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14314__A2 _07972_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16068_ _02748_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__buf_2
X_15019_ _04805_ _01885_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__nor2_1
XANTENNA__12190__S _06555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08890_ _03644_ _03648_ _03650_ _03651_ _03653_ _03654_ VGND VGND VPWR VPWR _03655_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09065__A _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16597__S _03026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12089__A0 _06114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09511_ _04168_ _04241_ _04242_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11534__S _06086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09442_ _04173_ _04174_ _04077_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_2_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09373_ count_cycle\[1\] _04014_ _04107_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09009__A1 mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11489__B net262 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14553__A2 _07952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13761__B1 _07225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15189__S0 _03670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput250 net250 VGND VGND VPWR VPWR mem_la_wdata[3] sky130_fd_sc_hd__buf_1
XANTENNA__11119__A2 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput261 net261 VGND VGND VPWR VPWR mem_la_wstrb[3] sky130_fd_sc_hd__buf_1
XANTENNA__13196__S _07118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10590__A3 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput272 net272 VGND VGND VPWR VPWR mem_wdata[18] sky130_fd_sc_hd__buf_1
XFILLER_0_101_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput283 net283 VGND VGND VPWR VPWR mem_wdata[28] sky130_fd_sc_hd__clkbuf_1
XANTENNA__10327__B1 net301 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput294 net294 VGND VGND VPWR VPWR mem_wdata[9] sky130_fd_sc_hd__buf_1
XANTENNA__09193__A0 _03940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16058__A2 decoded_imm_j\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09732__A2 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09709_ cpuregs.regs\[8\]\[9\] cpuregs.regs\[9\]\[9\] cpuregs.regs\[10\]\[9\] cpuregs.regs\[11\]\[9\]
+ _04274_ _04317_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__mux4_1
XANTENNA__09703__A _04369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10981_ _03573_ _04848_ _05663_ _05323_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12720_ _06297_ cpuregs.regs\[12\]\[25\] _06847_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12651_ _06297_ cpuregs.regs\[30\]\[25\] _06810_ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__mux2_1
XANTENNA__09248__A1 _03987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11602_ _06166_ cpuregs.regs\[10\]\[9\] _06086_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__mux2_1
X_15370_ _02208_ _02210_ _02213_ _02088_ _02020_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__a221o_1
X_12582_ _06779_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14321_ _03366_ _03319_ VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__nor2_4
XANTENNA__15416__S1 _02047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11533_ _06104_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__buf_2
XANTENNA__10584__A _05244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17040_ clknet_leaf_164_clk _00214_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11464_ _06041_ irq_pending\[20\] _06050_ net13 VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__a31o_1
X_14252_ reg_pc\[17\] _07926_ _07943_ _07935_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11358__A2 _03636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13203_ _07126_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__clkbuf_1
X_10415_ cpuregs.regs\[28\]\[29\] cpuregs.regs\[29\]\[29\] cpuregs.regs\[30\]\[29\]
+ cpuregs.regs\[31\]\[29\] _04579_ _04284_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__mux4_1
X_14183_ count_instr\[61\] _07890_ _07877_ VGND VGND VPWR VPWR _07894_ sky130_fd_sc_hd__o21ai_1
X_11395_ _03822_ _05996_ _06004_ _05976_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10030__A2 _04008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13134_ _06957_ cpuregs.regs\[4\]\[7\] _07082_ VGND VGND VPWR VPWR _07090_ sky130_fd_sc_hd__mux2_1
X_10346_ _05053_ _05054_ _04211_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__mux2_1
XANTENNA__13504__A0 _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12307__A1 _06586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_312 VGND VGND VPWR VPWR alphacore_312/HI cpi_insn[10] sky130_fd_sc_hd__conb_1
Xalphacore_323 VGND VGND VPWR VPWR alphacore_323/HI cpi_insn[21] sky130_fd_sc_hd__conb_1
X_17942_ clknet_leaf_67_clk _08383_ VGND VGND VPWR VPWR reg_out\[22\] sky130_fd_sc_hd__dfxtp_1
X_13065_ _07053_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__clkbuf_1
X_10277_ _04984_ _04987_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10318__B1 _04080_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_334 VGND VGND VPWR VPWR alphacore_334/HI cpi_valid sky130_fd_sc_hd__conb_1
XFILLER_0_29_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xalphacore_345 VGND VGND VPWR VPWR alphacore_345/HI trace_data[6] sky130_fd_sc_hd__conb_1
Xalphacore_356 VGND VGND VPWR VPWR alphacore_356/HI trace_data[17] sky130_fd_sc_hd__conb_1
X_12016_ _06461_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__clkbuf_1
Xalphacore_367 VGND VGND VPWR VPWR alphacore_367/HI trace_data[28] sky130_fd_sc_hd__conb_1
XANTENNA__09723__A2 _04447_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17873_ clknet_leaf_88_clk _01042_ VGND VGND VPWR VPWR count_cycle\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15257__B1 _02006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11530__A2 reg_next_pc\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16824_ _03155_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16755_ _06538_ cpuregs.regs\[13\]\[2\] _03116_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__mux2_1
X_13967_ _03341_ _07727_ _07728_ net150 VGND VGND VPWR VPWR _07744_ sky130_fd_sc_hd__a22o_1
XANTENNA__14480__A1 _07986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10716__S1 _05414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15706_ _08335_ _02517_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__nor2_1
X_12918_ _06183_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__buf_2
XANTENNA__16757__A0 _06540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16686_ _03081_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13898_ _03321_ _07678_ _07682_ net159 VGND VGND VPWR VPWR _07696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15024__A3 _04871_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18425_ clknet_leaf_187_clk _01490_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15637_ _03298_ _03410_ _03400_ _03277_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12849_ _06224_ cpuregs.regs\[6\]\[16\] _06917_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14232__A1 reg_next_pc\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16446__A _02931_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18356_ clknet_leaf_52_clk _00063_ VGND VGND VPWR VPWR reg_sh\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15568_ cpuregs.regs\[8\]\[28\] cpuregs.regs\[9\]\[28\] cpuregs.regs\[10\]\[28\]
+ cpuregs.regs\[11\]\[28\] _02030_ _02031_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15980__A1 _03891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_173_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08998__A0 mem_rdata_q\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17307_ clknet_leaf_13_clk _00481_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10254__C1 _04328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14519_ _08176_ _08179_ VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__or2_2
XFILLER_0_127_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18287_ clknet_leaf_38_clk _01355_ VGND VGND VPWR VPWR mem_state\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08462__A2 irq_active VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15499_ _01989_ _02334_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17238_ clknet_leaf_125_clk _00412_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15732__A1 _04806_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14535__A2 _07904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11349__A2 _03767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17169_ clknet_leaf_115_clk _00343_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09991_ net40 _04710_ _04667_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08942_ _03638_ _03703_ _03705_ _03400_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__o22a_1
XANTENNA__12214__A _06533_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08873_ _03637_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15248__B1 _01963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15343__S0 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12665__A_N _06081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09425_ _04157_ _04158_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15260__A _03664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13699__B decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09356_ _04058_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11588__A2 _03359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09287_ _04023_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12095__S _06496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10608__S _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16790__S _03127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15184__C1 _01969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12537__A1 _06540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10200_ net47 _04745_ _04666_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__a21o_1
X_11180_ reg_next_pc\[2\] reg_out\[2\] _03189_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__mux2_2
XANTENNA__08602__A _03378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10131_ count_cycle\[20\] _04014_ _04846_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__a21o_1
XANTENNA__11760__A2 reg_pc\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10062_ _04268_ _04757_ _04779_ _03302_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__o211a_1
XFILLER_0_100_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14870_ count_cycle\[58\] _01798_ _01800_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13821_ cpuregs.regs\[0\]\[7\] VGND VGND VPWR VPWR _07650_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_35_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16540_ _03003_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__clkbuf_8
X_13752_ _05044_ _05260_ _07560_ _07279_ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__o211a_1
X_10964_ _05377_ _05603_ _05645_ _05251_ _05648_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_63_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12703_ _06232_ cpuregs.regs\[12\]\[17\] _06836_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16471_ cpuregs.waddr\[2\] _06082_ _06601_ _06081_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__and4bb_4
X_13683_ _07511_ _07515_ _07526_ _03311_ VGND VGND VPWR VPWR _07528_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10895_ _03619_ _05583_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18210_ clknet_leaf_43_clk _01281_ VGND VGND VPWR VPWR instr_sltu sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15422_ cpuregs.regs\[28\]\[19\] cpuregs.regs\[29\]\[19\] cpuregs.regs\[30\]\[19\]
+ cpuregs.regs\[31\]\[19\] _03661_ _03662_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__mux4_1
X_12634_ _06232_ cpuregs.regs\[30\]\[17\] _06799_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18141_ clknet_leaf_47_clk alu_out\[15\] VGND VGND VPWR VPWR alu_out_q\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15353_ decoded_imm\[15\] _02009_ _02197_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__a21o_1
X_12565_ _06770_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14304_ irq_pending\[0\] irq_pending\[1\] irq_pending\[2\] irq_pending\[3\] VGND
+ VGND VPWR VPWR _07981_ sky130_fd_sc_hd__or4_1
XFILLER_0_163_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18072_ clknet_leaf_73_clk _01177_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dfxtp_2
X_11516_ _06071_ reg_next_pc\[1\] _03351_ _06072_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15284_ _02020_ _02124_ _02132_ _01960_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__o211a_2
X_12496_ _06733_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17023_ clknet_leaf_181_clk _00197_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14235_ reg_next_pc\[12\] _05858_ _07901_ _07931_ VGND VGND VPWR VPWR _07932_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_150_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11447_ _03305_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output88_A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14166_ _07881_ _07882_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11378_ cpuregs.raddr2\[4\] _03636_ _05986_ _05988_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__o22a_1
X_10329_ irq_mask\[26\] _04448_ timer\[26\] _04187_ _04027_ VGND VGND VPWR VPWR _05039_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13117_ _07080_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_111_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _06053_ VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15573__S0 _01918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ clknet_leaf_61_clk _08396_ VGND VGND VPWR VPWR reg_out\[5\] sky130_fd_sc_hd__dfxtp_1
X_13048_ cpuregs.regs\[3\]\[31\] _06598_ _07009_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11873__A cpuregs.waddr\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17856_ clknet_leaf_101_clk _01025_ VGND VGND VPWR VPWR count_cycle\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15325__S0 _02085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09343__A _04077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16807_ _06590_ cpuregs.regs\[13\]\[27\] _03138_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__mux2_1
XANTENNA__14989__C1 _08335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17787_ clknet_leaf_84_clk _00956_ VGND VGND VPWR VPWR count_instr\[58\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__16875__S _03174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14999_ _01862_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16738_ _03108_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08407__A_N _03191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09555__S1 _04285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16669_ cpuregs.regs\[1\]\[29\] _06327_ _03062_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__mux2_1
XANTENNA__14205__A1 reg_next_pc\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09880__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09880__B2 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11019__A1 _05458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09210_ _03953_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__clkbuf_1
X_18408_ clknet_leaf_149_clk _01473_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10227__C1 _04100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09141_ _03895_ _03863_ _03870_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18339_ clknet_leaf_37_clk _01407_ VGND VGND VPWR VPWR mem_16bit_buffer\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10428__S _04320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08435__A2 _03219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08406__B mem_do_prefetch VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09072_ _03818_ _03770_ _03833_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__or3b_1
XANTENNA__15705__A1 _04561_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12643__S _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_153_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09974_ cpuregs.regs\[8\]\[16\] cpuregs.regs\[9\]\[16\] cpuregs.regs\[10\]\[16\]
+ cpuregs.regs\[11\]\[16\] _04057_ _04060_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10950__B1 _05213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09148__B1 _03878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13982__B decoder_trigger VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08925_ cpuregs.regs\[4\]\[3\] cpuregs.regs\[5\]\[3\] cpuregs.regs\[6\]\[3\] cpuregs.regs\[7\]\[3\]
+ _03658_ _03659_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__mux4_1
XANTENNA__13495__A2 decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09699__B2 _04426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11783__A _06327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08856_ _03616_ _03526_ _03620_ _03621_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__and4bb_1
XANTENNA__15316__S0 _01985_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09794__S1 _04285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_168_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08787_ net100 net68 VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__and2b_1
XANTENNA__10399__A _05106_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14995__A2 _01863_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16197__A1 net257 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12818__S _06906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09871__B2 _04024_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09408_ _04127_ _04131_ _04133_ _04141_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__o211ai_4
X_10680_ _05379_ _05380_ _05242_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_80_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14318__B _07994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09339_ _04073_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10233__A2 _04745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12350_ _06655_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11301_ _05920_ _05923_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__nor2_1
X_12281_ _06618_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11232_ reg_next_pc\[11\] reg_out\[11\] _05858_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__mux2_2
X_14020_ count_instr\[11\] count_instr\[10\] count_instr\[9\] _07773_ VGND VGND VPWR
+ VPWR _07781_ sky130_fd_sc_hd__and4_2
XANTENNA__09428__A _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11163_ _05816_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16121__A1 _05324_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15555__S0 _02111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09139__B1 _03895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10114_ cpuregs.regs\[4\]\[20\] cpuregs.regs\[5\]\[20\] cpuregs.regs\[6\]\[20\] cpuregs.regs\[7\]\[20\]
+ _04275_ _04278_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_73_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11094_ _05219_ _05762_ _05769_ VGND VGND VPWR VPWR alu_out\[28\] sky130_fd_sc_hd__o21ai_2
X_15971_ mem_rdata_q\[25\] _02610_ _02671_ _02689_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_73_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17710_ clknet_leaf_75_clk _00879_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dfxtp_1
XANTENNA__11693__A _06247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10045_ _04430_ _04760_ _04762_ _04070_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__o211a_1
X_14922_ net196 net165 _01835_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_10_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15307__S0 _01990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17641_ clknet_leaf_46_clk _00810_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_1
X_14853_ count_cycle\[52\] count_cycle\[53\] _01786_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16695__S _03076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output126_A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13804_ _07232_ _07637_ _07638_ _07639_ _07640_ VGND VGND VPWR VPWR _07641_ sky130_fd_sc_hd__o41a_1
X_17572_ clknet_leaf_16_clk _00741_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10102__A reg_pc\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14784_ _01741_ _08350_ _01742_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__and3b_1
XFILLER_0_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11996_ _06450_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09311__B1 _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16523_ cpuregs.regs\[17\]\[24\] _06584_ _02990_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__mux2_1
X_13735_ _05013_ _07576_ _07224_ VGND VGND VPWR VPWR _07577_ sky130_fd_sc_hd__mux2_1
XANTENNA__16188__A1 net257 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10947_ _04754_ _04744_ _05230_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__mux2_1
XANTENNA__12728__S _06847_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_119_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11632__S _06176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13413__A _05209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14199__B1 _07906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16454_ _02958_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__clkbuf_1
X_13666_ net80 decoded_imm\[21\] VGND VGND VPWR VPWR _07512_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10878_ _03560_ _05567_ _05363_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08507__A _03276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12749__A1 _06536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15405_ _02245_ _02246_ _03713_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12617_ _06166_ cpuregs.regs\[30\]\[9\] _06788_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16385_ _06991_ cpuregs.regs\[16\]\[23\] _02918_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__mux2_1
X_13597_ _07418_ _07422_ _07432_ VGND VGND VPWR VPWR _07448_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18124_ clknet_leaf_40_clk _01228_ VGND VGND VPWR VPWR latched_is_lb sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15336_ decoded_imm\[14\] _02009_ _01963_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__a21o_1
X_12548_ _06761_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18055_ clknet_leaf_59_clk _01160_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_113_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15267_ _02109_ _02113_ _02116_ _02037_ _01969_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__a221o_1
X_12479_ _06724_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_2 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17006_ clknet_leaf_123_clk _00180_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_14218_ _05856_ _06143_ VGND VGND VPWR VPWR _07920_ sky130_fd_sc_hd__or2_1
XANTENNA__09917__A2 _04049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15198_ cpuregs.regs\[20\]\[7\] cpuregs.regs\[21\]\[7\] cpuregs.regs\[22\]\[7\] cpuregs.regs\[23\]\[7\]
+ _03649_ _03643_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14149_ _07869_ _07815_ _07870_ VGND VGND VPWR VPWR _07871_ sky130_fd_sc_hd__and3b_1
XANTENNA__10083__S1 _04283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14898__B net257 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08710_ net109 net77 VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__nor2_1
XANTENNA__11807__S _06348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11488__A1 _06054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17908_ clknet_leaf_85_clk _01077_ VGND VGND VPWR VPWR count_cycle\[53\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10711__S _05390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09690_ _04268_ _04397_ _04417_ _04149_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09073__A _03215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08641_ irq_state\[1\] VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17839_ clknet_leaf_61_clk _01008_ VGND VGND VPWR VPWR reg_next_pc\[16\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_117_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08572_ irq_mask\[1\] irq_pending\[1\] VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__and2b_2
XFILLER_0_88_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09801__A _04227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16179__A1 net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12638__S _06799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10999__B1 _05218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15926__A1 _02625_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09124_ _03779_ _03789_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__nor2_1
XANTENNA__10846__S0 _05413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09055_ _03790_ _03816_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11176__B1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15537__S0 _02046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14114__B1 _07834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09957_ _04535_ _04598_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__or2b_1
X_08908_ _03664_ _03672_ _00067_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__o21a_1
X_09888_ _04608_ _04609_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_51_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08839_ _03474_ _03489_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_51_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11018__A _05219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11850_ _06371_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15090__A1 _03719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10801_ _03515_ _05495_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11781_ _06252_ _03337_ _06253_ _06325_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13520_ net69 decoded_imm\[11\] VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__nand2_1
X_10732_ _05428_ _05429_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13451_ _07310_ _07311_ VGND VGND VPWR VPWR _07312_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10663_ _03540_ _05362_ _05363_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12402_ _06683_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__clkbuf_1
X_16170_ _02803_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__clkbuf_1
X_10594_ _05292_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__or2_1
X_13382_ _07243_ _07244_ _07246_ VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15121_ _01918_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_11_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12333_ _06646_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15052_ _03666_ _01911_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_75_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12264_ _06609_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_75_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15594__S _02110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14003_ count_instr\[6\] _07767_ VGND VGND VPWR VPWR _07769_ sky130_fd_sc_hd__and2_1
X_11215_ _05852_ _05853_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__nor2_1
X_12195_ _06207_ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__buf_2
XANTENNA__09592__S _04321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput72 net72 VGND VGND VPWR VPWR cpi_rs1[14] sky130_fd_sc_hd__clkbuf_1
Xoutput83 net83 VGND VGND VPWR VPWR cpi_rs1[24] sky130_fd_sc_hd__buf_1
X_11146_ _03407_ net127 net104 _04422_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__a22o_2
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput94 net94 VGND VGND VPWR VPWR cpi_rs1[5] sky130_fd_sc_hd__buf_1
XANTENNA_output243_A net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14656__A1 _03294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13408__A _07224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11077_ _05323_ _05753_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__nor2_1
X_15954_ _03196_ net299 VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09758__S1 _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09532__A0 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10028_ _03637_ _04744_ _04673_ _04746_ _04266_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__a221o_1
X_14905_ net218 net187 _01824_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__mux2_1
X_15885_ _02611_ _02620_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__and2_1
XANTENNA__14408__A1 _03378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14408__B2 _03293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14836_ count_cycle\[46\] _01774_ count_cycle\[47\] VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17624_ clknet_leaf_109_clk _00793_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13616__C1 _07217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08936__S _03664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_127_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ clknet_leaf_154_clk _00724_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_14767_ count_cycle\[25\] _01729_ _01717_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14239__A _03294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09835__A1 _04068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11979_ _06441_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16506_ cpuregs.regs\[17\]\[16\] _06567_ _02979_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__mux2_1
XANTENNA__10445__A2 _04104_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13718_ _04945_ _05258_ _07517_ _07237_ VGND VGND VPWR VPWR _07561_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17486_ clknet_leaf_136_clk _00655_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14698_ count_cycle\[3\] _08337_ _07877_ VGND VGND VPWR VPWR _08341_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09930__S1 _04233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16437_ _02949_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13649_ _04708_ _05261_ _07495_ _07274_ VGND VGND VPWR VPWR _07496_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13797__B decoded_imm\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16368_ _06974_ cpuregs.regs\[16\]\[15\] _02907_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18107_ clknet_leaf_89_clk _01211_ VGND VGND VPWR VPWR timer\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13289__S _07165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15319_ _02153_ _02157_ _02027_ _02165_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__o211a_4
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_12 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12193__S _06555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16299_ _06974_ cpuregs.regs\[15\]\[15\] _02870_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_120_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_120_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18038_ clknet_leaf_80_clk _00015_ VGND VGND VPWR VPWR irq_pending\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11158__A0 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11110__B _05143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15519__S0 _02085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09811_ reg_pc\[12\] decoded_imm\[12\] VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__nand2_1
XANTENNA__09771__B1 _03252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10381__A1 _04105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14421__B _07988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09742_ _04420_ _04467_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__or2_2
XANTENNA__09523__B1 _04254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10133__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09673_ cpuregs.regs\[8\]\[8\] cpuregs.regs\[9\]\[8\] cpuregs.regs\[10\]\[8\] cpuregs.regs\[11\]\[8\]
+ _04056_ _04091_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_187_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_187_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_143_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16629__A _03039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _03309_ _03385_ _03237_ _03251_ _03398_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__a41o_1
XANTENNA__15533__A _03709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09531__A _03524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13083__A0 _06974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08555_ _03330_ _03331_ _03332_ _03333_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__or4_1
XANTENNA__12368__S _06663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13622__A2 _04777_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12830__A0 _06150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08486_ _03269_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13988__A _06053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13386__A1 _07209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_746 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09107_ _03832_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10295__S1 _04277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_111_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_115_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09038_ _03799_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09437__S0 _04056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13689__A2 _04909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10047__S1 _04473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16303__S _02870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16088__B1 _02634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11000_ net81 _04880_ _05236_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08610__A _03384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _06988_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_178_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_178_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__10124__A1 _04215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11902_ _06400_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10675__A2 _04039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15670_ timer\[2\] _02483_ timer\[3\] VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__o21ai_1
X_12882_ _06077_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__buf_2
XFILLER_0_169_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15063__A1 _01907_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14621_ _08272_ _08273_ VGND VGND VPWR VPWR _08274_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11833_ _06362_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12278__S _06615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ clknet_leaf_16_clk _00087_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__dfxtp_4
X_14552_ _08208_ _08209_ VGND VGND VPWR VPWR _08210_ sky130_fd_sc_hd__nor2_1
X_11764_ _06116_ reg_next_pc\[27\] _06308_ _06310_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13503_ _07356_ _07357_ _07359_ _07360_ VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__o31a_1
X_10715_ _05292_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__buf_4
X_17271_ clknet_leaf_155_clk _00445_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14483_ _08012_ _08142_ _08143_ _08146_ VGND VGND VPWR VPWR _08147_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_101_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11695_ _06249_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16222_ _02835_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__clkbuf_1
X_13434_ _07287_ _07292_ VGND VGND VPWR VPWR _07296_ sky130_fd_sc_hd__or2_1
X_10646_ _05347_ _05262_ _05235_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output193_A net193 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16153_ _02794_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__clkbuf_1
X_13365_ _04037_ decoded_imm\[0\] _07227_ _07228_ VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_102_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_102_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10286__S1 _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10577_ _03612_ _05219_ _05253_ _05280_ VGND VGND VPWR VPWR alu_out\[0\] sky130_fd_sc_hd__o22a_1
X_15104_ _03677_ _01960_ _01961_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12316_ _06636_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__clkbuf_1
X_16084_ _03767_ _03935_ _02751_ _03816_ _03215_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__a32o_1
X_13296_ _07175_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__clkbuf_1
X_15035_ _05069_ _01885_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12247_ _06342_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__buf_2
XANTENNA__14522__A _07998_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output70_A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12178_ _06551_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11560__B1 _06098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15826__B1 _03747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11129_ _03433_ _05440_ _05357_ _03434_ _05801_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__o221a_1
XANTENNA__10261__S _04222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16986_ clknet_leaf_189_clk _00160_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_169_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_169_clk sky130_fd_sc_hd__clkbuf_2
X_15937_ mem_rdata_q\[5\] mem_rdata_q\[4\] mem_rdata_q\[6\] VGND VGND VPWR VPWR _02663_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_160_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11312__B1 _05932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09600__S0 _04329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15868_ _02624_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__buf_2
XANTENNA__16251__A0 mem_rdata_q\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14819_ _01765_ _01753_ _01766_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__and3b_1
X_17607_ clknet_leaf_178_clk _00776_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09808__A1 _04149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18587_ clknet_leaf_187_clk _01652_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_15799_ _02583_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09808__B2 _04532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17538_ clknet_leaf_188_clk _00707_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11091__A2 _05220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17469_ clknet_leaf_114_clk _00638_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15800__B _07994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12916__S _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13368__A1 _04160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14565__B1 _07952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15109__A2 _01963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16334__D _06081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12217__A _06265_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08890__S1 _03654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__16123__S _02771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12651__S _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13540__A1 _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_985 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09725_ reg_pc\[9\] decoded_imm\[9\] VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__nor2_1
XANTENNA__12887__A _06095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10657__A2 _05222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09656_ count_instr\[39\] instr_rdinstrh instr_rdinstr count_instr\[7\] VGND VGND
+ VPWR VPWR _04385_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08607_ _03250_ _03381_ _00865_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__or3_1
XANTENNA__13056__A0 _06947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09587_ _04283_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__buf_4
XANTENNA__16793__S _03138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14399__A3 _07992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15596__A2 _02216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10409__A2 decoded_imm\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08538_ cpu_state\[3\] VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__inv_2
XANTENNA__11606__A1 _06116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08469_ instr_rdinstrh instr_rdinstr instr_rdcycleh VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__nor3_4
XTAP_TAPCELL_ROW_34_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12826__S _06906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10500_ net91 VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__buf_4
XFILLER_0_135_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11480_ _06054_ irq_pending\[27\] _06059_ net20 VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__a31o_1
XANTENNA__08605__A _03277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14326__B _07997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10431_ _05125_ _05129_ _04100_ _05137_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__a211o_2
XANTENNA__10346__S _04211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13150_ _07098_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__clkbuf_1
X_10362_ irq_mask\[27\] _04448_ timer\[27\] _04187_ _04188_ VGND VGND VPWR VPWR _05071_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11790__B1 _06098_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12101_ _06166_ cpuregs.regs\[23\]\[9\] _06496_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13081_ _06972_ cpuregs.regs\[7\]\[14\] _07057_ VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__mux2_1
X_10293_ _04430_ _05003_ _04214_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12032_ _06469_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09830__S0 _04329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16840_ _06554_ cpuregs.regs\[14\]\[10\] _03163_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__mux2_1
XANTENNA__15284__A1 _02020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16771_ _03115_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__buf_6
X_13983_ _03363_ _07754_ cpu_state\[1\] _03376_ VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__and4b_2
X_15722_ timer\[16\] _02524_ timer\[17\] VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__o21a_1
XANTENNA__11905__S _06398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18510_ clknet_leaf_107_clk _01575_ VGND VGND VPWR VPWR cpuregs.regs\[18\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15173__A _01959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10648__A2 _04198_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12934_ _06976_ cpuregs.regs\[31\]\[16\] _06964_ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16233__A0 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15653_ _02476_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__clkbuf_4
X_18441_ clknet_leaf_98_clk _01506_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12865_ _06932_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_103_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output206_A net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14604_ _08257_ _08246_ VGND VGND VPWR VPWR _08258_ sky130_fd_sc_hd__nor2_1
X_11816_ _06353_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__clkbuf_1
X_18372_ clknet_leaf_129_clk _01437_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_15584_ cpuregs.regs\[0\]\[29\] cpuregs.regs\[1\]\[29\] cpuregs.regs\[2\]\[29\] cpuregs.regs\[3\]\[29\]
+ _01908_ _01909_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_83_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _06895_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09897__S0 _04216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17323_ clknet_leaf_151_clk _00497_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14535_ reg_next_pc\[18\] _07904_ _08121_ _08192_ _08194_ VGND VGND VPWR VPWR _08195_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__11073__A2 _05357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11747_ _06226_ reg_next_pc\[25\] _06293_ _06295_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__a211o_2
XFILLER_0_28_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14517__A decoded_imm_j\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13421__A _07283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17254_ clknet_leaf_137_clk _00428_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14466_ _08126_ _08127_ _08130_ VGND VGND VPWR VPWR _08131_ sky130_fd_sc_hd__a21oi_2
X_11678_ reg_pc\[18\] reg_pc\[17\] _06218_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09649__S0 _04216_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16205_ _03187_ net33 net44 _02823_ clear_prefetched_high_word VGND VGND VPWR VPWR
+ _02825_ sky130_fd_sc_hd__a41o_1
XFILLER_0_52_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13417_ _04262_ _07277_ _07278_ _07279_ VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__o211a_1
X_10629_ _05295_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__clkbuf_4
X_17185_ clknet_leaf_189_clk _00359_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10259__S1 _04218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14397_ _07921_ _07994_ _08067_ VGND VGND VPWR VPWR _08068_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_153_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16136_ _02785_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__clkbuf_1
X_13348_ cpu_state\[4\] _03399_ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15198__S1 _03643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16067_ _02610_ _02747_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__and2_1
X_13279_ _06966_ cpuregs.regs\[5\]\[11\] _07165_ VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__mux2_1
X_15018_ irq_mask\[18\] _01880_ _01890_ _01891_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__a211o_1
XANTENNA__09346__A _04080_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10336__A1 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10336__B2 _05045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09821__S0 _04085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10887__A2 _05357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16969_ clknet_leaf_142_clk _00143_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11815__S _06348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09510_ irq_mask\[4\] _04021_ timer\[4\] _04187_ _04188_ VGND VGND VPWR VPWR _04242_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09081__A _03841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09441_ cpuregs.regs\[16\]\[3\] cpuregs.regs\[17\]\[3\] cpuregs.regs\[18\]\[3\] cpuregs.regs\[19\]\[3\]
+ _04071_ _04073_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__mux4_1
X_18639_ clknet_leaf_180_clk _01699_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14786__B1 _01717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09372_ count_instr\[1\] _04012_ _04009_ _04106_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12261__A1 _06540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16527__A1 _06588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10976__A1_N _05404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11489__C _03305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14553__A3 _08050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13761__A1 _03631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15189__S1 _03671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10690__A _05323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput240 net240 VGND VGND VPWR VPWR mem_la_wdata[23] sky130_fd_sc_hd__buf_1
Xoutput251 net251 VGND VGND VPWR VPWR mem_la_wdata[4] sky130_fd_sc_hd__buf_1
XANTENNA__13513__A1 _07274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput262 net262 VGND VGND VPWR VPWR mem_valid sky130_fd_sc_hd__buf_1
Xoutput273 net273 VGND VGND VPWR VPWR mem_wdata[19] sky130_fd_sc_hd__clkbuf_1
XANTENNA__16788__S _03127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput284 net284 VGND VGND VPWR VPWR mem_wdata[29] sky130_fd_sc_hd__clkbuf_1
Xoutput295 net295 VGND VGND VPWR VPWR mem_wstrb[0] sky130_fd_sc_hd__clkbuf_1
XANTENNA__09193__A1 _03891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13506__A _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09708_ cpuregs.regs\[12\]\[9\] cpuregs.regs\[13\]\[9\] cpuregs.regs\[14\]\[9\] cpuregs.regs\[15\]\[9\]
+ _04274_ _04317_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10980_ _03466_ _03572_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__nor2_1
XANTENNA__16215__A0 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09639_ cpuregs.regs\[12\]\[7\] cpuregs.regs\[13\]\[7\] cpuregs.regs\[14\]\[7\] cpuregs.regs\[15\]\[7\]
+ _04290_ _04276_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14777__B1 _01717_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12650_ _06815_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11601_ _06165_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__buf_2
XANTENNA__11055__A2 _05397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12556__S _06763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12581_ cpuregs.regs\[2\]\[24\] _06584_ _06774_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14320_ _07996_ VGND VGND VPWR VPWR _07997_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_61_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11532_ _06100_ _06102_ _06103_ _06093_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__o22a_2
XFILLER_0_147_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14251_ _05909_ _06229_ _07942_ _05893_ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__o211a_2
XFILLER_0_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11463_ irq_mask\[20\] _06042_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13202_ _06957_ cpuregs.regs\[8\]\[7\] _07118_ VGND VGND VPWR VPWR _07126_ sky130_fd_sc_hd__mux2_1
XANTENNA__13752__A1 _05044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10414_ _04018_ count_cycle\[61\] _04014_ count_cycle\[29\] _05120_ VGND VGND VPWR
+ VPWR _05121_ sky130_fd_sc_hd__a221o_1
X_14182_ count_instr\[61\] count_instr\[60\] count_instr\[59\] _07887_ VGND VGND VPWR
+ VPWR _07893_ sky130_fd_sc_hd__and4_2
XFILLER_0_33_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11394_ _03781_ _06003_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10110__S0 _04275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13387__S _05257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13133_ _07089_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15168__A _01936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10345_ cpuregs.regs\[24\]\[27\] cpuregs.regs\[25\]\[27\] cpuregs.regs\[26\]\[27\]
+ cpuregs.regs\[27\]\[27\] _04758_ _04759_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__mux4_1
XFILLER_0_104_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xalphacore_302 VGND VGND VPWR VPWR alphacore_302/HI cpi_insn[0] sky130_fd_sc_hd__conb_1
Xalphacore_313 VGND VGND VPWR VPWR alphacore_313/HI cpi_insn[11] sky130_fd_sc_hd__conb_1
X_17941_ clknet_leaf_67_clk _08382_ VGND VGND VPWR VPWR reg_out\[21\] sky130_fd_sc_hd__dfxtp_1
X_13064_ _06955_ cpuregs.regs\[7\]\[6\] _07046_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__mux2_1
Xalphacore_324 VGND VGND VPWR VPWR alphacore_324/HI cpi_insn[22] sky130_fd_sc_hd__conb_1
X_10276_ _04985_ _04986_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__nor2_1
XANTENNA__10318__A1 _04068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_335 VGND VGND VPWR VPWR alphacore_335/HI mem_addr[0] sky130_fd_sc_hd__conb_1
XANTENNA__16698__S _03087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xalphacore_346 VGND VGND VPWR VPWR alphacore_346/HI trace_data[7] sky130_fd_sc_hd__conb_1
X_12015_ _06078_ cpuregs.regs\[22\]\[0\] _06460_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__mux2_1
XANTENNA__09184__B2 _03888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_357 VGND VGND VPWR VPWR alphacore_357/HI trace_data[18] sky130_fd_sc_hd__conb_1
Xalphacore_368 VGND VGND VPWR VPWR alphacore_368/HI trace_data[29] sky130_fd_sc_hd__conb_1
X_17872_ clknet_leaf_90_clk _01041_ VGND VGND VPWR VPWR count_cycle\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15257__A1 _02020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16823_ _06538_ cpuregs.regs\[14\]\[2\] _03152_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13966_ _07743_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__clkbuf_1
X_16754_ _03118_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10177__S0 _04281_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15705_ _04561_ _02476_ _02515_ _02516_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__a22o_1
X_12917_ _06965_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__clkbuf_1
X_16685_ _06951_ cpuregs.regs\[19\]\[4\] _03076_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__mux2_1
X_13897_ _07695_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_100_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18424_ clknet_leaf_12_clk _01489_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_15636_ cpu_state\[2\] _03254_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__nand2_1
X_12848_ _06923_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18355_ clknet_leaf_52_clk _00062_ VGND VGND VPWR VPWR reg_sh\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12466__S _06715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15567_ cpuregs.regs\[12\]\[28\] cpuregs.regs\[13\]\[28\] cpuregs.regs\[14\]\[28\]
+ cpuregs.regs\[15\]\[28\] _01979_ _01980_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12779_ _06886_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15980__A2 _03767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08998__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17306_ clknet_leaf_188_clk _00480_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_14518_ _08177_ _08178_ VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18286_ clknet_leaf_38_clk _01354_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dfxtp_2
X_15498_ cpuregs.regs\[8\]\[24\] cpuregs.regs\[9\]\[24\] cpuregs.regs\[10\]\[24\]
+ cpuregs.regs\[11\]\[24\] _02013_ _02014_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17237_ clknet_leaf_115_clk _00411_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_14449_ _08113_ _08114_ VGND VGND VPWR VPWR _08115_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14940__A0 net205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17168_ clknet_leaf_110_clk _00342_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16119_ mem_state\[0\] _02774_ _02777_ _02768_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__o22a_1
XANTENNA__15078__A _03646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09990_ _04668_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__clkbuf_4
X_17099_ clknet_leaf_177_clk _00273_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08941_ reg_sh\[3\] reg_sh\[2\] _03704_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_50_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08872_ _03312_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__buf_2
XANTENNA__16401__S _02895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15248__A1 decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15343__S1 _01997_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_91_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_2
X_09424_ _04152_ _04153_ _04155_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__a21o_1
XANTENNA__10493__B1 _04237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11037__A2 _05220_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09355_ _04088_ _04089_ _04078_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__mux2_1
XANTENNA__10685__A _05254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12376__S _06663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09286_ instr_timer VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13734__A1 _07232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_896 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09938__B1 _04100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10548__B2 _05251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08602__B _03379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13000__S _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08829__A_N net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10130_ count_instr\[20\] _04012_ _04009_ _04845_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__a211o_1
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10061_ _04271_ _04777_ _04778_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__a21o_1
XANTENNA__15716__A _02476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16436__A0 _06974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13820_ _07649_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__clkbuf_1
X_13751_ _07591_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__clkbuf_1
X_10963_ _03478_ _05357_ _05647_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_82_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_2
X_12702_ _06843_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16470_ _02966_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_63_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13682_ _07511_ _07515_ _07526_ VGND VGND VPWR VPWR _07527_ sky130_fd_sc_hd__a21oi_1
X_10894_ _03562_ _05582_ _05390_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__mux2_1
XANTENNA__14214__A2 _07906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15421_ _02260_ _02261_ _03653_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12633_ _06806_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12286__S _06615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18140_ clknet_leaf_46_clk alu_out\[14\] VGND VGND VPWR VPWR alu_out_q\[14\] sky130_fd_sc_hd__dfxtp_1
X_15352_ _01934_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12564_ cpuregs.regs\[2\]\[16\] _06567_ _06763_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__mux2_1
XANTENNA__10787__A1 _05225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11984__A0 _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14303_ irq_pending\[4\] irq_pending\[5\] irq_pending\[6\] irq_pending\[7\] VGND
+ VGND VPWR VPWR _07980_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_18071_ clknet_leaf_72_clk _01176_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_170_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11515_ reg_out\[1\] alu_out_q\[1\] latched_stalu VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__mux2_1
X_15283_ _02126_ _02128_ _02131_ _03683_ _02018_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12495_ _06224_ cpuregs.regs\[28\]\[16\] _06726_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17022_ clknet_leaf_171_clk _00196_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_14234_ _05856_ _06190_ VGND VGND VPWR VPWR _07931_ sky130_fd_sc_hd__or2_1
XANTENNA__14922__A0 net196 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09929__B1 _04082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11446_ _06029_ irq_pending\[12\] _06040_ net4 VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_150_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14165_ count_instr\[55\] _07879_ _07877_ VGND VGND VPWR VPWR _07882_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_78_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11377_ _05969_ _03900_ _05987_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13116_ _07007_ cpuregs.regs\[7\]\[31\] _07045_ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__mux2_1
X_10328_ _04051_ _05037_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__nor2_1
XANTENNA__13489__B1 _03631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14096_ count_instr\[35\] _07831_ VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_111_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15573__S1 _01919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09157__A1 _03910_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17924_ clknet_leaf_56_clk _08395_ VGND VGND VPWR VPWR reg_out\[4\] sky130_fd_sc_hd__dfxtp_1
X_13047_ _07043_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__clkbuf_1
X_10259_ cpuregs.regs\[28\]\[24\] cpuregs.regs\[29\]\[24\] cpuregs.regs\[30\]\[24\]
+ cpuregs.regs\[31\]\[24\] _04329_ _04218_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__mux4_1
XANTENNA__11873__B cpuregs.waddr\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17855_ clknet_leaf_102_clk _01024_ VGND VGND VPWR VPWR count_cycle\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__15325__S1 _02086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16806_ _03145_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13336__S0 _04579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17786_ clknet_leaf_84_clk _00955_ VGND VGND VPWR VPWR count_instr\[57\] sky130_fd_sc_hd__dfxtp_1
X_14998_ irq_mask\[10\] _01864_ _01879_ _01876_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__a211o_1
XANTENNA__15650__B2 mem_do_wdata VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16737_ _07003_ cpuregs.regs\[19\]\[29\] _03098_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__mux2_1
X_13949_ _07714_ _07731_ VGND VGND VPWR VPWR _07732_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_73_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16668_ _03071_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18407_ clknet_leaf_156_clk _01472_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12196__S _06555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15619_ _02446_ _02447_ _03653_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16599_ _07001_ cpuregs.regs\[18\]\[28\] _03026_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09140_ _03891_ _03892_ _03880_ _03896_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18338_ clknet_leaf_37_clk _01406_ VGND VGND VPWR VPWR mem_16bit_buffer\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13964__B2 net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10322__S0 _04055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09071_ _03827_ _03832_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__nor2_2
XFILLER_0_126_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15705__A2 _02476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18269_ clknet_leaf_26_clk _01340_ VGND VGND VPWR VPWR decoded_imm\[27\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_32_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14913__A0 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09973_ _04070_ _04692_ _04082_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_168_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08924_ _03685_ _03686_ _03687_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__mux2_1
XANTENNA__16131__S _02771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08855_ _03535_ _03496_ _03499_ _03529_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__and4b_1
XANTENNA__15316__S1 _01986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08786_ _03550_ _03510_ _03515_ _03551_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_146_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15641__A1 _07992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_64_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_138_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16197__A2 net261 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09871__A2 _04448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09407_ _04135_ _04137_ _04140_ _04052_ _00073_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10218__B1 _04296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09338_ _00070_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__buf_4
XFILLER_0_75_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10769__A1 _05361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16091__A_N _03878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09269_ cpu_state\[3\] cpu_state\[6\] _03410_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__or3_4
XFILLER_0_118_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12834__S _06906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14615__A _07942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11300_ reg_out\[24\] _05909_ _05922_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__o21a_1
X_12280_ cpuregs.regs\[25\]\[12\] _06559_ _06615_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11231_ _05829_ _05865_ _05866_ _05867_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__a31o_4
XFILLER_0_121_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10354__S _04211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09428__B _04038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11162_ net128 net114 _04668_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15555__S1 _02004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10113_ _04272_ _04828_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__nand2_1
X_11093_ _05540_ _05700_ _05763_ _05768_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__o211a_1
XANTENNA__12143__A0 _06328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ mem_rdata_q\[2\] mem_rdata_q\[28\] VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__nor2_1
XANTENNA__16409__A0 _06947_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10044_ _04575_ _04761_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__or2_1
X_14921_ _01823_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__15307__S1 _01992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17640_ clknet_leaf_51_clk _00809_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfxtp_2
X_14852_ count_cycle\[52\] _01786_ _01788_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__o21a_1
X_13803_ _07304_ _05170_ _07305_ reg_pc\[30\] _07221_ VGND VGND VPWR VPWR _07640_
+ sky130_fd_sc_hd__a221o_1
X_14783_ count_cycle\[28\] count_cycle\[29\] _01736_ count_cycle\[30\] VGND VGND VPWR
+ VPWR _01742_ sky130_fd_sc_hd__a31o_1
X_17571_ clknet_leaf_15_clk _00740_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10102__B decoded_imm\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11995_ _06281_ cpuregs.regs\[21\]\[23\] _06446_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__mux2_1
XANTENNA_output119_A net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__11913__S _06398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13734_ _07232_ _07572_ _07573_ _07574_ _07575_ VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__o41a_1
XANTENNA__09311__B2 _04046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16522_ _02994_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10946_ _03482_ _05630_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16188__A2 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14199__A1 _07899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13665_ _04880_ decoded_imm\[21\] VGND VGND VPWR VPWR _07511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16453_ _06991_ cpuregs.regs\[29\]\[23\] _02954_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__mux2_1
X_10877_ _03494_ _03497_ _05550_ _03495_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__o31a_1
XFILLER_0_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10209__B1 _04011_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15404_ cpuregs.regs\[24\]\[18\] cpuregs.regs\[25\]\[18\] cpuregs.regs\[26\]\[18\]
+ cpuregs.regs\[27\]\[18\] _03640_ _03642_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__mux4_1
X_12616_ _06797_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16384_ _02921_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__clkbuf_1
X_13596_ _07445_ _07446_ VGND VGND VPWR VPWR _07447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11957__A0 _06132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18123_ clknet_leaf_41_clk _01227_ VGND VGND VPWR VPWR latched_is_lh sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15335_ _01969_ _02172_ _02180_ _01960_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__o211a_4
X_12547_ cpuregs.regs\[2\]\[8\] _06550_ _06752_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15243__S0 _01999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15266_ _02114_ _02115_ _02002_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__mux2_1
X_18054_ clknet_leaf_20_clk _01159_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dfxtp_4
X_12478_ _06157_ cpuregs.regs\[28\]\[8\] _06715_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08523__A _03302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_3 _01973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17005_ clknet_leaf_120_clk _00179_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_14217_ reg_pc\[6\] _07906_ _07919_ _07912_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10264__S _04077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14371__A1 _08035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11429_ irq_mask\[4\] _06030_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_130_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15197_ _02005_ _02043_ _02045_ _02049_ _03639_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__a221o_2
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14148_ count_instr\[49\] _07865_ count_instr\[50\] VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__a21o_1
XANTENNA__10932__A1 _05255_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09025__B_N _03206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__15320__B1 _01963_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14079_ count_instr\[30\] count_instr\[29\] _07818_ VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__and3_1
X_17907_ clknet_leaf_85_clk _01076_ VGND VGND VPWR VPWR count_cycle\[52\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08640_ _03407_ _03299_ _03408_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_128_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17838_ clknet_leaf_61_clk _01007_ VGND VGND VPWR VPWR reg_next_pc\[15\] sky130_fd_sc_hd__dfxtp_1
X_08571_ _03346_ _03347_ _03348_ _03349_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__or4_1
XANTENNA__12437__A1 _06578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17769_ clknet_leaf_95_clk _00938_ VGND VGND VPWR VPWR count_instr\[40\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12919__S _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_46_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_2
XANTENNA__11823__S _06348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13937__A1 _03336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15482__S0 _02046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09066__A0 mem_rdata_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09123_ _03854_ _03870_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__and2b_1
XFILLER_0_162_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15139__B1 _03692_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10846__S1 _05414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09054_ _03800_ _03804_ _03815_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__nor3_4
XFILLER_0_32_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11176__A1 _04038_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__16650__A _03039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11176__B2 _03297_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15537__S1 _02047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10902__S _05244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09956_ _04607_ _04639_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__or2_1
XANTENNA__12125__A0 _06257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08907_ cpuregs.regs\[28\]\[2\] cpuregs.regs\[29\]\[2\] cpuregs.regs\[30\]\[2\] cpuregs.regs\[31\]\[2\]
+ _03670_ _03671_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__mux4_1
X_09887_ _04597_ _04600_ _04607_ _04156_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__a31o_1
X_08838_ _03446_ _03453_ _03456_ _03459_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_51_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15075__C1 _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12428__A1 _06569_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08769_ net78 net110 VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__xor2_2
XFILLER_0_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_37_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_169_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10800_ _05323_ _05492_ _05493_ _05494_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__a22o_1
XANTENNA__13514__A _04493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11780_ reg_out\[29\] alu_out_q\[29\] _06069_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__mux2_1
XANTENNA__10534__S0 _05235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10731_ _03606_ _03527_ _05388_ _03528_ _03525_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__o311a_1
XFILLER_0_95_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15917__A2 _02617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13928__A1 _03356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13450_ net95 decoded_imm\[6\] VGND VGND VPWR VPWR _07311_ sky130_fd_sc_hd__or2_1
XANTENNA__09057__A0 mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10662_ _05323_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__buf_4
XFILLER_0_165_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14050__B1 _07790_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12401_ cpuregs.regs\[27\]\[4\] _06542_ _06678_ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13381_ net67 decoded_imm\[0\] _07228_ _07245_ VGND VGND VPWR VPWR _07246_ sky130_fd_sc_hd__a31o_1
XANTENNA__12564__S _06763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10593_ _05293_ _05294_ _05295_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15120_ cpuregs.regs\[0\]\[5\] cpuregs.regs\[1\]\[5\] cpuregs.regs\[2\]\[5\] cpuregs.regs\[3\]\[5\]
+ _01973_ _01974_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12332_ cpuregs.regs\[26\]\[4\] _06542_ _06641_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09439__A _04053_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15051_ cpuregs.regs\[8\]\[0\] cpuregs.regs\[9\]\[0\] cpuregs.regs\[10\]\[0\] cpuregs.regs\[11\]\[0\]
+ _03658_ _03659_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12263_ cpuregs.regs\[25\]\[4\] _06542_ _06604_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11167__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14002_ _07767_ _07768_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11214_ _05844_ _05848_ _05851_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__a21oi_1
X_12194_ _06562_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15176__A _03649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput73 net73 VGND VGND VPWR VPWR cpi_rs1[15] sky130_fd_sc_hd__buf_1
X_11145_ _03407_ net126 net103 _04422_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__a22o_2
XANTENNA__15302__B1 _02148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput84 net84 VGND VGND VPWR VPWR cpi_rs1[25] sky130_fd_sc_hd__clkbuf_1
Xoutput95 net95 VGND VGND VPWR VPWR cpi_rs1[6] sky130_fd_sc_hd__clkbuf_1
XANTENNA__14656__A2 _07968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11076_ _03452_ _05736_ _03588_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10127__C1 _04027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15953_ mem_state\[0\] mem_state\[1\] VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__nand2_1
XANTENNA__08547__A_N irq_mask\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09532__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10027_ net41 _04745_ _04666_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__a21o_1
X_14904_ _01826_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10113__A _04272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15884_ instr_lb _02635_ _02636_ is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR _01261_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17623_ clknet_leaf_118_clk _00792_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14835_ count_cycle\[46\] count_cycle\[47\] _01774_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_28_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_106_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13424__A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ clknet_leaf_140_clk _00723_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_14766_ _01729_ _01730_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__nor2_1
X_11978_ _06216_ cpuregs.regs\[21\]\[15\] _06435_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16505_ _02985_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09391__S0 _04123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10929_ _03488_ _05615_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__xor2_1
X_13717_ _05086_ _05227_ VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_152_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14697_ count_cycle\[0\] count_cycle\[1\] count_cycle\[2\] count_cycle\[3\] VGND
+ VGND VPWR VPWR _08340_ sky130_fd_sc_hd__and4_2
X_17485_ clknet_leaf_153_clk _00654_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15464__S0 _01973_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16436_ _06974_ cpuregs.regs\[29\]\[15\] _02943_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__mux2_1
X_13648_ _04959_ _07277_ VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13579_ _07431_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16367_ _02912_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12474__S _06715_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10602__A0 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__16869__A0 _06584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18106_ clknet_leaf_90_clk _01210_ VGND VGND VPWR VPWR timer\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_167_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15318_ _02159_ _02161_ _02164_ _02004_ _01969_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16298_ _02875_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18037_ clknet_leaf_79_clk _00014_ VGND VGND VPWR VPWR irq_pending\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15249_ net130 _02081_ _02098_ _02099_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__o22a_1
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11158__A1 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10366__C1 _03302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15519__S1 _02086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16097__A1 _03747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09810_ _04391_ _04504_ _04505_ _04534_ VGND VGND VPWR VPWR _08371_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_165_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09771__A1 _04017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09741_ net51 _04030_ _04034_ net34 _04423_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__o221a_1
XANTENNA__10669__A0 _04532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09523__A1 _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09523__B2 _03226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09672_ _04398_ _04399_ _04078_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__mux2_1
XANTENNA__10133__A2 _04745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08623_ is_sb_sh_sw _03391_ _03397_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13607__A0 _04708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12649__S _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08554_ irq_mask\[10\] irq_pending\[10\] VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__and2b_2
XFILLER_0_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08428__A _03206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14149__B _07815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08485_ _03254_ _03256_ _03268_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_18_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__16021__A1 decoded_imm\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15455__S0 _01999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09039__A0 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08862__S _03599_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13386__A2 _07250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14583__A1 _08071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12384__S _06663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09106_ _03780_ _03748_ _03743_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__or3b_1
XFILLER_0_115_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_758 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11301__B _05923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09037_ _03794_ _03798_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_92_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09437__S1 _04086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09240__A1_N _03979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16088__A1 is_alu_reg_imm VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12413__A _06677_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15835__A1 decoded_imm_j\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09939_ _04051_ _04659_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__nor2_1
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__15724__A _04737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08948__S0 _03661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12950_ _06987_ cpuregs.regs\[31\]\[21\] _06985_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _06184_ cpuregs.regs\[20\]\[11\] _06398_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12881_ _06940_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10675__A3 _04036_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11832_ _06193_ cpuregs.regs\[11\]\[12\] _06359_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__mux2_1
X_14620_ _08267_ _08271_ VGND VGND VPWR VPWR _08273_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14551_ _07952_ _08206_ VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__and2_1
X_11763_ _06252_ _03341_ _06253_ _06309_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16012__A1 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15446__S0 _01979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16012__B2 mem_rdata_q\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10714_ _05331_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__buf_6
X_13502_ _07304_ _04447_ _07305_ reg_pc\[9\] _07283_ VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17270_ clknet_leaf_125_clk _00444_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_14482_ _07937_ _07992_ _08145_ _06863_ VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14023__B1 _07775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11694_ _06248_ cpuregs.regs\[10\]\[19\] _06176_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13433_ _04342_ _07277_ _07294_ _07279_ VGND VGND VPWR VPWR _07295_ sky130_fd_sc_hd__o211a_1
XANTENNA__11699__A _06065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16221_ net43 mem_16bit_buffer\[3\] _02831_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__mux2_1
XANTENNA__14574__A1 reg_next_pc\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10645_ net72 net73 _05229_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__mux2_1
XANTENNA__12294__S _06615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16152_ net269 net231 _02786_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__mux2_1
X_13364_ _07229_ VGND VGND VPWR VPWR _07230_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10576_ _05255_ _05261_ _05279_ is_compare _03630_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__a32o_1
XANTENNA__09450__B1 _00073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12315_ cpuregs.regs\[25\]\[29\] _06594_ _06626_ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__mux2_1
X_15103_ is_slli_srli_srai cpuregs.raddr2\[2\] decoded_imm\[2\] _01932_ _01934_ VGND
+ VGND VPWR VPWR _01961_ sky130_fd_sc_hd__a221o_1
XANTENNA__10060__B2 _04023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16083_ _03213_ _03833_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__nand2_1
X_13295_ _06982_ cpuregs.regs\[5\]\[19\] _07165_ VGND VGND VPWR VPWR _07175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15034_ irq_mask\[26\] _01865_ _01899_ _01891_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__a211o_1
XFILLER_0_139_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12246_ _06597_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08801__A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08588__B_N decoder_trigger VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16079__A1 decoded_imm\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16079__B2 mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13419__A _07211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12177_ cpuregs.regs\[24\]\[8\] _06550_ _06534_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__mux2_1
XANTENNA__12323__A _06640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10363__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15826__A1 decoded_imm_j\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11128_ _03432_ _05301_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__nand2_1
X_16985_ clknet_leaf_172_clk _00159_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15634__A _07778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11059_ _03455_ _03457_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__or2_1
X_15936_ mem_rdata_q\[16\] mem_rdata_q\[17\] _02660_ _02661_ VGND VGND VPWR VPWR _02662_
+ sky130_fd_sc_hd__or4_1
XANTENNA__08947__S _03709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09600__S1 _04218_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09632__A net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ _02613_ _03940_ _02612_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__and3b_1
XANTENNA__16251__A1 _03864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_17606_ clknet_leaf_18_clk _00775_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_14818_ count_cycle\[40\] _01762_ count_cycle\[41\] VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__a21o_1
X_18586_ clknet_leaf_10_clk _01651_ VGND VGND VPWR VPWR cpuregs.regs\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15798_ latched_compr compressed_instr _08033_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17537_ clknet_leaf_15_clk _00706_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14749_ count_cycle\[19\] _01715_ _01718_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17468_ clknet_leaf_112_clk _00637_ VGND VGND VPWR VPWR cpuregs.regs\[31\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16419_ _06957_ cpuregs.regs\[29\]\[7\] _02932_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__mux2_1
XANTENNA__14565__A1 decoded_imm_j\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17399_ clknet_leaf_121_clk _00568_ VGND VGND VPWR VPWR cpuregs.regs\[9\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15514__B1 _02197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_140_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09807__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08711__A net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11000__A0 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13540__A2 decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__15817__A1 _03892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15817__B2 _03994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09724_ _04010_ _04429_ _04450_ _04150_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__o211a_1
XANTENNA__09542__A _04055_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09655_ irq_mask\[7\] _04308_ timer\[7\] _04023_ _04026_ VGND VGND VPWR VPWR _04384_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08606_ _03382_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__buf_1
X_09586_ _04215_ _04315_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08537_ _03314_ _03315_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12803__A1 _06590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08468_ instr_timer instr_maskirq instr_retirq VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_34_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10430_ _04054_ _05132_ _05136_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08786__A2 _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10361_ _04051_ _05069_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16314__S _02881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11790__A1 _06072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12100_ _06505_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__clkbuf_1
X_13080_ _07061_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10292_ cpuregs.regs\[0\]\[25\] cpuregs.regs\[1\]\[25\] cpuregs.regs\[2\]\[25\] cpuregs.regs\[3\]\[25\]
+ _04217_ _04219_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12031_ _06157_ cpuregs.regs\[22\]\[8\] _06460_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_155_Left_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09830__S1 _04376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11542__B2 _06093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16770_ _03126_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__clkbuf_1
X_13982_ instr_waitirq decoder_trigger VGND VGND VPWR VPWR _07754_ sky130_fd_sc_hd__and2b_2
XFILLER_0_137_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15721_ _02526_ _02527_ _02528_ _02481_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__o211a_1
XANTENNA__09594__S0 _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12933_ _06223_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__buf_2
XANTENNA__10598__A _05213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10502__C1 _04202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10648__A3 _03524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15036__A2 _01865_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18440_ clknet_leaf_151_clk _01505_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_15652_ _02475_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_103_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _06281_ cpuregs.regs\[6\]\[23\] _06928_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14603_ _05941_ _06286_ _07944_ _05922_ VGND VGND VPWR VPWR _08257_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_84_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18371_ clknet_leaf_146_clk _01436_ VGND VGND VPWR VPWR cpuregs.regs\[15\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_11815_ _06125_ cpuregs.regs\[11\]\[4\] _06348_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__mux2_1
XANTENNA_output101_A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12795_ cpuregs.regs\[9\]\[23\] _06582_ _06891_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__mux2_1
X_15583_ cpuregs.regs\[4\]\[29\] cpuregs.regs\[5\]\[29\] cpuregs.regs\[6\]\[29\] cpuregs.regs\[7\]\[29\]
+ _01908_ _01909_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__mux4_1
XFILLER_0_157_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_164_Left_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__15419__S0 _03649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09897__S1 _04376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17322_ clknet_leaf_139_clk _00496_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11746_ _06252_ _03347_ _06253_ _06294_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__a22o_1
X_14534_ _03293_ _07944_ _07946_ _08193_ VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__and4_1
XANTENNA__14517__B _07943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10281__B2 _04165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17253_ clknet_leaf_148_clk _00427_ VGND VGND VPWR VPWR cpuregs.regs\[28\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11677_ _06233_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__clkbuf_1
X_14465_ _08128_ _08129_ VGND VGND VPWR VPWR _08130_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09649__S1 _04376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16204_ prefetched_high_word _02823_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__nor2_1
X_10628_ _05269_ _05271_ _05232_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__mux2_1
X_13416_ _07238_ VGND VGND VPWR VPWR _07279_ sky130_fd_sc_hd__buf_2
XANTENNA__09423__B1 _04156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17184_ clknet_leaf_174_clk _00358_ VGND VGND VPWR VPWR cpuregs.regs\[26\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14396_ _08063_ _08065_ _08066_ _08035_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__o22a_1
X_13347_ _04037_ decoded_imm\[0\] _07213_ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16135_ net292 net128 _02771_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__mux2_1
X_10559_ _03609_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11781__A1 _06252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13278_ _07166_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__clkbuf_1
X_16066_ instr_jal _08232_ _02726_ mem_rdata_q\[31\] VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08531__A cpu_state\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_173_Left_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15017_ _03240_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__clkbuf_4
X_12229_ _06296_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__buf_2
XANTENNA__10336__A2 _05044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12730__A0 _06336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09821__S1 _04087_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09065__C _03822_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15364__A _02066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16968_ clknet_leaf_129_clk _00142_ VGND VGND VPWR VPWR cpuregs.regs\[11\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15919_ _02633_ _02646_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_140_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12199__S _06555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16899_ clknet_leaf_30_clk _00044_ VGND VGND VPWR VPWR mem_rdata_q\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09440_ cpuregs.regs\[20\]\[3\] cpuregs.regs\[21\]\[3\] cpuregs.regs\[22\]\[3\] cpuregs.regs\[23\]\[3\]
+ _04071_ _04073_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__mux4_1
XFILLER_0_91_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09081__B _03237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18638_ clknet_leaf_178_clk _01698_ VGND VGND VPWR VPWR cpuregs.regs\[14\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13038__A1 _06588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14235__B1 _07901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09371_ count_instr\[33\] _04104_ _04105_ count_cycle\[33\] VGND VGND VPWR VPWR _04106_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18569_ clknet_leaf_99_clk _01634_ VGND VGND VPWR VPWR cpuregs.regs\[19\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09662__B1 _04390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10272__B2 _03385_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11772__A1 _06252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09537__A _04009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput230 net230 VGND VGND VPWR VPWR mem_la_wdata[14] sky130_fd_sc_hd__clkbuf_1
XANTENNA__08441__A cpu_state\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput241 net241 VGND VGND VPWR VPWR mem_la_wdata[24] sky130_fd_sc_hd__clkbuf_1
Xoutput252 net252 VGND VGND VPWR VPWR mem_la_wdata[5] sky130_fd_sc_hd__buf_1
Xoutput263 net263 VGND VGND VPWR VPWR mem_wdata[0] sky130_fd_sc_hd__clkbuf_1
Xoutput274 net274 VGND VGND VPWR VPWR mem_wdata[1] sky130_fd_sc_hd__clkbuf_1
Xoutput285 net285 VGND VGND VPWR VPWR mem_wdata[2] sky130_fd_sc_hd__clkbuf_1
Xoutput296 net296 VGND VGND VPWR VPWR mem_wstrb[1] sky130_fd_sc_hd__buf_1
XANTENNA__10910__S _05230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14474__B1 _07905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09272__A _03252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09707_ _04211_ _04433_ _04069_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__o21a_1
XANTENNA__13506__B decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09638_ cpuregs.regs\[8\]\[7\] cpuregs.regs\[9\]\[7\] cpuregs.regs\[10\]\[7\] cpuregs.regs\[11\]\[7\]
+ _04290_ _04276_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__mux4_1
XFILLER_0_167_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09569_ cpuregs.regs\[24\]\[5\] cpuregs.regs\[25\]\[5\] cpuregs.regs\[26\]\[5\] cpuregs.regs\[27\]\[5\]
+ _04275_ _04278_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_65_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12837__S _06917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11600_ _06161_ _06164_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__nor2_2
XFILLER_0_37_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12580_ _06778_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11531_ reg_pc\[2\] _06090_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__xor2_1
XANTENNA__11460__B1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10357__S _04065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11042__A instr_sub VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14250_ _07922_ VGND VGND VPWR VPWR _07942_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11462_ _06041_ irq_pending\[19\] _06049_ net11 VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13201_ _07125_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10413_ count_instr\[61\] _04016_ _04145_ count_instr\[29\] VGND VGND VPWR VPWR _05120_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14181_ _07892_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13752__A2 _05260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11393_ _03633_ _06002_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__nand2_2
XFILLER_0_33_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11763__A1 _06252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10110__S1 _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13132_ _06955_ cpuregs.regs\[4\]\[6\] _07082_ VGND VGND VPWR VPWR _07089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10344_ cpuregs.regs\[28\]\[27\] cpuregs.regs\[29\]\[27\] cpuregs.regs\[30\]\[27\]
+ cpuregs.regs\[31\]\[27\] _04758_ _04759_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14072__B _07815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_303 VGND VGND VPWR VPWR alphacore_303/HI cpi_insn[1] sky130_fd_sc_hd__conb_1
X_17940_ clknet_leaf_67_clk _08381_ VGND VGND VPWR VPWR reg_out\[20\] sky130_fd_sc_hd__dfxtp_1
X_13063_ _07052_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__clkbuf_1
Xalphacore_314 VGND VGND VPWR VPWR alphacore_314/HI cpi_insn[12] sky130_fd_sc_hd__conb_1
X_10275_ reg_pc\[25\] decoded_imm\[25\] VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xalphacore_325 VGND VGND VPWR VPWR alphacore_325/HI cpi_insn[23] sky130_fd_sc_hd__conb_1
XANTENNA__12712__A0 _06266_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xalphacore_336 VGND VGND VPWR VPWR alphacore_336/HI mem_addr[1] sky130_fd_sc_hd__conb_1
X_12014_ _06459_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__clkbuf_8
Xalphacore_347 VGND VGND VPWR VPWR alphacore_347/HI trace_data[8] sky130_fd_sc_hd__conb_1
Xalphacore_358 VGND VGND VPWR VPWR alphacore_358/HI trace_data[19] sky130_fd_sc_hd__conb_1
X_17871_ clknet_leaf_88_clk _01040_ VGND VGND VPWR VPWR count_cycle\[16\] sky130_fd_sc_hd__dfxtp_1
Xalphacore_369 VGND VGND VPWR VPWR alphacore_369/HI trace_data[30] sky130_fd_sc_hd__conb_1
XANTENNA__10105__B decoded_imm\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output149_A net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16822_ _03154_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11279__A0 reg_next_pc\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16753_ _06536_ cpuregs.regs\[13\]\[1\] _03116_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13965_ _07737_ _07742_ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_85_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10177__S1 _04470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15704_ timer\[12\] _02514_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__or2_1
X_12916_ _06963_ cpuregs.regs\[31\]\[10\] _06964_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__mux2_1
X_16684_ _03080_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__clkbuf_1
X_13896_ _07691_ _07694_ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__and2_1
XANTENNA__09910__A _04051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18423_ clknet_leaf_14_clk _01488_ VGND VGND VPWR VPWR cpuregs.regs\[29\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15635_ _02462_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12847_ _06216_ cpuregs.regs\[6\]\[15\] _06917_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__mux2_1
XANTENNA__12747__S _06869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14528__A decoded_imm_j\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13432__A _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18354_ clknet_leaf_53_clk _00061_ VGND VGND VPWR VPWR reg_sh\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15566_ net118 _01905_ _02397_ _02398_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__o22a_1
XANTENNA__13440__A1 _04040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12778_ cpuregs.regs\[9\]\[15\] _06565_ _06880_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10254__A1 _04211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17305_ clknet_leaf_15_clk _00479_ VGND VGND VPWR VPWR cpuregs.regs\[30\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_14517_ decoded_imm_j\[17\] _07943_ VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_155_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18285_ clknet_leaf_42_clk _01353_ VGND VGND VPWR VPWR is_compare sky130_fd_sc_hd__dfxtp_1
X_11729_ _06226_ reg_next_pc\[23\] _06277_ _06279_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__a211o_2
XFILLER_0_83_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15497_ cpuregs.regs\[12\]\[24\] cpuregs.regs\[13\]\[24\] cpuregs.regs\[14\]\[24\]
+ cpuregs.regs\[15\]\[24\] _01970_ _01971_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17236_ clknet_leaf_120_clk _00410_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08960__S _03713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14448_ decoded_imm_j\[12\] _07932_ VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13578__S _07374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17167_ clknet_leaf_124_clk _00341_ VGND VGND VPWR VPWR cpuregs.regs\[25\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14379_ _07986_ _08047_ _08049_ _08050_ _07919_ VGND VGND VPWR VPWR _08051_ sky130_fd_sc_hd__a32o_1
XANTENNA__11754__A1 _06252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16118_ _02776_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17098_ clknet_leaf_139_clk _00272_ VGND VGND VPWR VPWR cpuregs.regs\[23\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08940_ reg_sh\[3\] reg_sh\[2\] reg_sh\[4\] VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__or3b_1
XFILLER_0_0_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_16049_ decoded_imm\[12\] _02720_ _02736_ _02737_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08871_ _03630_ _03632_ _01226_ _03636_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15248__A2 _02009_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09580__C1 _03302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10031__A reg_pc\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09423_ _04152_ _04153_ _04155_ _04156_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__a31o_1
XANTENNA__10493__A1 _04328_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12657__S _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16129__S _02771_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11117__S0 _05286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14438__A decoded_imm_j\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09354_ cpuregs.regs\[0\]\[1\] cpuregs.regs\[1\]\[1\] cpuregs.regs\[2\]\[1\] cpuregs.regs\[3\]\[1\]
+ _04085_ _04087_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__mux4_1
XANTENNA__13431__A1 _04251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10685__B _05260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11442__B1 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09285_ _04021_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_43_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16381__A0 _06987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15184__B2 _02037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11745__A1 alu_out_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16799__S _03138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10060_ irq_mask\[18\] _04021_ timer\[18\] _04023_ _04026_ VGND VGND VPWR VPWR _04778_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__09797__S0 _04325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08799__B_N net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10962_ _03477_ _05398_ _05221_ _03476_ _05646_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__o221a_1
X_13750_ _05044_ _07590_ _07224_ VGND VGND VPWR VPWR _07591_ sky130_fd_sc_hd__mux2_1
XANTENNA__11136__A1_N _04040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_355 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12701_ _06224_ cpuregs.regs\[12\]\[16\] _06836_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10893_ _03491_ _05567_ _03492_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__o21a_1
X_13681_ _07524_ _07525_ VGND VGND VPWR VPWR _07526_ sky130_fd_sc_hd__nand2_1
XANTENNA__15947__B1 _02667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15420_ cpuregs.regs\[16\]\[19\] cpuregs.regs\[17\]\[19\] cpuregs.regs\[18\]\[19\]
+ cpuregs.regs\[19\]\[19\] _03645_ _01991_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_80_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12632_ _06224_ cpuregs.regs\[30\]\[16\] _06799_ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__mux2_1
XANTENNA__13422__B2 reg_pc\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10236__A1 _04391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12563_ _06769_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__clkbuf_1
X_15351_ _02020_ _02187_ _02195_ _01960_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__o211a_4
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_866 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14302_ irq_pending\[12\] irq_pending\[13\] irq_pending\[14\] irq_pending\[15\] VGND
+ VGND VPWR VPWR _07979_ sky130_fd_sc_hd__or4_1
X_11514_ _06087_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__clkbuf_1
X_18070_ clknet_leaf_73_clk _01175_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11203__C _05840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ _06732_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__clkbuf_1
X_15282_ _02129_ _02130_ _02002_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17021_ clknet_leaf_1_clk _00195_ VGND VGND VPWR VPWR cpuregs.regs\[21\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09929__A1 _04231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11445_ irq_mask\[12\] _06030_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__or2_1
X_14233_ reg_pc\[11\] _07926_ _07930_ _07912_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_150_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11736__A1 alu_out_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_706 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11500__A _03195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14164_ count_instr\[55\] count_instr\[54\] count_instr\[53\] _07874_ VGND VGND VPWR
+ VPWR _07881_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_78_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11376_ _05970_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13115_ _07079_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__clkbuf_1
X_10327_ _05024_ _05028_ net301 _05036_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__a211o_4
X_14095_ _07831_ _07832_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__nor2_1
XANTENNA__15907__A mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16502__S _02979_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ cpuregs.regs\[3\]\[30\] _06596_ _07009_ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__mux2_1
X_17923_ clknet_leaf_54_clk _08394_ VGND VGND VPWR VPWR reg_out\[3\] sky130_fd_sc_hd__dfxtp_1
X_10258_ _04214_ _04969_ _04237_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__a21o_1
X_17854_ clknet_leaf_64_clk _01023_ VGND VGND VPWR VPWR reg_next_pc\[31\] sky130_fd_sc_hd__dfxtp_1
X_10189_ cpuregs.regs\[12\]\[22\] cpuregs.regs\[13\]\[22\] cpuregs.regs\[14\]\[22\]
+ cpuregs.regs\[15\]\[22\] _04084_ _04086_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__mux4_1
X_16805_ _06588_ cpuregs.regs\[13\]\[26\] _03138_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__mux2_1
XANTENNA__13336__S1 _04284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17785_ clknet_leaf_85_clk _00954_ VGND VGND VPWR VPWR count_instr\[56\] sky130_fd_sc_hd__dfxtp_1
X_14997_ _04493_ _01869_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09314__C1 _04049_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16736_ _03107_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__clkbuf_1
X_13948_ _03346_ _07727_ _07728_ net144 VGND VGND VPWR VPWR _07731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_46 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09640__A _00071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16667_ cpuregs.regs\[1\]\[28\] _06319_ _03062_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__mux2_1
X_13879_ _03338_ _07678_ _07682_ net131 VGND VGND VPWR VPWR _07683_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18406_ clknet_leaf_140_clk _01471_ VGND VGND VPWR VPWR cpuregs.regs\[16\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15618_ cpuregs.regs\[0\]\[31\] cpuregs.regs\[1\]\[31\] cpuregs.regs\[2\]\[31\] cpuregs.regs\[3\]\[31\]
+ _02046_ _02047_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__mux4_1
XFILLER_0_173_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16598_ _03034_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11424__B1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09712__S0 _04217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18337_ clknet_leaf_35_clk _01405_ VGND VGND VPWR VPWR mem_16bit_buffer\[8\] sky130_fd_sc_hd__dfxtp_1
X_15549_ net117 _02382_ _03272_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10322__S1 _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09070_ mem_16bit_buffer\[8\] _03831_ _03728_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__mux2_1
X_18268_ clknet_leaf_25_clk _01339_ VGND VGND VPWR VPWR decoded_imm\[26\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_114_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15089__A _03666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17219_ clknet_leaf_133_clk _00393_ VGND VGND VPWR VPWR cpuregs.regs\[27\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18199_ clknet_leaf_43_clk _01270_ VGND VGND VPWR VPWR instr_sltiu sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09518__C _03384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10026__A _04668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09972_ _04690_ _04691_ _04121_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__mux2_1
XANTENNA__12940__S _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08923_ _03666_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__buf_6
XANTENNA__11556__S _06086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10460__S _04064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08854_ _03534_ _03493_ _03619_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__and3_1
XANTENNA__12241__A _06327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08785_ net130 net98 VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_146_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09550__A _04280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10466__A1 _04271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10010__S0 _04477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13072__A _07045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09406_ _04138_ _04139_ _04077_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13404__A1 _07232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09608__B1 instr_rdinstr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10218__A1 _04483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09337_ _04071_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__buf_6
XFILLER_0_35_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13800__A _03631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09268_ _03840_ _04001_ _04005_ _03751_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13168__A0 _06991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09199_ _03842_ _03810_ _03845_ _03945_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__a31o_1
XANTENNA__13011__S _07021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08613__B _03387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11230_ _04466_ _03841_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__and2_1
XANTENNA__10077__S0 _04579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__16657__A1 _06280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11161_ _05815_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_2
XFILLER_0_140_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16322__S _02881_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10112_ _04826_ _04827_ _04287_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__mux2_1
X_11092_ _05601_ _05659_ _05767_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_73_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10043_ cpuregs.regs\[20\]\[18\] cpuregs.regs\[21\]\[18\] cpuregs.regs\[22\]\[18\]
+ cpuregs.regs\[23\]\[18\] _04057_ _04060_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__mux4_1
X_14920_ _01834_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12151__A cpuregs.waddr\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10154__B1 _04082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14851_ count_cycle\[52\] _01786_ _01714_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__a21oi_1
X_13802_ _05044_ _05260_ _07614_ VGND VGND VPWR VPWR _07639_ sky130_fd_sc_hd__o21ba_1
X_17570_ clknet_leaf_189_clk _00739_ VGND VGND VPWR VPWR cpuregs.regs\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_14782_ count_cycle\[28\] count_cycle\[29\] count_cycle\[30\] _01736_ VGND VGND VPWR
+ VPWR _01741_ sky130_fd_sc_hd__and4_2
XFILLER_0_97_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11994_ _06449_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14840__B1 _01723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16521_ cpuregs.regs\[17\]\[23\] _06582_ _02990_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__mux2_1
X_13733_ _07304_ _05009_ _07305_ reg_pc\[25\] _07283_ VGND VGND VPWR VPWR _07575_
+ sky130_fd_sc_hd__a221o_1
X_10945_ _03482_ _05630_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12297__S _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16042__C1 _02634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16452_ _02957_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13664_ _04848_ _07271_ _07498_ _07510_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__o22a_1
X_10876_ _05219_ _05553_ _05566_ VGND VGND VPWR VPWR alu_out\[13\] sky130_fd_sc_hd__o21ai_2
XFILLER_0_128_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15403_ cpuregs.regs\[28\]\[18\] cpuregs.regs\[29\]\[18\] cpuregs.regs\[30\]\[18\]
+ cpuregs.regs\[31\]\[18\] _03661_ _03662_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12615_ _06157_ cpuregs.regs\[30\]\[8\] _06788_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__mux2_1
X_16383_ _06989_ cpuregs.regs\[16\]\[22\] _02918_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__mux2_1
X_13595_ net74 decoded_imm\[16\] VGND VGND VPWR VPWR _07446_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_152_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18122_ clknet_leaf_27_clk _01226_ VGND VGND VPWR VPWR decoder_pseudo_trigger sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15334_ _02174_ _02176_ _02179_ _02037_ _02006_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__a221o_1
X_12546_ _06760_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10090__C1 _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15243__S1 _02000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18053_ clknet_leaf_20_clk _01158_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15265_ cpuregs.regs\[16\]\[10\] cpuregs.regs\[17\]\[10\] cpuregs.regs\[18\]\[10\]
+ cpuregs.regs\[19\]\[10\] _01985_ _01986_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12477_ _06723_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11230__A _04466_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17004_ clknet_leaf_180_clk _00178_ VGND VGND VPWR VPWR cpuregs.regs\[20\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_4 _01990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output93_A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14216_ reg_next_pc\[6\] _05834_ _07901_ _07918_ VGND VGND VPWR VPWR _07919_ sky130_fd_sc_hd__o211a_2
XFILLER_0_151_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11428_ _06029_ irq_pending\[3\] _06031_ net26 VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15196_ _03709_ _02048_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__or2_1
XANTENNA__08586__B1 _03308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16648__A1 _06247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14147_ _07865_ _07868_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__and2_1
X_11359_ _05970_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__buf_2
XFILLER_0_67_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15320__A1 decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14078_ count_instr\[29\] _07818_ _07820_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__o21a_1
X_17906_ clknet_leaf_87_clk _01075_ VGND VGND VPWR VPWR count_cycle\[51\] sky130_fd_sc_hd__dfxtp_1
X_13029_ _07034_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13882__A1 _03351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17837_ clknet_leaf_60_clk _01006_ VGND VGND VPWR VPWR reg_next_pc\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15372__A _01932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08570_ irq_mask\[7\] irq_pending\[7\] VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__and2b_2
X_17768_ clknet_leaf_94_clk _00937_ VGND VGND VPWR VPWR count_instr\[39\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__14831__B1 _01723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09370__A instr_rdcycleh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16719_ _06984_ cpuregs.regs\[19\]\[20\] _03098_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09933__S0 _04487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17699_ clknet_leaf_75_clk _00868_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08819__A_N net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15482__S1 _02047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09066__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16407__S _02932_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09122_ _03862_ _03879_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__and2_2
XFILLER_0_115_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15139__A1 _01989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08714__A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09053_ _03810_ _03814_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11176__A2 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13570__B1 _03275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09774__C1 _04499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12670__S _06825_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09545__A _04058_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09955_ irq_pending\[15\] _04049_ _04641_ _03385_ _04675_ VGND VGND VPWR VPWR _08375_
+ sky130_fd_sc_hd__a221o_1
X_08906_ _03646_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__buf_4
XANTENNA__10136__B1 _04851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09886_ _04597_ _04600_ _04607_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10687__A1 _05361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11884__A0 _06114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08837_ _03602_ _03600_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_51_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16378__A _02895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15075__B1 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08768_ _03532_ _03533_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__nand2_2
XANTENNA__15170__S0 _02022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14822__B1 _01723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09280__A instr_rdcycleh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08699_ net111 net79 VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10534__S1 _05237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10730_ _03523_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_24_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10661_ _05300_ _03532_ _05338_ _05355_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__a31o_1
XANTENNA__09057__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12845__S _06917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14626__A _08035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12400_ _06682_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_97_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13380_ net78 decoded_imm\[1\] VGND VGND VPWR VPWR _07245_ sky130_fd_sc_hd__and2_1
X_10592_ _05242_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12331_ _06645_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12262_ _06608_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__clkbuf_1
X_15050_ cpuregs.regs\[12\]\[0\] cpuregs.regs\[13\]\[0\] cpuregs.regs\[14\]\[0\] cpuregs.regs\[15\]\[0\]
+ _01908_ _01909_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11167__A2 _04710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11213_ _05844_ _05848_ _05851_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__and3_1
X_14001_ count_instr\[5\] _07765_ _07759_ VGND VGND VPWR VPWR _07768_ sky130_fd_sc_hd__o21ai_1
X_12193_ cpuregs.regs\[24\]\[13\] _06561_ _06555_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10914__A2 instr_slli VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11144_ _03407_ _05254_ net102 _04422_ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__a22o_2
XANTENNA__15302__A1 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput74 net74 VGND VGND VPWR VPWR cpi_rs1[16] sky130_fd_sc_hd__buf_1
Xoutput85 net85 VGND VGND VPWR VPWR cpi_rs1[26] sky130_fd_sc_hd__buf_1
Xoutput96 net96 VGND VGND VPWR VPWR cpi_rs1[7] sky130_fd_sc_hd__buf_1
X_11075_ _03450_ _05738_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__or2_1
X_15952_ net66 net299 VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__nand2_1
X_10026_ _04668_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__clkbuf_4
X_14903_ net217 net186 _01824_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__mux2_1
XANTENNA__10222__S0 _04280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11209__B _05848_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15883_ _02611_ _02614_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__and2_1
XANTENNA_output229_A net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11924__S _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17622_ clknet_leaf_97_clk _00791_ VGND VGND VPWR VPWR cpuregs.regs\[5\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_14834_ count_cycle\[46\] _01774_ _01776_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__o21a_1
XANTENNA__13616__A1 _04602_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15161__S0 _02013_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14813__B1 _01723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09190__A _03935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13424__B decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17553_ clknet_leaf_136_clk _00722_ VGND VGND VPWR VPWR cpuregs.regs\[4\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ count_cycle\[24\] _01726_ _01723_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_106_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ _06440_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11225__A _04456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16504_ cpuregs.regs\[17\]\[15\] _06565_ _02979_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13716_ _07554_ _07557_ VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_123_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15920__A mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__16566__A0 _06968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10928_ _05517_ _05612_ _03565_ _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__a31o_1
X_17484_ clknet_leaf_160_clk _00653_ VGND VGND VPWR VPWR cpuregs.regs\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09391__S1 _04124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14696_ _08339_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16435_ _02948_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15464__S1 _01974_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13647_ _04810_ _05260_ _07465_ _07279_ VGND VGND VPWR VPWR _07494_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12755__S _06869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10859_ _03498_ _05534_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12052__A0 _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16366_ _06972_ cpuregs.regs\[16\]\[14\] _02907_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__mux2_1
X_13578_ _04611_ _07430_ _07374_ VGND VGND VPWR VPWR _07431_ sky130_fd_sc_hd__mux2_1
XANTENNA__10063__C1 _04780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18105_ clknet_leaf_90_clk _01209_ VGND VGND VPWR VPWR timer\[20\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10602__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15317_ _02162_ _02163_ _02002_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12529_ _06639_ _06750_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__nor2_4
XFILLER_0_14_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16297_ _06972_ cpuregs.regs\[15\]\[14\] _02870_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__mux2_1
X_18036_ clknet_leaf_79_clk _00013_ VGND VGND VPWR VPWR irq_pending\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15248_ decoded_imm\[9\] _02009_ _01963_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12355__A1 _06565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15179_ _01989_ _02032_ _02017_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10905__A2 _05440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09365__A net300 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__16097__A2 _03781_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13304__A0 _06991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09740_ net68 VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__clkbuf_4
.ends

