module simpleuart (clk,
    reg_dat_re,
    reg_dat_wait,
    reg_dat_we,
    resetn,
    ser_rx,
    ser_tx,
    reg_dat_di,
    reg_dat_do,
    reg_div_di,
    reg_div_do,
    reg_div_we);
 input clk;
 input reg_dat_re;
 output reg_dat_wait;
 input reg_dat_we;
 input resetn;
 input ser_rx;
 output ser_tx;
 input [31:0] reg_dat_di;
 output [31:0] reg_dat_do;
 input [31:0] reg_div_di;
 output [31:0] reg_div_do;
 input [3:0] reg_div_we;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire \recv_buf_data[0] ;
 wire \recv_buf_data[1] ;
 wire \recv_buf_data[2] ;
 wire \recv_buf_data[3] ;
 wire \recv_buf_data[4] ;
 wire \recv_buf_data[5] ;
 wire \recv_buf_data[6] ;
 wire \recv_buf_data[7] ;
 wire recv_buf_valid;
 wire \recv_divcnt[0] ;
 wire \recv_divcnt[10] ;
 wire \recv_divcnt[11] ;
 wire \recv_divcnt[12] ;
 wire \recv_divcnt[13] ;
 wire \recv_divcnt[14] ;
 wire \recv_divcnt[15] ;
 wire \recv_divcnt[16] ;
 wire \recv_divcnt[17] ;
 wire \recv_divcnt[18] ;
 wire \recv_divcnt[19] ;
 wire \recv_divcnt[1] ;
 wire \recv_divcnt[20] ;
 wire \recv_divcnt[21] ;
 wire \recv_divcnt[22] ;
 wire \recv_divcnt[23] ;
 wire \recv_divcnt[24] ;
 wire \recv_divcnt[25] ;
 wire \recv_divcnt[26] ;
 wire \recv_divcnt[27] ;
 wire \recv_divcnt[28] ;
 wire \recv_divcnt[29] ;
 wire \recv_divcnt[2] ;
 wire \recv_divcnt[30] ;
 wire \recv_divcnt[31] ;
 wire \recv_divcnt[3] ;
 wire \recv_divcnt[4] ;
 wire \recv_divcnt[5] ;
 wire \recv_divcnt[6] ;
 wire \recv_divcnt[7] ;
 wire \recv_divcnt[8] ;
 wire \recv_divcnt[9] ;
 wire \recv_pattern[0] ;
 wire \recv_pattern[1] ;
 wire \recv_pattern[2] ;
 wire \recv_pattern[3] ;
 wire \recv_pattern[4] ;
 wire \recv_pattern[5] ;
 wire \recv_pattern[6] ;
 wire \recv_pattern[7] ;
 wire \recv_state[0] ;
 wire \recv_state[1] ;
 wire \recv_state[2] ;
 wire \recv_state[3] ;
 wire \send_bitcnt[0] ;
 wire \send_bitcnt[1] ;
 wire \send_bitcnt[2] ;
 wire \send_bitcnt[3] ;
 wire \send_divcnt[0] ;
 wire \send_divcnt[10] ;
 wire \send_divcnt[11] ;
 wire \send_divcnt[12] ;
 wire \send_divcnt[13] ;
 wire \send_divcnt[14] ;
 wire \send_divcnt[15] ;
 wire \send_divcnt[16] ;
 wire \send_divcnt[17] ;
 wire \send_divcnt[18] ;
 wire \send_divcnt[19] ;
 wire \send_divcnt[1] ;
 wire \send_divcnt[20] ;
 wire \send_divcnt[21] ;
 wire \send_divcnt[22] ;
 wire \send_divcnt[23] ;
 wire \send_divcnt[24] ;
 wire \send_divcnt[25] ;
 wire \send_divcnt[26] ;
 wire \send_divcnt[27] ;
 wire \send_divcnt[28] ;
 wire \send_divcnt[29] ;
 wire \send_divcnt[2] ;
 wire \send_divcnt[30] ;
 wire \send_divcnt[31] ;
 wire \send_divcnt[3] ;
 wire \send_divcnt[4] ;
 wire \send_divcnt[5] ;
 wire \send_divcnt[6] ;
 wire \send_divcnt[7] ;
 wire \send_divcnt[8] ;
 wire \send_divcnt[9] ;
 wire send_dummy;
 wire \send_pattern[1] ;
 wire \send_pattern[2] ;
 wire \send_pattern[3] ;
 wire \send_pattern[4] ;
 wire \send_pattern[5] ;
 wire \send_pattern[6] ;
 wire \send_pattern[7] ;
 wire \send_pattern[8] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sky130_fd_sc_hd__or3_2 _0769_ (.A(\send_bitcnt[2] ),
    .B(\send_bitcnt[1] ),
    .C(\send_bitcnt[0] ),
    .X(_0204_));
 sky130_fd_sc_hd__or3_1 _0770_ (.A(send_dummy),
    .B(\send_bitcnt[3] ),
    .C(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__and2_1 _0771_ (.A(net10),
    .B(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__clkbuf_1 _0772_ (.A(_0206_),
    .X(net81));
 sky130_fd_sc_hd__clkinv_8 _0773_ (.A(recv_buf_valid),
    .Y(net73));
 sky130_fd_sc_hd__or2_1 _0774_ (.A(\recv_buf_data[0] ),
    .B(net73),
    .X(_0207_));
 sky130_fd_sc_hd__clkbuf_1 _0775_ (.A(_0207_),
    .X(net49));
 sky130_fd_sc_hd__or2_1 _0776_ (.A(\recv_buf_data[1] ),
    .B(net73),
    .X(_0208_));
 sky130_fd_sc_hd__clkbuf_1 _0777_ (.A(_0208_),
    .X(net60));
 sky130_fd_sc_hd__or2_1 _0778_ (.A(\recv_buf_data[2] ),
    .B(net73),
    .X(_0209_));
 sky130_fd_sc_hd__clkbuf_1 _0779_ (.A(_0209_),
    .X(net71));
 sky130_fd_sc_hd__or2_1 _0780_ (.A(\recv_buf_data[3] ),
    .B(net73),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_1 _0781_ (.A(_0210_),
    .X(net74));
 sky130_fd_sc_hd__or2_1 _0782_ (.A(\recv_buf_data[4] ),
    .B(net73),
    .X(_0211_));
 sky130_fd_sc_hd__clkbuf_1 _0783_ (.A(_0211_),
    .X(net75));
 sky130_fd_sc_hd__or2_1 _0784_ (.A(\recv_buf_data[5] ),
    .B(net73),
    .X(_0212_));
 sky130_fd_sc_hd__clkbuf_1 _0785_ (.A(_0212_),
    .X(net76));
 sky130_fd_sc_hd__or2_1 _0786_ (.A(\recv_buf_data[6] ),
    .B(net73),
    .X(_0213_));
 sky130_fd_sc_hd__clkbuf_1 _0787_ (.A(_0213_),
    .X(net77));
 sky130_fd_sc_hd__or2_1 _0788_ (.A(\recv_buf_data[7] ),
    .B(net73),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_1 _0789_ (.A(_0214_),
    .X(net78));
 sky130_fd_sc_hd__nor2_1 _0790_ (.A(net73),
    .B(net9),
    .Y(_0215_));
 sky130_fd_sc_hd__inv_2 _0791_ (.A(\recv_state[3] ),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_2 _0792_ (.A(\recv_state[1] ),
    .Y(_0217_));
 sky130_fd_sc_hd__or4_1 _0793_ (.A(_0216_),
    .B(\recv_state[2] ),
    .C(_0217_),
    .D(\recv_state[0] ),
    .X(_0218_));
 sky130_fd_sc_hd__clkbuf_4 _0794_ (.A(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__inv_2 _0795_ (.A(\recv_divcnt[29] ),
    .Y(_0220_));
 sky130_fd_sc_hd__xor2_1 _0796_ (.A(net105),
    .B(\recv_divcnt[30] ),
    .X(_0221_));
 sky130_fd_sc_hd__inv_2 _0797_ (.A(net106),
    .Y(_0222_));
 sky130_fd_sc_hd__and2_1 _0798_ (.A(_0222_),
    .B(\recv_divcnt[31] ),
    .X(_0223_));
 sky130_fd_sc_hd__nor2_1 _0799_ (.A(_0222_),
    .B(\recv_divcnt[31] ),
    .Y(_0224_));
 sky130_fd_sc_hd__a2111o_1 _0800_ (.A1(net103),
    .A2(_0220_),
    .B1(_0221_),
    .C1(_0223_),
    .D1(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__inv_2 _0801_ (.A(\recv_divcnt[28] ),
    .Y(_0226_));
 sky130_fd_sc_hd__o22a_1 _0802_ (.A1(net103),
    .A2(_0220_),
    .B1(_0226_),
    .B2(net102),
    .X(_0227_));
 sky130_fd_sc_hd__or2_1 _0803_ (.A(_0225_),
    .B(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__inv_2 _0804_ (.A(net111),
    .Y(_0229_));
 sky130_fd_sc_hd__nand2_1 _0805_ (.A(_0229_),
    .B(\recv_divcnt[7] ),
    .Y(_0230_));
 sky130_fd_sc_hd__inv_2 _0806_ (.A(net109),
    .Y(_0231_));
 sky130_fd_sc_hd__inv_2 _0807_ (.A(net108),
    .Y(_0232_));
 sky130_fd_sc_hd__a22o_1 _0808_ (.A1(_0231_),
    .A2(\recv_divcnt[5] ),
    .B1(\recv_divcnt[4] ),
    .B2(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__inv_2 _0809_ (.A(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _0810_ (.A(net107),
    .Y(_0235_));
 sky130_fd_sc_hd__inv_2 _0811_ (.A(net104),
    .Y(_0236_));
 sky130_fd_sc_hd__a22o_1 _0812_ (.A1(_0235_),
    .A2(\recv_divcnt[3] ),
    .B1(\recv_divcnt[2] ),
    .B2(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__inv_2 _0813_ (.A(net93),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_2 _0814_ (.A(net82),
    .Y(_0239_));
 sky130_fd_sc_hd__o22a_1 _0815_ (.A1(_0238_),
    .A2(\recv_divcnt[1] ),
    .B1(\recv_divcnt[0] ),
    .B2(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__and2_1 _0816_ (.A(_0238_),
    .B(\recv_divcnt[1] ),
    .X(_0241_));
 sky130_fd_sc_hd__o22a_1 _0817_ (.A1(_0236_),
    .A2(\recv_divcnt[2] ),
    .B1(_0240_),
    .B2(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__o22a_1 _0818_ (.A1(_0232_),
    .A2(\recv_divcnt[4] ),
    .B1(\recv_divcnt[3] ),
    .B2(_0235_),
    .X(_0243_));
 sky130_fd_sc_hd__o21ai_1 _0819_ (.A1(_0237_),
    .A2(_0242_),
    .B1(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__nor2_1 _0820_ (.A(_0231_),
    .B(\recv_divcnt[5] ),
    .Y(_0245_));
 sky130_fd_sc_hd__clkinv_2 _0821_ (.A(net110),
    .Y(_0246_));
 sky130_fd_sc_hd__inv_2 _0822_ (.A(\recv_divcnt[6] ),
    .Y(_0247_));
 sky130_fd_sc_hd__nor2_1 _0823_ (.A(_0229_),
    .B(\recv_divcnt[7] ),
    .Y(_0248_));
 sky130_fd_sc_hd__a21o_1 _0824_ (.A1(net110),
    .A2(_0247_),
    .B1(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__a21o_1 _0825_ (.A1(_0246_),
    .A2(\recv_divcnt[6] ),
    .B1(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__a211o_1 _0826_ (.A1(_0234_),
    .A2(_0244_),
    .B1(_0245_),
    .C1(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__or3_1 _0827_ (.A(net110),
    .B(_0247_),
    .C(_0248_),
    .X(_0252_));
 sky130_fd_sc_hd__inv_2 _0828_ (.A(net88),
    .Y(_0253_));
 sky130_fd_sc_hd__inv_2 _0829_ (.A(\recv_divcnt[14] ),
    .Y(_0254_));
 sky130_fd_sc_hd__nor2_1 _0830_ (.A(net87),
    .B(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__a21o_1 _0831_ (.A1(_0253_),
    .A2(\recv_divcnt[15] ),
    .B1(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__inv_2 _0832_ (.A(net86),
    .Y(_0257_));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(net85),
    .Y(_0258_));
 sky130_fd_sc_hd__a22o_1 _0834_ (.A1(_0257_),
    .A2(\recv_divcnt[13] ),
    .B1(\recv_divcnt[12] ),
    .B2(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__inv_2 _0835_ (.A(\recv_divcnt[9] ),
    .Y(_0260_));
 sky130_fd_sc_hd__inv_2 _0836_ (.A(\recv_divcnt[8] ),
    .Y(_0261_));
 sky130_fd_sc_hd__o22a_1 _0837_ (.A1(net113),
    .A2(_0260_),
    .B1(_0261_),
    .B2(net112),
    .X(_0262_));
 sky130_fd_sc_hd__or3b_1 _0838_ (.A(_0256_),
    .B(_0259_),
    .C_N(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__inv_2 _0839_ (.A(\recv_divcnt[13] ),
    .Y(_0264_));
 sky130_fd_sc_hd__or2_1 _0840_ (.A(_0253_),
    .B(\recv_divcnt[15] ),
    .X(_0265_));
 sky130_fd_sc_hd__inv_2 _0841_ (.A(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__a221o_1 _0842_ (.A1(net87),
    .A2(_0254_),
    .B1(_0264_),
    .B2(net86),
    .C1(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__inv_2 _0843_ (.A(net83),
    .Y(_0268_));
 sky130_fd_sc_hd__a2bb2o_1 _0844_ (.A1_N(_0268_),
    .A2_N(\recv_divcnt[10] ),
    .B1(_0260_),
    .B2(net113),
    .X(_0269_));
 sky130_fd_sc_hd__inv_2 _0845_ (.A(net84),
    .Y(_0270_));
 sky130_fd_sc_hd__nor2_1 _0846_ (.A(_0270_),
    .B(\recv_divcnt[11] ),
    .Y(_0271_));
 sky130_fd_sc_hd__a211o_1 _0847_ (.A1(_0268_),
    .A2(\recv_divcnt[10] ),
    .B1(_0269_),
    .C1(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__nor2_1 _0848_ (.A(_0258_),
    .B(\recv_divcnt[12] ),
    .Y(_0273_));
 sky130_fd_sc_hd__a221o_1 _0849_ (.A1(_0270_),
    .A2(\recv_divcnt[11] ),
    .B1(_0261_),
    .B2(net112),
    .C1(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__or4_1 _0850_ (.A(_0263_),
    .B(_0267_),
    .C(_0272_),
    .D(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__a31o_1 _0851_ (.A1(_0230_),
    .A2(_0251_),
    .A3(_0252_),
    .B1(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__inv_2 _0852_ (.A(\recv_divcnt[11] ),
    .Y(_0277_));
 sky130_fd_sc_hd__or3b_1 _0853_ (.A(net83),
    .B(_0271_),
    .C_N(\recv_divcnt[10] ),
    .X(_0278_));
 sky130_fd_sc_hd__o221a_1 _0854_ (.A1(net84),
    .A2(_0277_),
    .B1(_0262_),
    .B2(_0272_),
    .C1(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__o21ba_1 _0855_ (.A1(_0273_),
    .A2(_0279_),
    .B1_N(_0259_),
    .X(_0280_));
 sky130_fd_sc_hd__or3_1 _0856_ (.A(_0255_),
    .B(_0267_),
    .C(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__nand2_1 _0857_ (.A(_0256_),
    .B(_0265_),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _0858_ (.A(net102),
    .Y(_0283_));
 sky130_fd_sc_hd__nor2_1 _0859_ (.A(_0283_),
    .B(\recv_divcnt[28] ),
    .Y(_0284_));
 sky130_fd_sc_hd__or3b_1 _0860_ (.A(_0225_),
    .B(_0284_),
    .C_N(_0227_),
    .X(_0285_));
 sky130_fd_sc_hd__inv_2 _0861_ (.A(net100),
    .Y(_0286_));
 sky130_fd_sc_hd__and2_1 _0862_ (.A(_0286_),
    .B(\recv_divcnt[26] ),
    .X(_0287_));
 sky130_fd_sc_hd__clkinv_2 _0863_ (.A(net101),
    .Y(_0288_));
 sky130_fd_sc_hd__nor2_1 _0864_ (.A(_0288_),
    .B(\recv_divcnt[27] ),
    .Y(_0289_));
 sky130_fd_sc_hd__inv_2 _0865_ (.A(net99),
    .Y(_0290_));
 sky130_fd_sc_hd__nand2_1 _0866_ (.A(_0288_),
    .B(\recv_divcnt[27] ),
    .Y(_0291_));
 sky130_fd_sc_hd__o221a_1 _0867_ (.A1(_0286_),
    .A2(\recv_divcnt[26] ),
    .B1(\recv_divcnt[25] ),
    .B2(_0290_),
    .C1(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__or3b_1 _0868_ (.A(_0287_),
    .B(_0289_),
    .C_N(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__inv_2 _0869_ (.A(net98),
    .Y(_0294_));
 sky130_fd_sc_hd__nor2_1 _0870_ (.A(_0294_),
    .B(\recv_divcnt[24] ),
    .Y(_0295_));
 sky130_fd_sc_hd__inv_2 _0871_ (.A(\recv_divcnt[25] ),
    .Y(_0296_));
 sky130_fd_sc_hd__inv_2 _0872_ (.A(\recv_divcnt[24] ),
    .Y(_0297_));
 sky130_fd_sc_hd__o22a_1 _0873_ (.A1(net99),
    .A2(_0296_),
    .B1(_0297_),
    .B2(net98),
    .X(_0298_));
 sky130_fd_sc_hd__or4b_1 _0874_ (.A(_0285_),
    .B(_0293_),
    .C(_0295_),
    .D_N(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__inv_2 _0875_ (.A(net89),
    .Y(_0300_));
 sky130_fd_sc_hd__clkinv_2 _0876_ (.A(\recv_divcnt[17] ),
    .Y(_0301_));
 sky130_fd_sc_hd__inv_2 _0877_ (.A(\recv_divcnt[16] ),
    .Y(_0302_));
 sky130_fd_sc_hd__o22a_1 _0878_ (.A1(net90),
    .A2(_0301_),
    .B1(_0302_),
    .B2(net89),
    .X(_0303_));
 sky130_fd_sc_hd__inv_2 _0879_ (.A(\recv_divcnt[20] ),
    .Y(_0304_));
 sky130_fd_sc_hd__inv_2 _0880_ (.A(\recv_divcnt[19] ),
    .Y(_0305_));
 sky130_fd_sc_hd__o22a_1 _0881_ (.A1(net94),
    .A2(_0304_),
    .B1(_0305_),
    .B2(net92),
    .X(_0306_));
 sky130_fd_sc_hd__nand2_1 _0882_ (.A(net90),
    .B(_0301_),
    .Y(_0307_));
 sky130_fd_sc_hd__o2111ai_1 _0883_ (.A1(_0300_),
    .A2(\recv_divcnt[16] ),
    .B1(_0303_),
    .C1(_0306_),
    .D1(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__and2b_1 _0884_ (.A_N(\recv_divcnt[19] ),
    .B(net92),
    .X(_0309_));
 sky130_fd_sc_hd__xor2_1 _0885_ (.A(net91),
    .B(\recv_divcnt[18] ),
    .X(_0310_));
 sky130_fd_sc_hd__or2_1 _0886_ (.A(_0309_),
    .B(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__inv_2 _0887_ (.A(\recv_divcnt[22] ),
    .Y(_0312_));
 sky130_fd_sc_hd__clkinv_2 _0888_ (.A(net97),
    .Y(_0313_));
 sky130_fd_sc_hd__nor2_1 _0889_ (.A(_0313_),
    .B(\recv_divcnt[23] ),
    .Y(_0314_));
 sky130_fd_sc_hd__clkinv_2 _0890_ (.A(net96),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_2 _0891_ (.A(\recv_divcnt[21] ),
    .Y(_0316_));
 sky130_fd_sc_hd__a22o_1 _0892_ (.A1(_0315_),
    .A2(\recv_divcnt[22] ),
    .B1(_0316_),
    .B2(net95),
    .X(_0317_));
 sky130_fd_sc_hd__a211o_1 _0893_ (.A1(net96),
    .A2(_0312_),
    .B1(_0314_),
    .C1(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__clkinv_2 _0894_ (.A(net95),
    .Y(_0319_));
 sky130_fd_sc_hd__clkinv_2 _0895_ (.A(net94),
    .Y(_0320_));
 sky130_fd_sc_hd__nor2_1 _0896_ (.A(_0320_),
    .B(\recv_divcnt[20] ),
    .Y(_0321_));
 sky130_fd_sc_hd__a221o_1 _0897_ (.A1(_0313_),
    .A2(\recv_divcnt[23] ),
    .B1(\recv_divcnt[21] ),
    .B2(_0319_),
    .C1(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__or3_1 _0898_ (.A(_0311_),
    .B(_0318_),
    .C(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__or3_1 _0899_ (.A(_0299_),
    .B(_0308_),
    .C(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__a31o_1 _0900_ (.A1(_0276_),
    .A2(_0281_),
    .A3(_0282_),
    .B1(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__or2b_1 _0901_ (.A(_0289_),
    .B_N(_0287_),
    .X(_0326_));
 sky130_fd_sc_hd__o211a_1 _0902_ (.A1(_0293_),
    .A2(_0298_),
    .B1(_0326_),
    .C1(_0291_),
    .X(_0327_));
 sky130_fd_sc_hd__inv_2 _0903_ (.A(\recv_divcnt[23] ),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _0904_ (.A(\recv_divcnt[18] ),
    .Y(_0329_));
 sky130_fd_sc_hd__or3b_1 _0905_ (.A(_0303_),
    .B(_0311_),
    .C_N(_0307_),
    .X(_0330_));
 sky130_fd_sc_hd__o311a_1 _0906_ (.A1(net91),
    .A2(_0329_),
    .A3(_0309_),
    .B1(_0330_),
    .C1(_0306_),
    .X(_0331_));
 sky130_fd_sc_hd__o22a_1 _0907_ (.A1(net95),
    .A2(_0316_),
    .B1(_0321_),
    .B2(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__or3_1 _0908_ (.A(net96),
    .B(_0312_),
    .C(_0314_),
    .X(_0333_));
 sky130_fd_sc_hd__o221a_1 _0909_ (.A1(net97),
    .A2(_0328_),
    .B1(_0318_),
    .B2(_0332_),
    .C1(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__inv_2 _0910_ (.A(net105),
    .Y(_0335_));
 sky130_fd_sc_hd__inv_2 _0911_ (.A(\recv_divcnt[30] ),
    .Y(_0336_));
 sky130_fd_sc_hd__nor2_1 _0912_ (.A(_0336_),
    .B(_0224_),
    .Y(_0337_));
 sky130_fd_sc_hd__a21oi_1 _0913_ (.A1(_0335_),
    .A2(_0337_),
    .B1(_0223_),
    .Y(_0338_));
 sky130_fd_sc_hd__o221a_1 _0914_ (.A1(_0285_),
    .A2(_0327_),
    .B1(_0334_),
    .B2(_0299_),
    .C1(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__nand2_1 _0915_ (.A(_0240_),
    .B(_0243_),
    .Y(_0340_));
 sky130_fd_sc_hd__inv_2 _0916_ (.A(\recv_divcnt[2] ),
    .Y(_0341_));
 sky130_fd_sc_hd__a221o_1 _0917_ (.A1(_0229_),
    .A2(\recv_divcnt[7] ),
    .B1(\recv_divcnt[0] ),
    .B2(_0239_),
    .C1(_0241_),
    .X(_0342_));
 sky130_fd_sc_hd__a2111o_1 _0918_ (.A1(net104),
    .A2(_0341_),
    .B1(_0342_),
    .C1(_0237_),
    .D1(_0245_),
    .X(_0343_));
 sky130_fd_sc_hd__or4_1 _0919_ (.A(_0233_),
    .B(_0340_),
    .C(_0250_),
    .D(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__nor3_1 _0920_ (.A(_0344_),
    .B(_0275_),
    .C(_0324_),
    .Y(_0345_));
 sky130_fd_sc_hd__a31o_1 _0921_ (.A1(_0228_),
    .A2(_0325_),
    .A3(_0339_),
    .B1(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_4 _0922_ (.A(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__nor2_4 _0923_ (.A(_0219_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__buf_4 _0924_ (.A(net47),
    .X(_0349_));
 sky130_fd_sc_hd__clkbuf_4 _0925_ (.A(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__o21a_1 _0926_ (.A1(_0215_),
    .A2(_0348_),
    .B1(_0350_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_4 _0927_ (.A(_0349_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _0928_ (.A0(net112),
    .A1(net41),
    .S(net44),
    .X(_0352_));
 sky130_fd_sc_hd__and2_1 _0929_ (.A(_0351_),
    .B(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_1 _0930_ (.A(_0353_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _0931_ (.A0(net113),
    .A1(net42),
    .S(net44),
    .X(_0354_));
 sky130_fd_sc_hd__and2_1 _0932_ (.A(_0351_),
    .B(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _0933_ (.A(_0355_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _0934_ (.A0(net83),
    .A1(net12),
    .S(net44),
    .X(_0356_));
 sky130_fd_sc_hd__and2_1 _0935_ (.A(_0351_),
    .B(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_1 _0936_ (.A(_0357_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _0937_ (.A0(net84),
    .A1(net13),
    .S(net44),
    .X(_0358_));
 sky130_fd_sc_hd__and2_1 _0938_ (.A(_0351_),
    .B(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_1 _0939_ (.A(_0359_),
    .X(_0004_));
 sky130_fd_sc_hd__clkbuf_2 _0940_ (.A(_0349_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _0941_ (.A0(net85),
    .A1(net14),
    .S(net44),
    .X(_0361_));
 sky130_fd_sc_hd__and2_1 _0942_ (.A(_0360_),
    .B(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_1 _0943_ (.A(_0362_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _0944_ (.A0(net86),
    .A1(net15),
    .S(net44),
    .X(_0363_));
 sky130_fd_sc_hd__and2_1 _0945_ (.A(_0360_),
    .B(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_1 _0946_ (.A(_0364_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _0947_ (.A0(net87),
    .A1(net16),
    .S(net44),
    .X(_0365_));
 sky130_fd_sc_hd__and2_1 _0948_ (.A(_0360_),
    .B(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_1 _0949_ (.A(_0366_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _0950_ (.A0(net88),
    .A1(net17),
    .S(net44),
    .X(_0367_));
 sky130_fd_sc_hd__and2_1 _0951_ (.A(_0360_),
    .B(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_1 _0952_ (.A(_0368_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _0953_ (.A0(net89),
    .A1(net18),
    .S(net45),
    .X(_0369_));
 sky130_fd_sc_hd__and2_1 _0954_ (.A(_0360_),
    .B(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_1 _0955_ (.A(_0370_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(net90),
    .A1(net19),
    .S(net45),
    .X(_0371_));
 sky130_fd_sc_hd__and2_1 _0957_ (.A(_0360_),
    .B(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__clkbuf_1 _0958_ (.A(_0372_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _0959_ (.A0(net91),
    .A1(net20),
    .S(net45),
    .X(_0373_));
 sky130_fd_sc_hd__and2_1 _0960_ (.A(_0360_),
    .B(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _0961_ (.A(_0374_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _0962_ (.A0(net92),
    .A1(net21),
    .S(net45),
    .X(_0375_));
 sky130_fd_sc_hd__and2_1 _0963_ (.A(_0360_),
    .B(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_1 _0964_ (.A(_0376_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _0965_ (.A0(net94),
    .A1(net23),
    .S(net45),
    .X(_0377_));
 sky130_fd_sc_hd__and2_1 _0966_ (.A(_0360_),
    .B(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_1 _0967_ (.A(_0378_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _0968_ (.A0(net95),
    .A1(net24),
    .S(net45),
    .X(_0379_));
 sky130_fd_sc_hd__and2_1 _0969_ (.A(_0360_),
    .B(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _0970_ (.A(_0380_),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_2 _0971_ (.A(net47),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _0972_ (.A0(net96),
    .A1(net25),
    .S(net45),
    .X(_0382_));
 sky130_fd_sc_hd__and2_1 _0973_ (.A(_0381_),
    .B(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_1 _0974_ (.A(_0383_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _0975_ (.A0(net97),
    .A1(net26),
    .S(net45),
    .X(_0384_));
 sky130_fd_sc_hd__and2_1 _0976_ (.A(_0381_),
    .B(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_1 _0977_ (.A(_0385_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0978_ (.A0(net98),
    .A1(net27),
    .S(net46),
    .X(_0386_));
 sky130_fd_sc_hd__and2_1 _0979_ (.A(_0381_),
    .B(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_1 _0980_ (.A(_0387_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _0981_ (.A0(net99),
    .A1(net28),
    .S(net46),
    .X(_0388_));
 sky130_fd_sc_hd__and2_1 _0982_ (.A(_0381_),
    .B(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_1 _0983_ (.A(_0389_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0984_ (.A0(net100),
    .A1(net29),
    .S(net46),
    .X(_0390_));
 sky130_fd_sc_hd__and2_1 _0985_ (.A(_0381_),
    .B(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_1 _0986_ (.A(_0391_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0987_ (.A0(net101),
    .A1(net30),
    .S(net46),
    .X(_0392_));
 sky130_fd_sc_hd__and2_1 _0988_ (.A(_0381_),
    .B(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _0989_ (.A(_0393_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _0990_ (.A0(net102),
    .A1(net31),
    .S(net46),
    .X(_0394_));
 sky130_fd_sc_hd__and2_1 _0991_ (.A(_0381_),
    .B(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _0992_ (.A(_0395_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _0993_ (.A0(net103),
    .A1(net32),
    .S(net46),
    .X(_0396_));
 sky130_fd_sc_hd__and2_1 _0994_ (.A(_0381_),
    .B(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_1 _0995_ (.A(_0397_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(net105),
    .A1(net34),
    .S(net46),
    .X(_0398_));
 sky130_fd_sc_hd__and2_1 _0997_ (.A(_0381_),
    .B(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_1 _0998_ (.A(_0399_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _0999_ (.A0(net106),
    .A1(net35),
    .S(net46),
    .X(_0400_));
 sky130_fd_sc_hd__and2_1 _1000_ (.A(_0381_),
    .B(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _1001_ (.A(_0401_),
    .X(_0024_));
 sky130_fd_sc_hd__o22a_1 _1002_ (.A1(_0313_),
    .A2(\send_divcnt[23] ),
    .B1(\send_divcnt[22] ),
    .B2(_0315_),
    .X(_0402_));
 sky130_fd_sc_hd__inv_2 _1003_ (.A(\send_divcnt[13] ),
    .Y(_0403_));
 sky130_fd_sc_hd__a2bb2o_1 _1004_ (.A1_N(\send_divcnt[12] ),
    .A2_N(_0258_),
    .B1(net86),
    .B2(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__inv_2 _1005_ (.A(\send_divcnt[14] ),
    .Y(_0405_));
 sky130_fd_sc_hd__o22a_1 _1006_ (.A1(net87),
    .A2(_0405_),
    .B1(_0403_),
    .B2(net86),
    .X(_0406_));
 sky130_fd_sc_hd__and2b_1 _1007_ (.A_N(_0404_),
    .B(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__inv_2 _1008_ (.A(\send_divcnt[10] ),
    .Y(_0408_));
 sky130_fd_sc_hd__a2bb2o_1 _1009_ (.A1_N(_0270_),
    .A2_N(\send_divcnt[11] ),
    .B1(_0408_),
    .B2(net83),
    .X(_0409_));
 sky130_fd_sc_hd__or2b_1 _1010_ (.A(net84),
    .B_N(\send_divcnt[11] ),
    .X(_0410_));
 sky130_fd_sc_hd__inv_2 _1011_ (.A(\send_divcnt[8] ),
    .Y(_0411_));
 sky130_fd_sc_hd__inv_2 _1012_ (.A(\send_divcnt[7] ),
    .Y(_0412_));
 sky130_fd_sc_hd__inv_2 _1013_ (.A(\send_divcnt[9] ),
    .Y(_0413_));
 sky130_fd_sc_hd__a22o_1 _1014_ (.A1(net113),
    .A2(_0413_),
    .B1(_0411_),
    .B2(net112),
    .X(_0414_));
 sky130_fd_sc_hd__inv_2 _1015_ (.A(net113),
    .Y(_0415_));
 sky130_fd_sc_hd__o21ai_1 _1016_ (.A1(net83),
    .A2(_0408_),
    .B1(_0410_),
    .Y(_0416_));
 sky130_fd_sc_hd__a211o_1 _1017_ (.A1(_0415_),
    .A2(\send_divcnt[9] ),
    .B1(_0409_),
    .C1(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__nor2_1 _1018_ (.A(_0414_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__o221a_1 _1019_ (.A1(net112),
    .A2(_0411_),
    .B1(_0412_),
    .B2(net111),
    .C1(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__nand2_1 _1020_ (.A(_0246_),
    .B(\send_divcnt[6] ),
    .Y(_0420_));
 sky130_fd_sc_hd__inv_2 _1021_ (.A(\send_divcnt[5] ),
    .Y(_0421_));
 sky130_fd_sc_hd__and2b_1 _1022_ (.A_N(net93),
    .B(\send_divcnt[1] ),
    .X(_0422_));
 sky130_fd_sc_hd__and2b_1 _1023_ (.A_N(net82),
    .B(\send_divcnt[0] ),
    .X(_0423_));
 sky130_fd_sc_hd__or2b_1 _1024_ (.A(\send_divcnt[1] ),
    .B_N(net93),
    .X(_0424_));
 sky130_fd_sc_hd__o221a_1 _1025_ (.A1(_0236_),
    .A2(\send_divcnt[2] ),
    .B1(_0422_),
    .B2(_0423_),
    .C1(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_1 _1026_ (.A1(_0235_),
    .A2(\send_divcnt[3] ),
    .B1(\send_divcnt[2] ),
    .B2(_0236_),
    .X(_0426_));
 sky130_fd_sc_hd__o22a_1 _1027_ (.A1(_0232_),
    .A2(\send_divcnt[4] ),
    .B1(\send_divcnt[3] ),
    .B2(_0235_),
    .X(_0427_));
 sky130_fd_sc_hd__o21ai_1 _1028_ (.A1(_0425_),
    .A2(_0426_),
    .B1(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__inv_2 _1029_ (.A(\send_divcnt[4] ),
    .Y(_0429_));
 sky130_fd_sc_hd__o22a_1 _1030_ (.A1(net109),
    .A2(_0421_),
    .B1(_0429_),
    .B2(net108),
    .X(_0430_));
 sky130_fd_sc_hd__nor2_1 _1031_ (.A(_0246_),
    .B(\send_divcnt[6] ),
    .Y(_0431_));
 sky130_fd_sc_hd__a221o_1 _1032_ (.A1(net109),
    .A2(_0421_),
    .B1(_0428_),
    .B2(_0430_),
    .C1(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__a22o_1 _1033_ (.A1(net111),
    .A2(_0412_),
    .B1(_0420_),
    .B2(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__and2b_1 _1034_ (.A_N(_0417_),
    .B(_0414_),
    .X(_0434_));
 sky130_fd_sc_hd__a221o_1 _1035_ (.A1(_0409_),
    .A2(_0410_),
    .B1(_0419_),
    .B2(_0433_),
    .C1(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__inv_2 _1036_ (.A(\send_divcnt[15] ),
    .Y(_0436_));
 sky130_fd_sc_hd__a22o_1 _1037_ (.A1(net88),
    .A2(_0436_),
    .B1(_0405_),
    .B2(net87),
    .X(_0437_));
 sky130_fd_sc_hd__nor2_1 _1038_ (.A(net88),
    .B(_0436_),
    .Y(_0438_));
 sky130_fd_sc_hd__a211oi_1 _1039_ (.A1(_0258_),
    .A2(\send_divcnt[12] ),
    .B1(_0437_),
    .C1(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__a21oi_1 _1040_ (.A1(_0404_),
    .A2(_0406_),
    .B1(_0437_),
    .Y(_0440_));
 sky130_fd_sc_hd__nor2_1 _1041_ (.A(_0438_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__a31o_1 _1042_ (.A1(_0407_),
    .A2(_0435_),
    .A3(_0439_),
    .B1(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__inv_2 _1043_ (.A(\send_divcnt[17] ),
    .Y(_0443_));
 sky130_fd_sc_hd__nor2_1 _1044_ (.A(net90),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__and2_1 _1045_ (.A(_0320_),
    .B(\send_divcnt[20] ),
    .X(_0445_));
 sky130_fd_sc_hd__nor2_1 _1046_ (.A(_0444_),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__xnor2_1 _1047_ (.A(net89),
    .B(\send_divcnt[16] ),
    .Y(_0447_));
 sky130_fd_sc_hd__nand2_1 _1048_ (.A(_0313_),
    .B(\send_divcnt[23] ),
    .Y(_0448_));
 sky130_fd_sc_hd__a22oi_1 _1049_ (.A1(_0315_),
    .A2(\send_divcnt[22] ),
    .B1(\send_divcnt[21] ),
    .B2(_0319_),
    .Y(_0449_));
 sky130_fd_sc_hd__o211a_1 _1050_ (.A1(_0319_),
    .A2(\send_divcnt[21] ),
    .B1(_0448_),
    .C1(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__inv_2 _1051_ (.A(\send_divcnt[19] ),
    .Y(_0451_));
 sky130_fd_sc_hd__inv_2 _1052_ (.A(\send_divcnt[18] ),
    .Y(_0452_));
 sky130_fd_sc_hd__inv_2 _1053_ (.A(net91),
    .Y(_0453_));
 sky130_fd_sc_hd__inv_2 _1054_ (.A(net90),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_2 _1055_ (.A(net92),
    .Y(_0455_));
 sky130_fd_sc_hd__o22a_1 _1056_ (.A1(_0320_),
    .A2(\send_divcnt[20] ),
    .B1(\send_divcnt[19] ),
    .B2(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__o221a_1 _1057_ (.A1(_0453_),
    .A2(\send_divcnt[18] ),
    .B1(\send_divcnt[17] ),
    .B2(_0454_),
    .C1(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__o221a_1 _1058_ (.A1(net92),
    .A2(_0451_),
    .B1(_0452_),
    .B2(net91),
    .C1(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__and4_1 _1059_ (.A(_0446_),
    .B(_0447_),
    .C(_0450_),
    .D(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__or3_1 _1060_ (.A(_0300_),
    .B(\send_divcnt[16] ),
    .C(_0444_),
    .X(_0460_));
 sky130_fd_sc_hd__a22o_1 _1061_ (.A1(_0455_),
    .A2(\send_divcnt[19] ),
    .B1(\send_divcnt[18] ),
    .B2(_0453_),
    .X(_0461_));
 sky130_fd_sc_hd__a221o_1 _1062_ (.A1(_0460_),
    .A2(_0457_),
    .B1(_0461_),
    .B2(_0456_),
    .C1(_0445_),
    .X(_0462_));
 sky130_fd_sc_hd__o21ai_1 _1063_ (.A1(_0319_),
    .A2(\send_divcnt[21] ),
    .B1(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__a21bo_1 _1064_ (.A1(_0449_),
    .A2(_0463_),
    .B1_N(_0402_),
    .X(_0464_));
 sky130_fd_sc_hd__a32o_2 _1065_ (.A1(_0402_),
    .A2(_0442_),
    .A3(_0459_),
    .B1(_0464_),
    .B2(_0448_),
    .X(_0465_));
 sky130_fd_sc_hd__inv_2 _1066_ (.A(\send_divcnt[25] ),
    .Y(_0466_));
 sky130_fd_sc_hd__o22a_1 _1067_ (.A1(_0290_),
    .A2(\send_divcnt[25] ),
    .B1(\send_divcnt[24] ),
    .B2(_0294_),
    .X(_0467_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(\send_divcnt[26] ),
    .Y(_0468_));
 sky130_fd_sc_hd__inv_2 _1069_ (.A(\send_divcnt[29] ),
    .Y(_0469_));
 sky130_fd_sc_hd__o2bb2a_1 _1070_ (.A1_N(\send_divcnt[28] ),
    .A2_N(_0283_),
    .B1(net103),
    .B2(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__o221a_1 _1071_ (.A1(_0288_),
    .A2(\send_divcnt[27] ),
    .B1(_0468_),
    .B2(net100),
    .C1(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__o221a_1 _1072_ (.A1(_0222_),
    .A2(\send_divcnt[31] ),
    .B1(\send_divcnt[30] ),
    .B2(_0335_),
    .C1(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__inv_2 _1073_ (.A(net103),
    .Y(_0473_));
 sky130_fd_sc_hd__nor2_1 _1074_ (.A(_0473_),
    .B(\send_divcnt[29] ),
    .Y(_0474_));
 sky130_fd_sc_hd__and2_1 _1075_ (.A(_0288_),
    .B(\send_divcnt[27] ),
    .X(_0475_));
 sky130_fd_sc_hd__nor2_1 _1076_ (.A(_0283_),
    .B(\send_divcnt[28] ),
    .Y(_0476_));
 sky130_fd_sc_hd__inv_2 _1077_ (.A(\send_divcnt[30] ),
    .Y(_0477_));
 sky130_fd_sc_hd__nand2_1 _1078_ (.A(_0222_),
    .B(\send_divcnt[31] ),
    .Y(_0478_));
 sky130_fd_sc_hd__o21ai_1 _1079_ (.A1(net105),
    .A2(_0477_),
    .B1(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__a2111o_1 _1080_ (.A1(_0294_),
    .A2(\send_divcnt[24] ),
    .B1(_0475_),
    .C1(_0476_),
    .D1(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__a211oi_1 _1081_ (.A1(net100),
    .A2(_0468_),
    .B1(_0474_),
    .C1(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__o2111a_1 _1082_ (.A1(net99),
    .A2(_0466_),
    .B1(_0467_),
    .C1(_0472_),
    .D1(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__inv_2 _1083_ (.A(\send_divcnt[31] ),
    .Y(_0483_));
 sky130_fd_sc_hd__nor2_1 _1084_ (.A(_0288_),
    .B(\send_divcnt[27] ),
    .Y(_0484_));
 sky130_fd_sc_hd__a221o_1 _1085_ (.A1(_0286_),
    .A2(\send_divcnt[26] ),
    .B1(\send_divcnt[25] ),
    .B2(_0290_),
    .C1(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__o22a_1 _1086_ (.A1(_0286_),
    .A2(\send_divcnt[26] ),
    .B1(_0467_),
    .B2(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__nor2_1 _1087_ (.A(_0475_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__o31a_1 _1088_ (.A1(_0484_),
    .A2(_0476_),
    .A3(_0487_),
    .B1(_0470_),
    .X(_0488_));
 sky130_fd_sc_hd__o22a_1 _1089_ (.A1(net105),
    .A2(_0477_),
    .B1(_0474_),
    .B2(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__a221o_1 _1090_ (.A1(net106),
    .A2(_0483_),
    .B1(_0477_),
    .B2(net105),
    .C1(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__nor2_2 _1091_ (.A(\send_bitcnt[3] ),
    .B(_0204_),
    .Y(_0491_));
 sky130_fd_sc_hd__a221oi_4 _1092_ (.A1(_0465_),
    .A2(_0482_),
    .B1(_0490_),
    .B2(_0478_),
    .C1(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__clkbuf_4 _1093_ (.A(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__and2_1 _1094_ (.A(net10),
    .B(_0491_),
    .X(_0494_));
 sky130_fd_sc_hd__clkbuf_4 _1095_ (.A(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__nor2_4 _1096_ (.A(_0492_),
    .B(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__inv_2 _1097_ (.A(net47),
    .Y(_0497_));
 sky130_fd_sc_hd__and2_1 _1098_ (.A(send_dummy),
    .B(_0491_),
    .X(_0498_));
 sky130_fd_sc_hd__or2_1 _1099_ (.A(_0497_),
    .B(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_4 _1100_ (.A(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__a221o_1 _1101_ (.A1(\send_pattern[1] ),
    .A2(_0493_),
    .B1(_0496_),
    .B2(net114),
    .C1(_0500_),
    .X(_0025_));
 sky130_fd_sc_hd__a221o_1 _1102_ (.A1(\send_pattern[2] ),
    .A2(_0493_),
    .B1(_0495_),
    .B2(net1),
    .C1(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__a21o_1 _1103_ (.A1(\send_pattern[1] ),
    .A2(_0496_),
    .B1(_0501_),
    .X(_0026_));
 sky130_fd_sc_hd__a221o_1 _1104_ (.A1(\send_pattern[3] ),
    .A2(_0493_),
    .B1(_0495_),
    .B2(net2),
    .C1(_0500_),
    .X(_0502_));
 sky130_fd_sc_hd__a21o_1 _1105_ (.A1(\send_pattern[2] ),
    .A2(_0496_),
    .B1(_0502_),
    .X(_0027_));
 sky130_fd_sc_hd__a221o_1 _1106_ (.A1(\send_pattern[4] ),
    .A2(_0493_),
    .B1(_0495_),
    .B2(net3),
    .C1(_0500_),
    .X(_0503_));
 sky130_fd_sc_hd__a21o_1 _1107_ (.A1(\send_pattern[3] ),
    .A2(_0496_),
    .B1(_0503_),
    .X(_0028_));
 sky130_fd_sc_hd__a221o_1 _1108_ (.A1(\send_pattern[5] ),
    .A2(_0493_),
    .B1(_0495_),
    .B2(net4),
    .C1(_0500_),
    .X(_0504_));
 sky130_fd_sc_hd__a21o_1 _1109_ (.A1(\send_pattern[4] ),
    .A2(_0496_),
    .B1(_0504_),
    .X(_0029_));
 sky130_fd_sc_hd__a221o_1 _1110_ (.A1(\send_pattern[6] ),
    .A2(_0493_),
    .B1(_0495_),
    .B2(net5),
    .C1(_0500_),
    .X(_0505_));
 sky130_fd_sc_hd__a21o_1 _1111_ (.A1(\send_pattern[5] ),
    .A2(_0496_),
    .B1(_0505_),
    .X(_0030_));
 sky130_fd_sc_hd__a221o_1 _1112_ (.A1(\send_pattern[7] ),
    .A2(_0493_),
    .B1(_0495_),
    .B2(net6),
    .C1(_0500_),
    .X(_0506_));
 sky130_fd_sc_hd__a21o_1 _1113_ (.A1(\send_pattern[6] ),
    .A2(_0496_),
    .B1(_0506_),
    .X(_0031_));
 sky130_fd_sc_hd__a221o_1 _1114_ (.A1(\send_pattern[8] ),
    .A2(_0493_),
    .B1(_0495_),
    .B2(net7),
    .C1(_0500_),
    .X(_0507_));
 sky130_fd_sc_hd__a21o_1 _1115_ (.A1(\send_pattern[7] ),
    .A2(_0496_),
    .B1(_0507_),
    .X(_0032_));
 sky130_fd_sc_hd__or3_2 _1116_ (.A(_0492_),
    .B(_0494_),
    .C(_0498_),
    .X(_0508_));
 sky130_fd_sc_hd__or2_4 _1117_ (.A(_0497_),
    .B(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__or3b_1 _1118_ (.A(_0500_),
    .B(net8),
    .C_N(_0495_),
    .X(_0510_));
 sky130_fd_sc_hd__o21a_1 _1119_ (.A1(\send_pattern[8] ),
    .A2(_0509_),
    .B1(_0510_),
    .X(_0033_));
 sky130_fd_sc_hd__inv_2 _1120_ (.A(\send_bitcnt[0] ),
    .Y(_0511_));
 sky130_fd_sc_hd__and2_1 _1121_ (.A(_0511_),
    .B(_0508_),
    .X(_0512_));
 sky130_fd_sc_hd__nor2_1 _1122_ (.A(_0497_),
    .B(_0508_),
    .Y(_0513_));
 sky130_fd_sc_hd__buf_4 _1123_ (.A(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__a32o_1 _1124_ (.A1(_0351_),
    .A2(_0205_),
    .A3(_0512_),
    .B1(_0514_),
    .B2(\send_bitcnt[0] ),
    .X(_0034_));
 sky130_fd_sc_hd__a21o_1 _1125_ (.A1(_0511_),
    .A2(_0508_),
    .B1(\send_bitcnt[1] ),
    .X(_0515_));
 sky130_fd_sc_hd__nand3_1 _1126_ (.A(\send_bitcnt[1] ),
    .B(_0511_),
    .C(_0508_),
    .Y(_0516_));
 sky130_fd_sc_hd__and3_1 _1127_ (.A(_0349_),
    .B(_0515_),
    .C(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_1 _1128_ (.A(_0517_),
    .X(_0035_));
 sky130_fd_sc_hd__o21ai_1 _1129_ (.A1(\send_bitcnt[1] ),
    .A2(\send_bitcnt[0] ),
    .B1(\send_bitcnt[2] ),
    .Y(_0518_));
 sky130_fd_sc_hd__nand2_1 _1130_ (.A(_0204_),
    .B(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__mux2_1 _1131_ (.A0(\send_bitcnt[2] ),
    .A1(_0519_),
    .S(_0493_),
    .X(_0520_));
 sky130_fd_sc_hd__o21a_1 _1132_ (.A1(_0498_),
    .A2(_0520_),
    .B1(_0350_),
    .X(_0036_));
 sky130_fd_sc_hd__and2_1 _1133_ (.A(_0491_),
    .B(_0508_),
    .X(_0521_));
 sky130_fd_sc_hd__o21a_1 _1134_ (.A1(_0204_),
    .A2(_0496_),
    .B1(\send_bitcnt[3] ),
    .X(_0522_));
 sky130_fd_sc_hd__o21a_1 _1135_ (.A1(_0521_),
    .A2(_0522_),
    .B1(_0350_),
    .X(_0037_));
 sky130_fd_sc_hd__or4_1 _1136_ (.A(net43),
    .B(send_dummy),
    .C(net46),
    .D(net44),
    .X(_0523_));
 sky130_fd_sc_hd__nor2_2 _1137_ (.A(net45),
    .B(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__o21ai_1 _1138_ (.A1(_0498_),
    .A2(_0524_),
    .B1(_0350_),
    .Y(_0038_));
 sky130_fd_sc_hd__or3_2 _1139_ (.A(\recv_state[3] ),
    .B(\recv_state[2] ),
    .C(\recv_state[1] ),
    .X(_0525_));
 sky130_fd_sc_hd__nor2_1 _1140_ (.A(\recv_state[0] ),
    .B(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__a22oi_2 _1141_ (.A1(_0347_),
    .A2(_0525_),
    .B1(_0526_),
    .B2(net48),
    .Y(_0527_));
 sky130_fd_sc_hd__o22a_1 _1142_ (.A1(_0283_),
    .A2(\recv_divcnt[27] ),
    .B1(\recv_divcnt[26] ),
    .B2(_0288_),
    .X(_0528_));
 sky130_fd_sc_hd__and2_1 _1143_ (.A(_0283_),
    .B(\recv_divcnt[27] ),
    .X(_0529_));
 sky130_fd_sc_hd__a21oi_1 _1144_ (.A1(_0288_),
    .A2(\recv_divcnt[26] ),
    .B1(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__o211a_1 _1145_ (.A1(net100),
    .A2(_0296_),
    .B1(_0528_),
    .C1(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__nand2_1 _1146_ (.A(_0313_),
    .B(\recv_divcnt[22] ),
    .Y(_0532_));
 sky130_fd_sc_hd__nand2_1 _1147_ (.A(net97),
    .B(_0312_),
    .Y(_0533_));
 sky130_fd_sc_hd__xnor2_1 _1148_ (.A(net98),
    .B(\recv_divcnt[23] ),
    .Y(_0534_));
 sky130_fd_sc_hd__and3_1 _1149_ (.A(_0532_),
    .B(_0533_),
    .C(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__nand2_1 _1150_ (.A(_0315_),
    .B(\recv_divcnt[21] ),
    .Y(_0536_));
 sky130_fd_sc_hd__nor2_1 _1151_ (.A(_0315_),
    .B(\recv_divcnt[21] ),
    .Y(_0537_));
 sky130_fd_sc_hd__a31o_1 _1152_ (.A1(net95),
    .A2(_0304_),
    .A3(_0536_),
    .B1(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__a21oi_1 _1153_ (.A1(_0294_),
    .A2(\recv_divcnt[23] ),
    .B1(_0533_),
    .Y(_0539_));
 sky130_fd_sc_hd__a221o_1 _1154_ (.A1(net98),
    .A2(_0328_),
    .B1(_0535_),
    .B2(_0538_),
    .C1(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__nor2_1 _1155_ (.A(_0320_),
    .B(\recv_divcnt[19] ),
    .Y(_0541_));
 sky130_fd_sc_hd__o211a_1 _1156_ (.A1(net94),
    .A2(_0305_),
    .B1(_0329_),
    .C1(net92),
    .X(_0542_));
 sky130_fd_sc_hd__a22o_1 _1157_ (.A1(net91),
    .A2(_0301_),
    .B1(_0302_),
    .B2(net90),
    .X(_0543_));
 sky130_fd_sc_hd__xnor2_1 _1158_ (.A(net92),
    .B(\recv_divcnt[18] ),
    .Y(_0544_));
 sky130_fd_sc_hd__nor2_1 _1159_ (.A(net94),
    .B(_0305_),
    .Y(_0545_));
 sky130_fd_sc_hd__nor2_1 _1160_ (.A(_0541_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__o2111a_1 _1161_ (.A1(net91),
    .A2(_0301_),
    .B1(_0543_),
    .C1(_0544_),
    .D1(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__a21oi_1 _1162_ (.A1(_0319_),
    .A2(\recv_divcnt[20] ),
    .B1(_0537_),
    .Y(_0548_));
 sky130_fd_sc_hd__o2111a_1 _1163_ (.A1(_0319_),
    .A2(\recv_divcnt[20] ),
    .B1(_0536_),
    .C1(_0535_),
    .D1(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__o31a_1 _1164_ (.A1(_0541_),
    .A2(_0542_),
    .A3(_0547_),
    .B1(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__or2b_1 _1165_ (.A(\recv_divcnt[1] ),
    .B_N(net104),
    .X(_0551_));
 sky130_fd_sc_hd__and2b_1 _1166_ (.A_N(net107),
    .B(\recv_divcnt[2] ),
    .X(_0552_));
 sky130_fd_sc_hd__and2b_1 _1167_ (.A_N(net104),
    .B(\recv_divcnt[1] ),
    .X(_0553_));
 sky130_fd_sc_hd__a311o_1 _1168_ (.A1(_0238_),
    .A2(\recv_divcnt[0] ),
    .A3(_0551_),
    .B1(_0552_),
    .C1(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__o22a_1 _1169_ (.A1(_0232_),
    .A2(\recv_divcnt[3] ),
    .B1(\recv_divcnt[2] ),
    .B2(_0235_),
    .X(_0555_));
 sky130_fd_sc_hd__a22o_1 _1170_ (.A1(_0231_),
    .A2(\recv_divcnt[4] ),
    .B1(\recv_divcnt[3] ),
    .B2(_0232_),
    .X(_0556_));
 sky130_fd_sc_hd__a21o_1 _1171_ (.A1(_0554_),
    .A2(_0555_),
    .B1(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__o22a_1 _1172_ (.A1(_0246_),
    .A2(\recv_divcnt[5] ),
    .B1(\recv_divcnt[4] ),
    .B2(_0231_),
    .X(_0558_));
 sky130_fd_sc_hd__a22o_1 _1173_ (.A1(_0229_),
    .A2(\recv_divcnt[6] ),
    .B1(\recv_divcnt[5] ),
    .B2(_0246_),
    .X(_0559_));
 sky130_fd_sc_hd__and2b_1 _1174_ (.A_N(net112),
    .B(\recv_divcnt[7] ),
    .X(_0560_));
 sky130_fd_sc_hd__a211o_1 _1175_ (.A1(net111),
    .A2(_0247_),
    .B1(_0559_),
    .C1(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__a21o_1 _1176_ (.A1(_0557_),
    .A2(_0558_),
    .B1(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__or3_1 _1177_ (.A(_0229_),
    .B(\recv_divcnt[6] ),
    .C(_0560_),
    .X(_0563_));
 sky130_fd_sc_hd__or2b_1 _1178_ (.A(\recv_divcnt[7] ),
    .B_N(net112),
    .X(_0564_));
 sky130_fd_sc_hd__o22a_1 _1179_ (.A1(_0258_),
    .A2(\recv_divcnt[11] ),
    .B1(\recv_divcnt[10] ),
    .B2(_0270_),
    .X(_0565_));
 sky130_fd_sc_hd__and2b_1 _1180_ (.A_N(net85),
    .B(\recv_divcnt[11] ),
    .X(_0566_));
 sky130_fd_sc_hd__a221oi_1 _1181_ (.A1(_0270_),
    .A2(\recv_divcnt[10] ),
    .B1(\recv_divcnt[9] ),
    .B2(_0268_),
    .C1(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_1 _1182_ (.A(_0565_),
    .B(_0567_),
    .Y(_0568_));
 sky130_fd_sc_hd__and2b_1 _1183_ (.A_N(net88),
    .B(\recv_divcnt[14] ),
    .X(_0569_));
 sky130_fd_sc_hd__and2b_1 _1184_ (.A_N(net87),
    .B(\recv_divcnt[13] ),
    .X(_0570_));
 sky130_fd_sc_hd__and2b_1 _1185_ (.A_N(net89),
    .B(\recv_divcnt[15] ),
    .X(_0571_));
 sky130_fd_sc_hd__a2111o_1 _1186_ (.A1(_0257_),
    .A2(\recv_divcnt[12] ),
    .B1(_0569_),
    .C1(_0570_),
    .D1(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__a2bb2o_1 _1187_ (.A1_N(_0300_),
    .A2_N(\recv_divcnt[15] ),
    .B1(_0254_),
    .B2(net88),
    .X(_0573_));
 sky130_fd_sc_hd__a2bb2o_1 _1188_ (.A1_N(\recv_divcnt[12] ),
    .A2_N(_0257_),
    .B1(net87),
    .B2(_0264_),
    .X(_0574_));
 sky130_fd_sc_hd__or3_1 _1189_ (.A(_0572_),
    .B(_0573_),
    .C(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__nor2_1 _1190_ (.A(net113),
    .B(_0261_),
    .Y(_0576_));
 sky130_fd_sc_hd__o22a_1 _1191_ (.A1(_0268_),
    .A2(\recv_divcnt[9] ),
    .B1(\recv_divcnt[8] ),
    .B2(_0415_),
    .X(_0577_));
 sky130_fd_sc_hd__or4b_1 _1192_ (.A(_0568_),
    .B(_0575_),
    .C(_0576_),
    .D_N(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__a31o_1 _1193_ (.A1(_0562_),
    .A2(_0563_),
    .A3(_0564_),
    .B1(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__o22a_1 _1194_ (.A1(_0565_),
    .A2(_0566_),
    .B1(_0568_),
    .B2(_0577_),
    .X(_0580_));
 sky130_fd_sc_hd__nor2_1 _1195_ (.A(_0569_),
    .B(_0570_),
    .Y(_0581_));
 sky130_fd_sc_hd__a21oi_1 _1196_ (.A1(_0581_),
    .A2(_0574_),
    .B1(_0573_),
    .Y(_0582_));
 sky130_fd_sc_hd__o22a_1 _1197_ (.A1(_0575_),
    .A2(_0580_),
    .B1(_0582_),
    .B2(_0571_),
    .X(_0583_));
 sky130_fd_sc_hd__o221a_1 _1198_ (.A1(net91),
    .A2(_0301_),
    .B1(_0302_),
    .B2(net90),
    .C1(_0544_),
    .X(_0584_));
 sky130_fd_sc_hd__nand4b_1 _1199_ (.A_N(_0543_),
    .B(_0549_),
    .C(_0546_),
    .D(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__a21o_1 _1200_ (.A1(_0579_),
    .A2(_0583_),
    .B1(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__or3b_1 _1201_ (.A(_0540_),
    .B(_0550_),
    .C_N(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__a22o_1 _1202_ (.A1(net100),
    .A2(_0296_),
    .B1(_0297_),
    .B2(net99),
    .X(_0588_));
 sky130_fd_sc_hd__a21oi_1 _1203_ (.A1(_0290_),
    .A2(\recv_divcnt[24] ),
    .B1(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__a2bb2o_1 _1204_ (.A1_N(_0529_),
    .A2_N(_0528_),
    .B1(_0531_),
    .B2(_0588_),
    .X(_0590_));
 sky130_fd_sc_hd__a31o_1 _1205_ (.A1(_0531_),
    .A2(_0587_),
    .A3(_0589_),
    .B1(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__o22a_1 _1206_ (.A1(_0335_),
    .A2(\recv_divcnt[29] ),
    .B1(\recv_divcnt[28] ),
    .B2(_0473_),
    .X(_0592_));
 sky130_fd_sc_hd__nand2_1 _1207_ (.A(_0335_),
    .B(\recv_divcnt[29] ),
    .Y(_0593_));
 sky130_fd_sc_hd__o211a_1 _1208_ (.A1(net103),
    .A2(_0226_),
    .B1(_0592_),
    .C1(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__and2b_1 _1209_ (.A_N(_0592_),
    .B(_0593_),
    .X(_0595_));
 sky130_fd_sc_hd__a221o_1 _1210_ (.A1(net106),
    .A2(_0336_),
    .B1(_0591_),
    .B2(_0594_),
    .C1(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__inv_2 _1211_ (.A(_0525_),
    .Y(_0597_));
 sky130_fd_sc_hd__o211a_1 _1212_ (.A1(net106),
    .A2(_0336_),
    .B1(_0597_),
    .C1(\recv_state[0] ),
    .X(_0598_));
 sky130_fd_sc_hd__a21boi_1 _1213_ (.A1(_0596_),
    .A2(_0598_),
    .B1_N(_0527_),
    .Y(_0599_));
 sky130_fd_sc_hd__nand2_1 _1214_ (.A(\recv_state[0] ),
    .B(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__o2111a_1 _1215_ (.A1(\recv_state[0] ),
    .A2(_0527_),
    .B1(_0600_),
    .C1(_0351_),
    .D1(_0219_),
    .X(_0039_));
 sky130_fd_sc_hd__inv_2 _1216_ (.A(\recv_state[2] ),
    .Y(_0601_));
 sky130_fd_sc_hd__a31o_1 _1217_ (.A1(\recv_state[3] ),
    .A2(_0601_),
    .A3(_0599_),
    .B1(_0217_),
    .X(_0602_));
 sky130_fd_sc_hd__and3_1 _1218_ (.A(\recv_state[1] ),
    .B(\recv_state[0] ),
    .C(_0527_),
    .X(_0603_));
 sky130_fd_sc_hd__a211oi_1 _1219_ (.A1(_0600_),
    .A2(_0602_),
    .B1(_0603_),
    .C1(_0497_),
    .Y(_0040_));
 sky130_fd_sc_hd__and4_1 _1220_ (.A(\recv_state[2] ),
    .B(\recv_state[1] ),
    .C(\recv_state[0] ),
    .D(_0527_),
    .X(_0604_));
 sky130_fd_sc_hd__o21ai_1 _1221_ (.A1(\recv_state[2] ),
    .A2(_0603_),
    .B1(_0351_),
    .Y(_0605_));
 sky130_fd_sc_hd__nor2_1 _1222_ (.A(_0604_),
    .B(_0605_),
    .Y(_0041_));
 sky130_fd_sc_hd__nand2_1 _1223_ (.A(_0218_),
    .B(_0525_),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2_1 _1224_ (.A(_0599_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__xnor2_1 _1225_ (.A(_0216_),
    .B(_0604_),
    .Y(_0608_));
 sky130_fd_sc_hd__and3_1 _1226_ (.A(_0349_),
    .B(_0607_),
    .C(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__clkbuf_1 _1227_ (.A(_0609_),
    .X(_0042_));
 sky130_fd_sc_hd__nor2_1 _1228_ (.A(\send_divcnt[0] ),
    .B(_0509_),
    .Y(_0043_));
 sky130_fd_sc_hd__or2_1 _1229_ (.A(\send_divcnt[1] ),
    .B(\send_divcnt[0] ),
    .X(_0610_));
 sky130_fd_sc_hd__nand2_1 _1230_ (.A(\send_divcnt[1] ),
    .B(\send_divcnt[0] ),
    .Y(_0611_));
 sky130_fd_sc_hd__and3_1 _1231_ (.A(_0514_),
    .B(_0610_),
    .C(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__clkbuf_1 _1232_ (.A(_0612_),
    .X(_0044_));
 sky130_fd_sc_hd__inv_2 _1233_ (.A(\send_divcnt[2] ),
    .Y(_0613_));
 sky130_fd_sc_hd__nor2_1 _1234_ (.A(_0613_),
    .B(_0611_),
    .Y(_0614_));
 sky130_fd_sc_hd__nand2_1 _1235_ (.A(_0613_),
    .B(_0611_),
    .Y(_0615_));
 sky130_fd_sc_hd__clkbuf_4 _1236_ (.A(_0513_),
    .X(_0616_));
 sky130_fd_sc_hd__buf_4 _1237_ (.A(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__and3b_1 _1238_ (.A_N(_0614_),
    .B(_0615_),
    .C(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__clkbuf_1 _1239_ (.A(_0618_),
    .X(_0045_));
 sky130_fd_sc_hd__and4_1 _1240_ (.A(\send_divcnt[3] ),
    .B(\send_divcnt[2] ),
    .C(\send_divcnt[1] ),
    .D(\send_divcnt[0] ),
    .X(_0619_));
 sky130_fd_sc_hd__or2_1 _1241_ (.A(\send_divcnt[3] ),
    .B(_0614_),
    .X(_0620_));
 sky130_fd_sc_hd__and3b_1 _1242_ (.A_N(_0619_),
    .B(_0620_),
    .C(_0617_),
    .X(_0621_));
 sky130_fd_sc_hd__clkbuf_1 _1243_ (.A(_0621_),
    .X(_0046_));
 sky130_fd_sc_hd__nand2_1 _1244_ (.A(\send_divcnt[4] ),
    .B(_0619_),
    .Y(_0622_));
 sky130_fd_sc_hd__or2_1 _1245_ (.A(\send_divcnt[4] ),
    .B(_0619_),
    .X(_0623_));
 sky130_fd_sc_hd__and3_1 _1246_ (.A(_0514_),
    .B(_0622_),
    .C(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__clkbuf_1 _1247_ (.A(_0624_),
    .X(_0047_));
 sky130_fd_sc_hd__nor2_1 _1248_ (.A(_0421_),
    .B(_0622_),
    .Y(_0625_));
 sky130_fd_sc_hd__nand2_1 _1249_ (.A(_0421_),
    .B(_0622_),
    .Y(_0626_));
 sky130_fd_sc_hd__and3b_1 _1250_ (.A_N(_0625_),
    .B(_0626_),
    .C(_0617_),
    .X(_0627_));
 sky130_fd_sc_hd__clkbuf_1 _1251_ (.A(_0627_),
    .X(_0048_));
 sky130_fd_sc_hd__and4_1 _1252_ (.A(\send_divcnt[6] ),
    .B(\send_divcnt[5] ),
    .C(\send_divcnt[4] ),
    .D(_0619_),
    .X(_0628_));
 sky130_fd_sc_hd__or2_1 _1253_ (.A(\send_divcnt[6] ),
    .B(_0625_),
    .X(_0629_));
 sky130_fd_sc_hd__and3b_1 _1254_ (.A_N(_0628_),
    .B(_0629_),
    .C(_0617_),
    .X(_0630_));
 sky130_fd_sc_hd__clkbuf_1 _1255_ (.A(_0630_),
    .X(_0049_));
 sky130_fd_sc_hd__nand2_1 _1256_ (.A(\send_divcnt[7] ),
    .B(_0628_),
    .Y(_0631_));
 sky130_fd_sc_hd__or2_1 _1257_ (.A(\send_divcnt[7] ),
    .B(_0628_),
    .X(_0632_));
 sky130_fd_sc_hd__and3_1 _1258_ (.A(_0514_),
    .B(_0631_),
    .C(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_1 _1259_ (.A(_0633_),
    .X(_0050_));
 sky130_fd_sc_hd__nor2_1 _1260_ (.A(_0411_),
    .B(_0631_),
    .Y(_0634_));
 sky130_fd_sc_hd__nand2_1 _1261_ (.A(_0411_),
    .B(_0631_),
    .Y(_0635_));
 sky130_fd_sc_hd__and3b_1 _1262_ (.A_N(_0634_),
    .B(_0635_),
    .C(_0617_),
    .X(_0636_));
 sky130_fd_sc_hd__clkbuf_1 _1263_ (.A(_0636_),
    .X(_0051_));
 sky130_fd_sc_hd__nand2_1 _1264_ (.A(\send_divcnt[9] ),
    .B(_0634_),
    .Y(_0637_));
 sky130_fd_sc_hd__or2_1 _1265_ (.A(\send_divcnt[9] ),
    .B(_0634_),
    .X(_0638_));
 sky130_fd_sc_hd__and3_1 _1266_ (.A(_0514_),
    .B(_0637_),
    .C(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__clkbuf_1 _1267_ (.A(_0639_),
    .X(_0052_));
 sky130_fd_sc_hd__nor2_1 _1268_ (.A(_0408_),
    .B(_0413_),
    .Y(_0640_));
 sky130_fd_sc_hd__and4_1 _1269_ (.A(\send_divcnt[8] ),
    .B(\send_divcnt[7] ),
    .C(_0628_),
    .D(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__a211oi_1 _1270_ (.A1(_0408_),
    .A2(_0637_),
    .B1(_0641_),
    .C1(_0509_),
    .Y(_0053_));
 sky130_fd_sc_hd__and2_1 _1271_ (.A(\send_divcnt[11] ),
    .B(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__or2_1 _1272_ (.A(\send_divcnt[11] ),
    .B(_0641_),
    .X(_0643_));
 sky130_fd_sc_hd__and3b_1 _1273_ (.A_N(_0642_),
    .B(_0643_),
    .C(_0617_),
    .X(_0644_));
 sky130_fd_sc_hd__clkbuf_1 _1274_ (.A(_0644_),
    .X(_0054_));
 sky130_fd_sc_hd__and3_1 _1275_ (.A(\send_divcnt[12] ),
    .B(\send_divcnt[11] ),
    .C(_0641_),
    .X(_0645_));
 sky130_fd_sc_hd__or2_1 _1276_ (.A(\send_divcnt[12] ),
    .B(_0642_),
    .X(_0646_));
 sky130_fd_sc_hd__and3b_1 _1277_ (.A_N(_0645_),
    .B(_0646_),
    .C(_0617_),
    .X(_0647_));
 sky130_fd_sc_hd__clkbuf_1 _1278_ (.A(_0647_),
    .X(_0055_));
 sky130_fd_sc_hd__and4_1 _1279_ (.A(\send_divcnt[13] ),
    .B(\send_divcnt[12] ),
    .C(\send_divcnt[11] ),
    .D(_0641_),
    .X(_0648_));
 sky130_fd_sc_hd__or2_1 _1280_ (.A(\send_divcnt[13] ),
    .B(_0645_),
    .X(_0649_));
 sky130_fd_sc_hd__and3b_1 _1281_ (.A_N(_0648_),
    .B(_0649_),
    .C(_0616_),
    .X(_0650_));
 sky130_fd_sc_hd__clkbuf_1 _1282_ (.A(_0650_),
    .X(_0056_));
 sky130_fd_sc_hd__nand2_1 _1283_ (.A(\send_divcnt[14] ),
    .B(_0648_),
    .Y(_0651_));
 sky130_fd_sc_hd__or2_1 _1284_ (.A(\send_divcnt[14] ),
    .B(_0648_),
    .X(_0652_));
 sky130_fd_sc_hd__and3_1 _1285_ (.A(_0514_),
    .B(_0651_),
    .C(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__clkbuf_1 _1286_ (.A(_0653_),
    .X(_0057_));
 sky130_fd_sc_hd__and3_1 _1287_ (.A(\send_divcnt[15] ),
    .B(\send_divcnt[14] ),
    .C(_0648_),
    .X(_0654_));
 sky130_fd_sc_hd__a21o_1 _1288_ (.A1(\send_divcnt[14] ),
    .A2(_0648_),
    .B1(\send_divcnt[15] ),
    .X(_0655_));
 sky130_fd_sc_hd__and3b_1 _1289_ (.A_N(_0654_),
    .B(_0655_),
    .C(_0616_),
    .X(_0656_));
 sky130_fd_sc_hd__clkbuf_1 _1290_ (.A(_0656_),
    .X(_0058_));
 sky130_fd_sc_hd__nand2_1 _1291_ (.A(\send_divcnt[16] ),
    .B(_0654_),
    .Y(_0657_));
 sky130_fd_sc_hd__or2_1 _1292_ (.A(\send_divcnt[16] ),
    .B(_0654_),
    .X(_0658_));
 sky130_fd_sc_hd__and3_1 _1293_ (.A(_0514_),
    .B(_0657_),
    .C(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__clkbuf_1 _1294_ (.A(_0659_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _1295_ (.A(\send_divcnt[17] ),
    .B(\send_divcnt[16] ),
    .X(_0660_));
 sky130_fd_sc_hd__and4_1 _1296_ (.A(\send_divcnt[15] ),
    .B(\send_divcnt[14] ),
    .C(_0648_),
    .D(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__a211oi_1 _1297_ (.A1(_0443_),
    .A2(_0657_),
    .B1(_0661_),
    .C1(_0509_),
    .Y(_0060_));
 sky130_fd_sc_hd__and2_1 _1298_ (.A(\send_divcnt[18] ),
    .B(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__or2_1 _1299_ (.A(\send_divcnt[18] ),
    .B(_0661_),
    .X(_0663_));
 sky130_fd_sc_hd__and3b_1 _1300_ (.A_N(_0662_),
    .B(_0663_),
    .C(_0616_),
    .X(_0664_));
 sky130_fd_sc_hd__clkbuf_1 _1301_ (.A(_0664_),
    .X(_0061_));
 sky130_fd_sc_hd__and3_1 _1302_ (.A(\send_divcnt[19] ),
    .B(\send_divcnt[18] ),
    .C(_0661_),
    .X(_0665_));
 sky130_fd_sc_hd__or2_1 _1303_ (.A(\send_divcnt[19] ),
    .B(_0662_),
    .X(_0666_));
 sky130_fd_sc_hd__and3b_1 _1304_ (.A_N(_0665_),
    .B(_0666_),
    .C(_0616_),
    .X(_0667_));
 sky130_fd_sc_hd__clkbuf_1 _1305_ (.A(_0667_),
    .X(_0062_));
 sky130_fd_sc_hd__and4_1 _1306_ (.A(\send_divcnt[20] ),
    .B(\send_divcnt[19] ),
    .C(\send_divcnt[18] ),
    .D(_0661_),
    .X(_0668_));
 sky130_fd_sc_hd__or2_1 _1307_ (.A(\send_divcnt[20] ),
    .B(_0665_),
    .X(_0669_));
 sky130_fd_sc_hd__and3b_1 _1308_ (.A_N(_0668_),
    .B(_0669_),
    .C(_0616_),
    .X(_0670_));
 sky130_fd_sc_hd__clkbuf_1 _1309_ (.A(_0670_),
    .X(_0063_));
 sky130_fd_sc_hd__nand2_1 _1310_ (.A(\send_divcnt[21] ),
    .B(_0668_),
    .Y(_0671_));
 sky130_fd_sc_hd__or2_1 _1311_ (.A(\send_divcnt[21] ),
    .B(_0668_),
    .X(_0672_));
 sky130_fd_sc_hd__and3_1 _1312_ (.A(_0514_),
    .B(_0671_),
    .C(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__clkbuf_1 _1313_ (.A(_0673_),
    .X(_0064_));
 sky130_fd_sc_hd__and3_1 _1314_ (.A(\send_divcnt[22] ),
    .B(\send_divcnt[21] ),
    .C(_0668_),
    .X(_0674_));
 sky130_fd_sc_hd__a21o_1 _1315_ (.A1(\send_divcnt[21] ),
    .A2(_0668_),
    .B1(\send_divcnt[22] ),
    .X(_0675_));
 sky130_fd_sc_hd__and3b_1 _1316_ (.A_N(_0674_),
    .B(_0675_),
    .C(_0616_),
    .X(_0676_));
 sky130_fd_sc_hd__clkbuf_1 _1317_ (.A(_0676_),
    .X(_0065_));
 sky130_fd_sc_hd__and4_1 _1318_ (.A(\send_divcnt[23] ),
    .B(\send_divcnt[22] ),
    .C(\send_divcnt[21] ),
    .D(_0668_),
    .X(_0677_));
 sky130_fd_sc_hd__or2_1 _1319_ (.A(\send_divcnt[23] ),
    .B(_0674_),
    .X(_0678_));
 sky130_fd_sc_hd__and3b_1 _1320_ (.A_N(_0677_),
    .B(_0678_),
    .C(_0616_),
    .X(_0679_));
 sky130_fd_sc_hd__clkbuf_1 _1321_ (.A(_0679_),
    .X(_0066_));
 sky130_fd_sc_hd__nand2_1 _1322_ (.A(\send_divcnt[24] ),
    .B(_0677_),
    .Y(_0680_));
 sky130_fd_sc_hd__or2_1 _1323_ (.A(\send_divcnt[24] ),
    .B(_0677_),
    .X(_0681_));
 sky130_fd_sc_hd__and3_1 _1324_ (.A(_0514_),
    .B(_0680_),
    .C(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__clkbuf_1 _1325_ (.A(_0682_),
    .X(_0067_));
 sky130_fd_sc_hd__nor2_1 _1326_ (.A(_0466_),
    .B(_0680_),
    .Y(_0683_));
 sky130_fd_sc_hd__nand2_1 _1327_ (.A(_0466_),
    .B(_0680_),
    .Y(_0684_));
 sky130_fd_sc_hd__and3b_1 _1328_ (.A_N(_0683_),
    .B(_0684_),
    .C(_0616_),
    .X(_0685_));
 sky130_fd_sc_hd__clkbuf_1 _1329_ (.A(_0685_),
    .X(_0068_));
 sky130_fd_sc_hd__and4_1 _1330_ (.A(\send_divcnt[26] ),
    .B(\send_divcnt[25] ),
    .C(\send_divcnt[24] ),
    .D(_0677_),
    .X(_0686_));
 sky130_fd_sc_hd__or2_1 _1331_ (.A(\send_divcnt[26] ),
    .B(_0683_),
    .X(_0687_));
 sky130_fd_sc_hd__and3b_1 _1332_ (.A_N(_0686_),
    .B(_0687_),
    .C(_0616_),
    .X(_0688_));
 sky130_fd_sc_hd__clkbuf_1 _1333_ (.A(_0688_),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _1334_ (.A(\send_divcnt[27] ),
    .B(_0686_),
    .X(_0689_));
 sky130_fd_sc_hd__or2_1 _1335_ (.A(\send_divcnt[27] ),
    .B(_0686_),
    .X(_0690_));
 sky130_fd_sc_hd__and3b_1 _1336_ (.A_N(_0689_),
    .B(_0617_),
    .C(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__clkbuf_1 _1337_ (.A(_0691_),
    .X(_0070_));
 sky130_fd_sc_hd__and3_1 _1338_ (.A(\send_divcnt[28] ),
    .B(\send_divcnt[27] ),
    .C(_0686_),
    .X(_0692_));
 sky130_fd_sc_hd__or2_1 _1339_ (.A(\send_divcnt[28] ),
    .B(_0689_),
    .X(_0693_));
 sky130_fd_sc_hd__and3b_1 _1340_ (.A_N(_0692_),
    .B(_0617_),
    .C(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__clkbuf_1 _1341_ (.A(_0694_),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _1342_ (.A(\send_divcnt[29] ),
    .B(_0692_),
    .X(_0695_));
 sky130_fd_sc_hd__or2_1 _1343_ (.A(\send_divcnt[29] ),
    .B(_0692_),
    .X(_0696_));
 sky130_fd_sc_hd__and3b_1 _1344_ (.A_N(_0695_),
    .B(_0617_),
    .C(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__clkbuf_1 _1345_ (.A(_0697_),
    .X(_0072_));
 sky130_fd_sc_hd__or3b_2 _1346_ (.A(_0477_),
    .B(_0469_),
    .C_N(_0692_),
    .X(_0698_));
 sky130_fd_sc_hd__o211a_1 _1347_ (.A1(\send_divcnt[30] ),
    .A2(_0695_),
    .B1(_0698_),
    .C1(_0514_),
    .X(_0073_));
 sky130_fd_sc_hd__a2111oi_1 _1348_ (.A1(_0483_),
    .A2(_0698_),
    .B1(_0500_),
    .C1(_0495_),
    .D1(_0493_),
    .Y(_0699_));
 sky130_fd_sc_hd__o21a_1 _1349_ (.A1(_0483_),
    .A2(_0698_),
    .B1(_0699_),
    .X(_0074_));
 sky130_fd_sc_hd__clkbuf_4 _1350_ (.A(net47),
    .X(_0700_));
 sky130_fd_sc_hd__or2_1 _1351_ (.A(_0346_),
    .B(_0606_),
    .X(_0701_));
 sky130_fd_sc_hd__clkbuf_4 _1352_ (.A(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _1353_ (.A0(\recv_pattern[1] ),
    .A1(\recv_pattern[0] ),
    .S(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__and2_1 _1354_ (.A(_0700_),
    .B(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__clkbuf_1 _1355_ (.A(_0704_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _1356_ (.A0(\recv_pattern[2] ),
    .A1(\recv_pattern[1] ),
    .S(_0702_),
    .X(_0705_));
 sky130_fd_sc_hd__and2_1 _1357_ (.A(_0700_),
    .B(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__clkbuf_1 _1358_ (.A(_0706_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1359_ (.A0(\recv_pattern[3] ),
    .A1(\recv_pattern[2] ),
    .S(_0702_),
    .X(_0707_));
 sky130_fd_sc_hd__and2_1 _1360_ (.A(_0700_),
    .B(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__clkbuf_1 _1361_ (.A(_0708_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1362_ (.A0(\recv_pattern[4] ),
    .A1(\recv_pattern[3] ),
    .S(_0702_),
    .X(_0709_));
 sky130_fd_sc_hd__and2_1 _1363_ (.A(_0700_),
    .B(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__clkbuf_1 _1364_ (.A(_0710_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _1365_ (.A0(\recv_pattern[5] ),
    .A1(\recv_pattern[4] ),
    .S(_0702_),
    .X(_0711_));
 sky130_fd_sc_hd__and2_1 _1366_ (.A(_0700_),
    .B(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__clkbuf_1 _1367_ (.A(_0712_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _1368_ (.A0(\recv_pattern[6] ),
    .A1(\recv_pattern[5] ),
    .S(_0702_),
    .X(_0713_));
 sky130_fd_sc_hd__and2_1 _1369_ (.A(_0700_),
    .B(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__clkbuf_1 _1370_ (.A(_0714_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _1371_ (.A0(\recv_pattern[7] ),
    .A1(\recv_pattern[6] ),
    .S(_0702_),
    .X(_0715_));
 sky130_fd_sc_hd__and2_1 _1372_ (.A(_0700_),
    .B(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__clkbuf_1 _1373_ (.A(_0716_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _1374_ (.A0(net48),
    .A1(\recv_pattern[7] ),
    .S(_0702_),
    .X(_0717_));
 sky130_fd_sc_hd__and2_1 _1375_ (.A(_0700_),
    .B(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__clkbuf_1 _1376_ (.A(_0718_),
    .X(_0082_));
 sky130_fd_sc_hd__or3_1 _1377_ (.A(\recv_pattern[0] ),
    .B(_0219_),
    .C(_0347_),
    .X(_0719_));
 sky130_fd_sc_hd__o211a_1 _1378_ (.A1(\recv_buf_data[0] ),
    .A2(_0348_),
    .B1(_0719_),
    .C1(_0350_),
    .X(_0083_));
 sky130_fd_sc_hd__or3_1 _1379_ (.A(\recv_pattern[1] ),
    .B(_0219_),
    .C(_0347_),
    .X(_0720_));
 sky130_fd_sc_hd__o211a_1 _1380_ (.A1(\recv_buf_data[1] ),
    .A2(_0348_),
    .B1(_0720_),
    .C1(_0350_),
    .X(_0084_));
 sky130_fd_sc_hd__or3_1 _1381_ (.A(\recv_pattern[2] ),
    .B(_0219_),
    .C(_0347_),
    .X(_0721_));
 sky130_fd_sc_hd__o211a_1 _1382_ (.A1(\recv_buf_data[2] ),
    .A2(_0348_),
    .B1(_0721_),
    .C1(_0350_),
    .X(_0085_));
 sky130_fd_sc_hd__or3_1 _1383_ (.A(\recv_pattern[3] ),
    .B(_0219_),
    .C(_0347_),
    .X(_0722_));
 sky130_fd_sc_hd__o211a_1 _1384_ (.A1(\recv_buf_data[3] ),
    .A2(_0348_),
    .B1(_0722_),
    .C1(_0350_),
    .X(_0086_));
 sky130_fd_sc_hd__or3_1 _1385_ (.A(\recv_pattern[4] ),
    .B(_0219_),
    .C(_0347_),
    .X(_0723_));
 sky130_fd_sc_hd__o211a_1 _1386_ (.A1(\recv_buf_data[4] ),
    .A2(_0348_),
    .B1(_0723_),
    .C1(_0350_),
    .X(_0087_));
 sky130_fd_sc_hd__or3_1 _1387_ (.A(\recv_pattern[5] ),
    .B(_0219_),
    .C(_0347_),
    .X(_0724_));
 sky130_fd_sc_hd__o211a_1 _1388_ (.A1(\recv_buf_data[5] ),
    .A2(_0348_),
    .B1(_0724_),
    .C1(_0350_),
    .X(_0088_));
 sky130_fd_sc_hd__or3_1 _1389_ (.A(\recv_pattern[6] ),
    .B(_0219_),
    .C(_0347_),
    .X(_0725_));
 sky130_fd_sc_hd__o211a_1 _1390_ (.A1(\recv_buf_data[6] ),
    .A2(_0348_),
    .B1(_0725_),
    .C1(_0351_),
    .X(_0089_));
 sky130_fd_sc_hd__or3_1 _1391_ (.A(\recv_pattern[7] ),
    .B(_0219_),
    .C(_0347_),
    .X(_0726_));
 sky130_fd_sc_hd__o211a_1 _1392_ (.A1(\recv_buf_data[7] ),
    .A2(_0348_),
    .B1(_0726_),
    .C1(_0351_),
    .X(_0090_));
 sky130_fd_sc_hd__and2_1 _1393_ (.A(_0596_),
    .B(_0598_),
    .X(_0727_));
 sky130_fd_sc_hd__o211a_2 _1394_ (.A1(_0525_),
    .A2(_0727_),
    .B1(_0702_),
    .C1(net47),
    .X(_0728_));
 sky130_fd_sc_hd__buf_4 _1395_ (.A(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__and2b_1 _1396_ (.A_N(\recv_divcnt[0] ),
    .B(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__clkbuf_1 _1397_ (.A(_0730_),
    .X(_0091_));
 sky130_fd_sc_hd__or2_1 _1398_ (.A(\recv_divcnt[1] ),
    .B(\recv_divcnt[0] ),
    .X(_0731_));
 sky130_fd_sc_hd__nand2_1 _1399_ (.A(\recv_divcnt[1] ),
    .B(\recv_divcnt[0] ),
    .Y(_0732_));
 sky130_fd_sc_hd__and3_1 _1400_ (.A(_0729_),
    .B(_0731_),
    .C(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__clkbuf_1 _1401_ (.A(_0733_),
    .X(_0092_));
 sky130_fd_sc_hd__nor2_1 _1402_ (.A(_0341_),
    .B(_0732_),
    .Y(_0734_));
 sky130_fd_sc_hd__clkbuf_4 _1403_ (.A(_0728_),
    .X(_0735_));
 sky130_fd_sc_hd__nand2_1 _1404_ (.A(_0341_),
    .B(_0732_),
    .Y(_0736_));
 sky130_fd_sc_hd__and3b_1 _1405_ (.A_N(_0734_),
    .B(_0735_),
    .C(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__clkbuf_1 _1406_ (.A(_0737_),
    .X(_0093_));
 sky130_fd_sc_hd__and4_2 _1407_ (.A(\recv_divcnt[3] ),
    .B(\recv_divcnt[2] ),
    .C(\recv_divcnt[1] ),
    .D(\recv_divcnt[0] ),
    .X(_0738_));
 sky130_fd_sc_hd__or2_1 _1408_ (.A(\recv_divcnt[3] ),
    .B(_0734_),
    .X(_0739_));
 sky130_fd_sc_hd__clkbuf_4 _1409_ (.A(_0728_),
    .X(_0740_));
 sky130_fd_sc_hd__and3b_1 _1410_ (.A_N(_0738_),
    .B(_0739_),
    .C(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__clkbuf_1 _1411_ (.A(_0741_),
    .X(_0094_));
 sky130_fd_sc_hd__nand2_1 _1412_ (.A(\recv_divcnt[4] ),
    .B(_0738_),
    .Y(_0742_));
 sky130_fd_sc_hd__or2_1 _1413_ (.A(\recv_divcnt[4] ),
    .B(_0738_),
    .X(_0743_));
 sky130_fd_sc_hd__and3_1 _1414_ (.A(_0729_),
    .B(_0742_),
    .C(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__clkbuf_1 _1415_ (.A(_0744_),
    .X(_0095_));
 sky130_fd_sc_hd__and3_1 _1416_ (.A(\recv_divcnt[5] ),
    .B(\recv_divcnt[4] ),
    .C(_0738_),
    .X(_0745_));
 sky130_fd_sc_hd__a21o_1 _1417_ (.A1(\recv_divcnt[4] ),
    .A2(_0738_),
    .B1(\recv_divcnt[5] ),
    .X(_0746_));
 sky130_fd_sc_hd__and3b_1 _1418_ (.A_N(_0745_),
    .B(_0746_),
    .C(_0740_),
    .X(_0747_));
 sky130_fd_sc_hd__clkbuf_1 _1419_ (.A(_0747_),
    .X(_0096_));
 sky130_fd_sc_hd__and4_1 _1420_ (.A(\recv_divcnt[6] ),
    .B(\recv_divcnt[5] ),
    .C(\recv_divcnt[4] ),
    .D(_0738_),
    .X(_0748_));
 sky130_fd_sc_hd__or2_1 _1421_ (.A(\recv_divcnt[6] ),
    .B(_0745_),
    .X(_0749_));
 sky130_fd_sc_hd__and3b_1 _1422_ (.A_N(_0748_),
    .B(_0749_),
    .C(_0740_),
    .X(_0750_));
 sky130_fd_sc_hd__clkbuf_1 _1423_ (.A(_0750_),
    .X(_0097_));
 sky130_fd_sc_hd__nand2_1 _1424_ (.A(\recv_divcnt[7] ),
    .B(_0748_),
    .Y(_0751_));
 sky130_fd_sc_hd__or2_1 _1425_ (.A(\recv_divcnt[7] ),
    .B(_0748_),
    .X(_0752_));
 sky130_fd_sc_hd__and3_1 _1426_ (.A(_0729_),
    .B(_0751_),
    .C(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__clkbuf_1 _1427_ (.A(_0753_),
    .X(_0098_));
 sky130_fd_sc_hd__nor2_1 _1428_ (.A(_0261_),
    .B(_0751_),
    .Y(_0754_));
 sky130_fd_sc_hd__nand2_1 _1429_ (.A(_0261_),
    .B(_0751_),
    .Y(_0755_));
 sky130_fd_sc_hd__and3b_1 _1430_ (.A_N(_0754_),
    .B(_0755_),
    .C(_0740_),
    .X(_0756_));
 sky130_fd_sc_hd__clkbuf_1 _1431_ (.A(_0756_),
    .X(_0099_));
 sky130_fd_sc_hd__and4_1 _1432_ (.A(\recv_divcnt[9] ),
    .B(\recv_divcnt[8] ),
    .C(\recv_divcnt[7] ),
    .D(_0748_),
    .X(_0757_));
 sky130_fd_sc_hd__or2_1 _1433_ (.A(\recv_divcnt[9] ),
    .B(_0754_),
    .X(_0758_));
 sky130_fd_sc_hd__and3b_1 _1434_ (.A_N(_0757_),
    .B(_0758_),
    .C(_0740_),
    .X(_0759_));
 sky130_fd_sc_hd__clkbuf_1 _1435_ (.A(_0759_),
    .X(_0100_));
 sky130_fd_sc_hd__nand2_1 _1436_ (.A(\recv_divcnt[10] ),
    .B(_0757_),
    .Y(_0760_));
 sky130_fd_sc_hd__or2_1 _1437_ (.A(\recv_divcnt[10] ),
    .B(_0757_),
    .X(_0761_));
 sky130_fd_sc_hd__and3_1 _1438_ (.A(_0729_),
    .B(_0760_),
    .C(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__clkbuf_1 _1439_ (.A(_0762_),
    .X(_0101_));
 sky130_fd_sc_hd__nor2_1 _1440_ (.A(_0277_),
    .B(_0760_),
    .Y(_0763_));
 sky130_fd_sc_hd__nand2_1 _1441_ (.A(_0277_),
    .B(_0760_),
    .Y(_0764_));
 sky130_fd_sc_hd__and3b_1 _1442_ (.A_N(_0763_),
    .B(_0764_),
    .C(_0740_),
    .X(_0765_));
 sky130_fd_sc_hd__clkbuf_1 _1443_ (.A(_0765_),
    .X(_0102_));
 sky130_fd_sc_hd__and4_1 _1444_ (.A(\recv_divcnt[12] ),
    .B(\recv_divcnt[11] ),
    .C(\recv_divcnt[10] ),
    .D(_0757_),
    .X(_0766_));
 sky130_fd_sc_hd__or2_1 _1445_ (.A(\recv_divcnt[12] ),
    .B(_0763_),
    .X(_0767_));
 sky130_fd_sc_hd__and3b_1 _1446_ (.A_N(_0766_),
    .B(_0767_),
    .C(_0740_),
    .X(_0768_));
 sky130_fd_sc_hd__clkbuf_1 _1447_ (.A(_0768_),
    .X(_0103_));
 sky130_fd_sc_hd__and2_1 _1448_ (.A(\recv_divcnt[13] ),
    .B(_0766_),
    .X(_0131_));
 sky130_fd_sc_hd__or2_1 _1449_ (.A(\recv_divcnt[13] ),
    .B(_0766_),
    .X(_0132_));
 sky130_fd_sc_hd__and3b_1 _1450_ (.A_N(_0131_),
    .B(_0132_),
    .C(_0740_),
    .X(_0133_));
 sky130_fd_sc_hd__clkbuf_1 _1451_ (.A(_0133_),
    .X(_0104_));
 sky130_fd_sc_hd__and3_1 _1452_ (.A(\recv_divcnt[14] ),
    .B(\recv_divcnt[13] ),
    .C(_0766_),
    .X(_0134_));
 sky130_fd_sc_hd__or2_1 _1453_ (.A(\recv_divcnt[14] ),
    .B(_0131_),
    .X(_0135_));
 sky130_fd_sc_hd__and3b_1 _1454_ (.A_N(_0134_),
    .B(_0135_),
    .C(_0740_),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_1 _1455_ (.A(_0136_),
    .X(_0105_));
 sky130_fd_sc_hd__and4_1 _1456_ (.A(\recv_divcnt[15] ),
    .B(\recv_divcnt[14] ),
    .C(\recv_divcnt[13] ),
    .D(_0766_),
    .X(_0137_));
 sky130_fd_sc_hd__or2_1 _1457_ (.A(\recv_divcnt[15] ),
    .B(_0134_),
    .X(_0138_));
 sky130_fd_sc_hd__and3b_1 _1458_ (.A_N(_0137_),
    .B(_0138_),
    .C(_0740_),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_1 _1459_ (.A(_0139_),
    .X(_0106_));
 sky130_fd_sc_hd__nand2_1 _1460_ (.A(\recv_divcnt[16] ),
    .B(_0137_),
    .Y(_0140_));
 sky130_fd_sc_hd__or2_1 _1461_ (.A(\recv_divcnt[16] ),
    .B(_0137_),
    .X(_0141_));
 sky130_fd_sc_hd__and3_1 _1462_ (.A(_0729_),
    .B(_0140_),
    .C(_0141_),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _1463_ (.A(_0142_),
    .X(_0107_));
 sky130_fd_sc_hd__nor2_1 _1464_ (.A(_0301_),
    .B(_0302_),
    .Y(_0143_));
 sky130_fd_sc_hd__and2_1 _1465_ (.A(_0137_),
    .B(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__nand2_1 _1466_ (.A(_0301_),
    .B(_0140_),
    .Y(_0145_));
 sky130_fd_sc_hd__and3b_1 _1467_ (.A_N(_0144_),
    .B(_0735_),
    .C(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _1468_ (.A(_0146_),
    .X(_0108_));
 sky130_fd_sc_hd__and3_1 _1469_ (.A(\recv_divcnt[18] ),
    .B(_0137_),
    .C(_0143_),
    .X(_0147_));
 sky130_fd_sc_hd__or2_1 _1470_ (.A(\recv_divcnt[18] ),
    .B(_0144_),
    .X(_0148_));
 sky130_fd_sc_hd__and3b_1 _1471_ (.A_N(_0147_),
    .B(_0735_),
    .C(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_1 _1472_ (.A(_0149_),
    .X(_0109_));
 sky130_fd_sc_hd__and4_1 _1473_ (.A(\recv_divcnt[19] ),
    .B(\recv_divcnt[18] ),
    .C(_0137_),
    .D(_0143_),
    .X(_0150_));
 sky130_fd_sc_hd__or2_1 _1474_ (.A(\recv_divcnt[19] ),
    .B(_0147_),
    .X(_0151_));
 sky130_fd_sc_hd__and3b_1 _1475_ (.A_N(_0150_),
    .B(_0151_),
    .C(_0728_),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_1 _1476_ (.A(_0152_),
    .X(_0110_));
 sky130_fd_sc_hd__or2_1 _1477_ (.A(\recv_divcnt[20] ),
    .B(_0150_),
    .X(_0153_));
 sky130_fd_sc_hd__nand2_1 _1478_ (.A(\recv_divcnt[20] ),
    .B(_0150_),
    .Y(_0154_));
 sky130_fd_sc_hd__and3_1 _1479_ (.A(_0729_),
    .B(_0153_),
    .C(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__clkbuf_1 _1480_ (.A(_0155_),
    .X(_0111_));
 sky130_fd_sc_hd__nand2_1 _1481_ (.A(_0316_),
    .B(_0154_),
    .Y(_0156_));
 sky130_fd_sc_hd__or2_1 _1482_ (.A(_0316_),
    .B(_0154_),
    .X(_0157_));
 sky130_fd_sc_hd__and3_1 _1483_ (.A(_0729_),
    .B(_0156_),
    .C(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_1 _1484_ (.A(_0158_),
    .X(_0112_));
 sky130_fd_sc_hd__and4_1 _1485_ (.A(\recv_divcnt[22] ),
    .B(\recv_divcnt[21] ),
    .C(\recv_divcnt[20] ),
    .D(_0150_),
    .X(_0159_));
 sky130_fd_sc_hd__nand2_1 _1486_ (.A(_0312_),
    .B(_0157_),
    .Y(_0160_));
 sky130_fd_sc_hd__and3b_1 _1487_ (.A_N(_0159_),
    .B(_0735_),
    .C(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__clkbuf_1 _1488_ (.A(_0161_),
    .X(_0113_));
 sky130_fd_sc_hd__or2_1 _1489_ (.A(\recv_divcnt[23] ),
    .B(_0159_),
    .X(_0162_));
 sky130_fd_sc_hd__nand2_1 _1490_ (.A(\recv_divcnt[23] ),
    .B(_0159_),
    .Y(_0163_));
 sky130_fd_sc_hd__and3_1 _1491_ (.A(_0729_),
    .B(_0162_),
    .C(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_1 _1492_ (.A(_0164_),
    .X(_0114_));
 sky130_fd_sc_hd__nor2_1 _1493_ (.A(_0297_),
    .B(_0163_),
    .Y(_0165_));
 sky130_fd_sc_hd__nand2_1 _1494_ (.A(_0297_),
    .B(_0163_),
    .Y(_0166_));
 sky130_fd_sc_hd__and3b_1 _1495_ (.A_N(_0165_),
    .B(_0166_),
    .C(_0728_),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_1 _1496_ (.A(_0167_),
    .X(_0115_));
 sky130_fd_sc_hd__and4_1 _1497_ (.A(\recv_divcnt[25] ),
    .B(\recv_divcnt[24] ),
    .C(\recv_divcnt[23] ),
    .D(_0159_),
    .X(_0168_));
 sky130_fd_sc_hd__or2_1 _1498_ (.A(\recv_divcnt[25] ),
    .B(_0165_),
    .X(_0169_));
 sky130_fd_sc_hd__and3b_1 _1499_ (.A_N(_0168_),
    .B(_0735_),
    .C(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_1 _1500_ (.A(_0170_),
    .X(_0116_));
 sky130_fd_sc_hd__or2_1 _1501_ (.A(\recv_divcnt[26] ),
    .B(_0168_),
    .X(_0171_));
 sky130_fd_sc_hd__nand2_1 _1502_ (.A(\recv_divcnt[26] ),
    .B(_0168_),
    .Y(_0172_));
 sky130_fd_sc_hd__and3_1 _1503_ (.A(_0729_),
    .B(_0171_),
    .C(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__clkbuf_1 _1504_ (.A(_0173_),
    .X(_0117_));
 sky130_fd_sc_hd__and3_1 _1505_ (.A(\recv_divcnt[27] ),
    .B(\recv_divcnt[26] ),
    .C(_0168_),
    .X(_0174_));
 sky130_fd_sc_hd__a21o_1 _1506_ (.A1(\recv_divcnt[26] ),
    .A2(_0168_),
    .B1(\recv_divcnt[27] ),
    .X(_0175_));
 sky130_fd_sc_hd__and3b_1 _1507_ (.A_N(_0174_),
    .B(_0735_),
    .C(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__clkbuf_1 _1508_ (.A(_0176_),
    .X(_0118_));
 sky130_fd_sc_hd__or2_1 _1509_ (.A(\recv_divcnt[28] ),
    .B(_0174_),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_1 _1510_ (.A(\recv_divcnt[28] ),
    .B(_0174_),
    .Y(_0178_));
 sky130_fd_sc_hd__and3_1 _1511_ (.A(_0735_),
    .B(_0177_),
    .C(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__clkbuf_1 _1512_ (.A(_0179_),
    .X(_0119_));
 sky130_fd_sc_hd__and3_1 _1513_ (.A(\recv_divcnt[29] ),
    .B(\recv_divcnt[28] ),
    .C(_0174_),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_1 _1514_ (.A(_0220_),
    .B(_0178_),
    .Y(_0181_));
 sky130_fd_sc_hd__and3b_1 _1515_ (.A_N(_0180_),
    .B(_0735_),
    .C(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__clkbuf_1 _1516_ (.A(_0182_),
    .X(_0120_));
 sky130_fd_sc_hd__and4_1 _1517_ (.A(\recv_divcnt[30] ),
    .B(\recv_divcnt[29] ),
    .C(\recv_divcnt[28] ),
    .D(_0174_),
    .X(_0183_));
 sky130_fd_sc_hd__or2_1 _1518_ (.A(\recv_divcnt[30] ),
    .B(_0180_),
    .X(_0184_));
 sky130_fd_sc_hd__and3b_1 _1519_ (.A_N(_0183_),
    .B(_0735_),
    .C(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__clkbuf_1 _1520_ (.A(_0185_),
    .X(_0121_));
 sky130_fd_sc_hd__or2_1 _1521_ (.A(\recv_divcnt[31] ),
    .B(_0183_),
    .X(_0186_));
 sky130_fd_sc_hd__nand2_1 _1522_ (.A(\recv_divcnt[31] ),
    .B(_0183_),
    .Y(_0187_));
 sky130_fd_sc_hd__and3_1 _1523_ (.A(_0735_),
    .B(_0186_),
    .C(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_1 _1524_ (.A(_0188_),
    .X(_0122_));
 sky130_fd_sc_hd__o21ai_1 _1525_ (.A1(net43),
    .A2(_0239_),
    .B1(_0351_),
    .Y(_0189_));
 sky130_fd_sc_hd__a21o_1 _1526_ (.A1(net43),
    .A2(net11),
    .B1(_0189_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _1527_ (.A0(net93),
    .A1(net22),
    .S(net43),
    .X(_0190_));
 sky130_fd_sc_hd__and2_1 _1528_ (.A(_0700_),
    .B(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__clkbuf_1 _1529_ (.A(_0191_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _1530_ (.A0(net104),
    .A1(net33),
    .S(net43),
    .X(_0192_));
 sky130_fd_sc_hd__and2_1 _1531_ (.A(_0700_),
    .B(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__clkbuf_1 _1532_ (.A(_0193_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _1533_ (.A0(net107),
    .A1(net36),
    .S(net43),
    .X(_0194_));
 sky130_fd_sc_hd__and2_1 _1534_ (.A(_0349_),
    .B(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__clkbuf_1 _1535_ (.A(_0195_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _1536_ (.A0(net108),
    .A1(net37),
    .S(net43),
    .X(_0196_));
 sky130_fd_sc_hd__and2_1 _1537_ (.A(_0349_),
    .B(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_1 _1538_ (.A(_0197_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _1539_ (.A0(net109),
    .A1(net38),
    .S(net43),
    .X(_0198_));
 sky130_fd_sc_hd__and2_1 _1540_ (.A(_0349_),
    .B(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_1 _1541_ (.A(_0199_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _1542_ (.A0(net110),
    .A1(net39),
    .S(net43),
    .X(_0200_));
 sky130_fd_sc_hd__and2_1 _1543_ (.A(_0349_),
    .B(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_1 _1544_ (.A(_0201_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _1545_ (.A0(net111),
    .A1(net40),
    .S(net43),
    .X(_0202_));
 sky130_fd_sc_hd__and2_1 _1546_ (.A(_0349_),
    .B(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_1 _1547_ (.A(_0203_),
    .X(_0130_));
 sky130_fd_sc_hd__dfxtp_1 _1548_ (.CLK(clknet_4_15_0_clk),
    .D(_0000_),
    .Q(recv_buf_valid));
 sky130_fd_sc_hd__dfxtp_4 _1549_ (.CLK(clknet_4_5_0_clk),
    .D(_0001_),
    .Q(net112));
 sky130_fd_sc_hd__dfxtp_4 _1550_ (.CLK(clknet_4_5_0_clk),
    .D(_0002_),
    .Q(net113));
 sky130_fd_sc_hd__dfxtp_2 _1551_ (.CLK(clknet_4_5_0_clk),
    .D(_0003_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_2 _1552_ (.CLK(clknet_4_5_0_clk),
    .D(_0004_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_2 _1553_ (.CLK(clknet_4_7_0_clk),
    .D(_0005_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_4 _1554_ (.CLK(clknet_4_7_0_clk),
    .D(_0006_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_4 _1555_ (.CLK(clknet_4_7_0_clk),
    .D(_0007_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_4 _1556_ (.CLK(clknet_4_7_0_clk),
    .D(_0008_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_4 _1557_ (.CLK(clknet_4_7_0_clk),
    .D(_0009_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_4 _1558_ (.CLK(clknet_4_7_0_clk),
    .D(_0010_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_4 _1559_ (.CLK(clknet_4_6_0_clk),
    .D(_0011_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_4 _1560_ (.CLK(clknet_4_7_0_clk),
    .D(_0012_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_2 _1561_ (.CLK(clknet_4_7_0_clk),
    .D(_0013_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_2 _1562_ (.CLK(clknet_4_7_0_clk),
    .D(_0014_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_2 _1563_ (.CLK(clknet_4_13_0_clk),
    .D(_0015_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_2 _1564_ (.CLK(clknet_4_13_0_clk),
    .D(_0016_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_2 _1565_ (.CLK(clknet_4_13_0_clk),
    .D(_0017_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_2 _1566_ (.CLK(clknet_4_13_0_clk),
    .D(_0018_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_2 _1567_ (.CLK(clknet_4_13_0_clk),
    .D(_0019_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_2 _1568_ (.CLK(clknet_4_12_0_clk),
    .D(_0020_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_2 _1569_ (.CLK(clknet_4_13_0_clk),
    .D(_0021_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_2 _1570_ (.CLK(clknet_4_12_0_clk),
    .D(_0022_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_2 _1571_ (.CLK(clknet_4_13_0_clk),
    .D(_0023_),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_2 _1572_ (.CLK(clknet_4_13_0_clk),
    .D(_0024_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_4 _1573_ (.CLK(clknet_4_9_0_clk),
    .D(_0025_),
    .Q(net114));
 sky130_fd_sc_hd__dfxtp_1 _1574_ (.CLK(clknet_4_11_0_clk),
    .D(_0026_),
    .Q(\send_pattern[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1575_ (.CLK(clknet_4_12_0_clk),
    .D(_0027_),
    .Q(\send_pattern[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1576_ (.CLK(clknet_4_13_0_clk),
    .D(_0028_),
    .Q(\send_pattern[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1577_ (.CLK(clknet_4_13_0_clk),
    .D(_0029_),
    .Q(\send_pattern[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1578_ (.CLK(clknet_4_13_0_clk),
    .D(_0030_),
    .Q(\send_pattern[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1579_ (.CLK(clknet_4_15_0_clk),
    .D(_0031_),
    .Q(\send_pattern[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1580_ (.CLK(clknet_4_15_0_clk),
    .D(_0032_),
    .Q(\send_pattern[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1581_ (.CLK(clknet_4_15_0_clk),
    .D(_0033_),
    .Q(\send_pattern[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1582_ (.CLK(clknet_4_11_0_clk),
    .D(_0034_),
    .Q(\send_bitcnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1583_ (.CLK(clknet_4_11_0_clk),
    .D(_0035_),
    .Q(\send_bitcnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1584_ (.CLK(clknet_4_14_0_clk),
    .D(_0036_),
    .Q(\send_bitcnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1585_ (.CLK(clknet_4_14_0_clk),
    .D(_0037_),
    .Q(\send_bitcnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1586_ (.CLK(clknet_4_15_0_clk),
    .D(_0038_),
    .Q(send_dummy));
 sky130_fd_sc_hd__dfxtp_2 _1587_ (.CLK(clknet_4_11_0_clk),
    .D(_0039_),
    .Q(\recv_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1588_ (.CLK(clknet_4_10_0_clk),
    .D(_0040_),
    .Q(\recv_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1589_ (.CLK(clknet_4_10_0_clk),
    .D(_0041_),
    .Q(\recv_state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1590_ (.CLK(clknet_4_10_0_clk),
    .D(_0042_),
    .Q(\recv_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1591_ (.CLK(clknet_4_5_0_clk),
    .D(_0043_),
    .Q(\send_divcnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1592_ (.CLK(clknet_4_5_0_clk),
    .D(_0044_),
    .Q(\send_divcnt[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1593_ (.CLK(clknet_4_4_0_clk),
    .D(_0045_),
    .Q(\send_divcnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1594_ (.CLK(clknet_4_4_0_clk),
    .D(_0046_),
    .Q(\send_divcnt[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1595_ (.CLK(clknet_4_4_0_clk),
    .D(_0047_),
    .Q(\send_divcnt[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1596_ (.CLK(clknet_4_1_0_clk),
    .D(_0048_),
    .Q(\send_divcnt[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1597_ (.CLK(clknet_4_1_0_clk),
    .D(_0049_),
    .Q(\send_divcnt[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1598_ (.CLK(clknet_4_1_0_clk),
    .D(_0050_),
    .Q(\send_divcnt[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1599_ (.CLK(clknet_4_0_0_clk),
    .D(_0051_),
    .Q(\send_divcnt[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1600_ (.CLK(clknet_4_0_0_clk),
    .D(_0052_),
    .Q(\send_divcnt[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1601_ (.CLK(clknet_4_0_0_clk),
    .D(_0053_),
    .Q(\send_divcnt[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1602_ (.CLK(clknet_4_0_0_clk),
    .D(_0054_),
    .Q(\send_divcnt[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1603_ (.CLK(clknet_4_0_0_clk),
    .D(_0055_),
    .Q(\send_divcnt[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1604_ (.CLK(clknet_4_0_0_clk),
    .D(_0056_),
    .Q(\send_divcnt[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1605_ (.CLK(clknet_4_2_0_clk),
    .D(_0057_),
    .Q(\send_divcnt[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1606_ (.CLK(clknet_4_2_0_clk),
    .D(_0058_),
    .Q(\send_divcnt[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1607_ (.CLK(clknet_4_2_0_clk),
    .D(_0059_),
    .Q(\send_divcnt[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1608_ (.CLK(clknet_4_2_0_clk),
    .D(_0060_),
    .Q(\send_divcnt[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1609_ (.CLK(clknet_4_2_0_clk),
    .D(_0061_),
    .Q(\send_divcnt[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1610_ (.CLK(clknet_4_2_0_clk),
    .D(_0062_),
    .Q(\send_divcnt[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1611_ (.CLK(clknet_4_8_0_clk),
    .D(_0063_),
    .Q(\send_divcnt[20] ));
 sky130_fd_sc_hd__dfxtp_2 _1612_ (.CLK(clknet_4_8_0_clk),
    .D(_0064_),
    .Q(\send_divcnt[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1613_ (.CLK(clknet_4_8_0_clk),
    .D(_0065_),
    .Q(\send_divcnt[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1614_ (.CLK(clknet_4_8_0_clk),
    .D(_0066_),
    .Q(\send_divcnt[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1615_ (.CLK(clknet_4_8_0_clk),
    .D(_0067_),
    .Q(\send_divcnt[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1616_ (.CLK(clknet_4_9_0_clk),
    .D(_0068_),
    .Q(\send_divcnt[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1617_ (.CLK(clknet_4_8_0_clk),
    .D(_0069_),
    .Q(\send_divcnt[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1618_ (.CLK(clknet_4_10_0_clk),
    .D(_0070_),
    .Q(\send_divcnt[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1619_ (.CLK(clknet_4_10_0_clk),
    .D(_0071_),
    .Q(\send_divcnt[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1620_ (.CLK(clknet_4_10_0_clk),
    .D(_0072_),
    .Q(\send_divcnt[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1621_ (.CLK(clknet_4_10_0_clk),
    .D(_0073_),
    .Q(\send_divcnt[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1622_ (.CLK(clknet_4_11_0_clk),
    .D(_0074_),
    .Q(\send_divcnt[31] ));
 sky130_fd_sc_hd__dfxtp_1 _1623_ (.CLK(clknet_4_14_0_clk),
    .D(_0075_),
    .Q(\recv_pattern[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1624_ (.CLK(clknet_4_14_0_clk),
    .D(_0076_),
    .Q(\recv_pattern[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1625_ (.CLK(clknet_4_14_0_clk),
    .D(_0077_),
    .Q(\recv_pattern[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1626_ (.CLK(clknet_4_14_0_clk),
    .D(_0078_),
    .Q(\recv_pattern[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1627_ (.CLK(clknet_4_14_0_clk),
    .D(_0079_),
    .Q(\recv_pattern[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1628_ (.CLK(clknet_4_14_0_clk),
    .D(_0080_),
    .Q(\recv_pattern[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1629_ (.CLK(clknet_4_11_0_clk),
    .D(_0081_),
    .Q(\recv_pattern[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1630_ (.CLK(clknet_4_11_0_clk),
    .D(_0082_),
    .Q(\recv_pattern[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1631_ (.CLK(clknet_4_14_0_clk),
    .D(_0083_),
    .Q(\recv_buf_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1632_ (.CLK(clknet_4_15_0_clk),
    .D(_0084_),
    .Q(\recv_buf_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1633_ (.CLK(clknet_4_15_0_clk),
    .D(_0085_),
    .Q(\recv_buf_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1634_ (.CLK(clknet_4_15_0_clk),
    .D(_0086_),
    .Q(\recv_buf_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1635_ (.CLK(clknet_4_15_0_clk),
    .D(_0087_),
    .Q(\recv_buf_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1636_ (.CLK(clknet_4_15_0_clk),
    .D(_0088_),
    .Q(\recv_buf_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1637_ (.CLK(clknet_4_15_0_clk),
    .D(_0089_),
    .Q(\recv_buf_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1638_ (.CLK(clknet_4_15_0_clk),
    .D(_0090_),
    .Q(\recv_buf_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1639_ (.CLK(clknet_4_6_0_clk),
    .D(_0091_),
    .Q(\recv_divcnt[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1640_ (.CLK(clknet_4_6_0_clk),
    .D(_0092_),
    .Q(\recv_divcnt[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1641_ (.CLK(clknet_4_6_0_clk),
    .D(_0093_),
    .Q(\recv_divcnt[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1642_ (.CLK(clknet_4_6_0_clk),
    .D(_0094_),
    .Q(\recv_divcnt[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1643_ (.CLK(clknet_4_4_0_clk),
    .D(_0095_),
    .Q(\recv_divcnt[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1644_ (.CLK(clknet_4_4_0_clk),
    .D(_0096_),
    .Q(\recv_divcnt[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1645_ (.CLK(clknet_4_4_0_clk),
    .D(_0097_),
    .Q(\recv_divcnt[6] ));
 sky130_fd_sc_hd__dfxtp_2 _1646_ (.CLK(clknet_4_4_0_clk),
    .D(_0098_),
    .Q(\recv_divcnt[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1647_ (.CLK(clknet_4_4_0_clk),
    .D(_0099_),
    .Q(\recv_divcnt[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1648_ (.CLK(clknet_4_1_0_clk),
    .D(_0100_),
    .Q(\recv_divcnt[9] ));
 sky130_fd_sc_hd__dfxtp_2 _1649_ (.CLK(clknet_4_1_0_clk),
    .D(_0101_),
    .Q(\recv_divcnt[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1650_ (.CLK(clknet_4_0_0_clk),
    .D(_0102_),
    .Q(\recv_divcnt[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1651_ (.CLK(clknet_4_3_0_clk),
    .D(_0103_),
    .Q(\recv_divcnt[12] ));
 sky130_fd_sc_hd__dfxtp_2 _1652_ (.CLK(clknet_4_2_0_clk),
    .D(_0104_),
    .Q(\recv_divcnt[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1653_ (.CLK(clknet_4_2_0_clk),
    .D(_0105_),
    .Q(\recv_divcnt[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1654_ (.CLK(clknet_4_3_0_clk),
    .D(_0106_),
    .Q(\recv_divcnt[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1655_ (.CLK(clknet_4_3_0_clk),
    .D(_0107_),
    .Q(\recv_divcnt[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1656_ (.CLK(clknet_4_3_0_clk),
    .D(_0108_),
    .Q(\recv_divcnt[17] ));
 sky130_fd_sc_hd__dfxtp_2 _1657_ (.CLK(clknet_4_3_0_clk),
    .D(_0109_),
    .Q(\recv_divcnt[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1658_ (.CLK(clknet_4_3_0_clk),
    .D(_0110_),
    .Q(\recv_divcnt[19] ));
 sky130_fd_sc_hd__dfxtp_2 _1659_ (.CLK(clknet_4_6_0_clk),
    .D(_0111_),
    .Q(\recv_divcnt[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1660_ (.CLK(clknet_4_12_0_clk),
    .D(_0112_),
    .Q(\recv_divcnt[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1661_ (.CLK(clknet_4_12_0_clk),
    .D(_0113_),
    .Q(\recv_divcnt[22] ));
 sky130_fd_sc_hd__dfxtp_2 _1662_ (.CLK(clknet_4_3_0_clk),
    .D(_0114_),
    .Q(\recv_divcnt[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1663_ (.CLK(clknet_4_9_0_clk),
    .D(_0115_),
    .Q(\recv_divcnt[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1664_ (.CLK(clknet_4_8_0_clk),
    .D(_0116_),
    .Q(\recv_divcnt[25] ));
 sky130_fd_sc_hd__dfxtp_2 _1665_ (.CLK(clknet_4_8_0_clk),
    .D(_0117_),
    .Q(\recv_divcnt[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1666_ (.CLK(clknet_4_9_0_clk),
    .D(_0118_),
    .Q(\recv_divcnt[27] ));
 sky130_fd_sc_hd__dfxtp_2 _1667_ (.CLK(clknet_4_12_0_clk),
    .D(_0119_),
    .Q(\recv_divcnt[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1668_ (.CLK(clknet_4_9_0_clk),
    .D(_0120_),
    .Q(\recv_divcnt[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1669_ (.CLK(clknet_4_12_0_clk),
    .D(_0121_),
    .Q(\recv_divcnt[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1670_ (.CLK(clknet_4_12_0_clk),
    .D(_0122_),
    .Q(\recv_divcnt[31] ));
 sky130_fd_sc_hd__dfxtp_1 _1671_ (.CLK(clknet_4_5_0_clk),
    .D(_0123_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_2 _1672_ (.CLK(clknet_4_5_0_clk),
    .D(_0124_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_2 _1673_ (.CLK(clknet_4_4_0_clk),
    .D(_0125_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_2 _1674_ (.CLK(clknet_4_5_0_clk),
    .D(_0126_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_2 _1675_ (.CLK(clknet_4_5_0_clk),
    .D(_0127_),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_4 _1676_ (.CLK(clknet_4_5_0_clk),
    .D(_0128_),
    .Q(net109));
 sky130_fd_sc_hd__dfxtp_2 _1677_ (.CLK(clknet_4_5_0_clk),
    .D(_0129_),
    .Q(net110));
 sky130_fd_sc_hd__dfxtp_4 _1678_ (.CLK(clknet_4_5_0_clk),
    .D(_0130_),
    .Q(net111));
 sky130_fd_sc_hd__clkbuf_1 _1679_ (.A(net73),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _1680_ (.A(net73),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _1681_ (.A(net73),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _1682_ (.A(net73),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 _1683_ (.A(net73),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _1684_ (.A(net73),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 _1685_ (.A(net73),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 _1686_ (.A(net73),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 _1687_ (.A(net73),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 _1688_ (.A(net73),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 _1689_ (.A(net73),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _1690_ (.A(net73),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 _1691_ (.A(net73),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _1692_ (.A(net73),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _1693_ (.A(net73),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _1694_ (.A(net73),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _1695_ (.A(net73),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _1696_ (.A(net73),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _1697_ (.A(net73),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _1698_ (.A(net73),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _1699_ (.A(net73),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _1700_ (.A(net73),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _1701_ (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2785 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(reg_dat_di[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(reg_dat_di[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(reg_dat_di[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(reg_dat_di[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(reg_dat_di[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(reg_dat_di[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(reg_dat_di[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(reg_dat_di[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(reg_dat_re),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(reg_dat_we),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(reg_div_di[0]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(reg_div_di[10]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(reg_div_di[11]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(reg_div_di[12]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(reg_div_di[13]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(reg_div_di[14]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(reg_div_di[15]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(reg_div_di[16]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(reg_div_di[17]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(reg_div_di[18]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(reg_div_di[19]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(reg_div_di[1]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(reg_div_di[20]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(reg_div_di[21]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(reg_div_di[22]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(reg_div_di[23]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(reg_div_di[24]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(reg_div_di[25]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(reg_div_di[26]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(reg_div_di[27]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(reg_div_di[28]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(reg_div_di[29]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(reg_div_di[2]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(reg_div_di[30]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(reg_div_di[31]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(reg_div_di[3]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(reg_div_di[4]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(reg_div_di[5]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(reg_div_di[6]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(reg_div_di[7]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(reg_div_di[8]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(reg_div_di[9]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 input43 (.A(reg_div_we[0]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 input44 (.A(reg_div_we[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(reg_div_we[2]),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(reg_div_we[3]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(resetn),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(ser_rx),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net49),
    .X(reg_dat_do[0]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net50),
    .X(reg_dat_do[10]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net51),
    .X(reg_dat_do[11]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net52),
    .X(reg_dat_do[12]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net53),
    .X(reg_dat_do[13]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net54),
    .X(reg_dat_do[14]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .X(reg_dat_do[15]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(reg_dat_do[16]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(reg_dat_do[17]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(reg_dat_do[18]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(reg_dat_do[19]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(reg_dat_do[1]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(reg_dat_do[20]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .X(reg_dat_do[21]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net63),
    .X(reg_dat_do[22]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net64),
    .X(reg_dat_do[23]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net65),
    .X(reg_dat_do[24]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(reg_dat_do[25]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(reg_dat_do[26]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(reg_dat_do[27]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .X(reg_dat_do[28]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(reg_dat_do[29]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .X(reg_dat_do[2]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .X(reg_dat_do[30]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .X(reg_dat_do[31]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net74),
    .X(reg_dat_do[3]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .X(reg_dat_do[4]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net76),
    .X(reg_dat_do[5]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net77),
    .X(reg_dat_do[6]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net78),
    .X(reg_dat_do[7]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net79),
    .X(reg_dat_do[8]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net80),
    .X(reg_dat_do[9]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net81),
    .X(reg_dat_wait));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net82),
    .X(reg_div_do[0]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net83),
    .X(reg_div_do[10]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net84),
    .X(reg_div_do[11]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net85),
    .X(reg_div_do[12]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net86),
    .X(reg_div_do[13]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net87),
    .X(reg_div_do[14]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net88),
    .X(reg_div_do[15]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net89),
    .X(reg_div_do[16]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net90),
    .X(reg_div_do[17]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net91),
    .X(reg_div_do[18]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net92),
    .X(reg_div_do[19]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net93),
    .X(reg_div_do[1]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net94),
    .X(reg_div_do[20]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net95),
    .X(reg_div_do[21]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net96),
    .X(reg_div_do[22]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net97),
    .X(reg_div_do[23]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net98),
    .X(reg_div_do[24]));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net99),
    .X(reg_div_do[25]));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net100),
    .X(reg_div_do[26]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net101),
    .X(reg_div_do[27]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net102),
    .X(reg_div_do[28]));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net103),
    .X(reg_div_do[29]));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net104),
    .X(reg_div_do[2]));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net105),
    .X(reg_div_do[30]));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net106),
    .X(reg_div_do[31]));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net107),
    .X(reg_div_do[3]));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net108),
    .X(reg_div_do[4]));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net109),
    .X(reg_div_do[5]));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net110),
    .X(reg_div_do[6]));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net111),
    .X(reg_div_do[7]));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net112),
    .X(reg_div_do[8]));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net113),
    .X(reg_div_do[9]));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net114),
    .X(ser_tx));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__D (.DIODE(_0150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__B (.DIODE(_0150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__B (.DIODE(_0150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1475__A_N (.DIODE(_0150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__D (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__C (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1510__B (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__B (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__A_N (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__A (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__B2 (.DIODE(_0246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__A1 (.DIODE(_0246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__A (.DIODE(_0246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1020__A (.DIODE(_0246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0825__A1 (.DIODE(_0246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__A (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1048__A (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1002__A1 (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0897__A1 (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0889__A (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__A (.DIODE(_0315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__A (.DIODE(_0315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__A1 (.DIODE(_0315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1002__B2 (.DIODE(_0315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0892__A1 (.DIODE(_0315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__A1 (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__A1 (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1063__A1 (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1050__A1 (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__B2 (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0897__B2 (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__A (.DIODE(_0320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1056__A1 (.DIODE(_0320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__A (.DIODE(_0320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__A (.DIODE(_0320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1351__A (.DIODE(_0346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0922__A (.DIODE(_0346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1391__C (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__C (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1387__C (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__C (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1383__C (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1381__C (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1379__C (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1377__C (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__A1 (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0923__B (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1546__A (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1543__A (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__A (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__A (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__A (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1226__A (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__A (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0940__A (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0927__A (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0925__A (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1388__C1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1386__C1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1384__C1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1382__C1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__C1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1378__C1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1138__B1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1135__B1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1132__B1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__B1 (.DIODE(_0350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__B1 (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__C1 (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1390__C1 (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1221__B1 (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1215__C1 (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1124__A1 (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__A (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0935__A (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0932__A (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0929__A (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1092__A1 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1348__D1 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1131__S (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__A2 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1112__A2 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__A2 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__A2 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__A2 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1104__A2 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__A2 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1101__A2 (.DIODE(_0493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1348__B1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__A (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__C1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1112__C1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__C1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__C1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__C1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1104__C1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__C1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1101__C1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__C1 (.DIODE(_0509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__C1 (.DIODE(_0509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1228__B (.DIODE(_0509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__A2 (.DIODE(_0509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1347__C1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1324__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1312__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1293__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1258__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1246__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1231__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1124__B1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1138__A2 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1332__C (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1328__C (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1320__C (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1316__C (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1308__C (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1304__C (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1300__C (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1289__C (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1281__C (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1237__A (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1344__B (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1340__B (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1336__B (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1277__C (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1273__C (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1262__C (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1254__C (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1250__C (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1242__C (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1238__C (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1528__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1375__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1369__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1366__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1363__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1360__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1357__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1354__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__B1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1371__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1368__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1365__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1356__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1353__S (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__C (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1475__C (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__A (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1403__A (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1395__A (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1503__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1479__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1438__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1426__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1414__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1400__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__A (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__B (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1515__B (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__A (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__B (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1499__B (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__B (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1471__B (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1467__B (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__B (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1458__C (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1454__C (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1450__C (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1446__C (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__C (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__C (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1430__C (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1422__C (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1418__C (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1410__C (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1136__B (.DIODE(send_dummy));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__A (.DIODE(send_dummy));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__A (.DIODE(send_dummy));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1533__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1530__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1526__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1136__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1137__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__0972__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__0968__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__0962__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__0956__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__0953__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1136__C (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__0993__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__0987__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__C1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__1350__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__0971__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1701__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1700__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1696__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1694__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1692__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1691__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1689__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1686__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1684__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1683__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1681__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1680__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1679__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0780__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0776__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__A_N (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0814__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0934__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0853__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0845__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1180__A_N (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0941__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0833__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__1006__B2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0944__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0842__B2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0832__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__1184__A_N (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__B2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__1006__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0947__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0842__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0830__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__A_N (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0950__A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__A_N (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0953__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1054__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1044__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0956__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0882__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__1058__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__1053__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0906__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0885__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__1158__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__1156__C1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__1058__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__1055__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0962__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0884__B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0881__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__B_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__0813__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1156__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__0895__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__0881__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0968__A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0907__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0894__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0892__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0972__A0 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0908__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0893__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__0890__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0909__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0888__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__A0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1145__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1081__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__A0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__0987__A0 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0802__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1208__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1073__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1070__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0993__A0 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0802__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0800__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__1530__A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__A_N (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__B_N (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1089__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__A0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1210__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__A0 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1533__A0 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1166__A_N (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__A0 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0807__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0806__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__A0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0827__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0824__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0821__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__A0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1019__B2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0804__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__B_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1174__A_N (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1019__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0928__A0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0849__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1190__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0931__A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0844__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1101__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1599__CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1600__CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1601__CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1602__CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1603__CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1604__CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1650__CLK (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1605__CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1606__CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1608__CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1652__CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1653__CLK (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1651__CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1654__CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1655__CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1656__CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1657__CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1658__CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1662__CLK (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1593__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1595__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1645__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1647__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__CLK (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1549__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1551__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1592__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1671__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1672__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1674__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1675__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1676__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1677__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1678__CLK (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1613__CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1614__CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1615__CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1664__CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1665__CLK (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1616__CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1663__CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1666__CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1668__CLK (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1574__CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__CLK (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1568__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1570__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1660__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1661__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1667__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1669__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1670__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1564__CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1566__CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1571__CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1576__CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1578__CLK (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1626__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1628__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__CLK (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1580__CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1586__CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1632__CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1633__CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1635__CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1636__CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1638__CLK (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net93));
endmodule
