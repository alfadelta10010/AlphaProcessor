* NGSPICE file created from simpleuart.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt simpleuart VGND VPWR clk reg_dat_di[0] reg_dat_di[10] reg_dat_di[11] reg_dat_di[12]
+ reg_dat_di[13] reg_dat_di[14] reg_dat_di[15] reg_dat_di[16] reg_dat_di[17] reg_dat_di[18]
+ reg_dat_di[19] reg_dat_di[1] reg_dat_di[20] reg_dat_di[21] reg_dat_di[22] reg_dat_di[23]
+ reg_dat_di[24] reg_dat_di[25] reg_dat_di[26] reg_dat_di[27] reg_dat_di[28] reg_dat_di[29]
+ reg_dat_di[2] reg_dat_di[30] reg_dat_di[31] reg_dat_di[3] reg_dat_di[4] reg_dat_di[5]
+ reg_dat_di[6] reg_dat_di[7] reg_dat_di[8] reg_dat_di[9] reg_dat_do[0] reg_dat_do[10]
+ reg_dat_do[11] reg_dat_do[12] reg_dat_do[13] reg_dat_do[14] reg_dat_do[15] reg_dat_do[16]
+ reg_dat_do[17] reg_dat_do[18] reg_dat_do[19] reg_dat_do[1] reg_dat_do[20] reg_dat_do[21]
+ reg_dat_do[22] reg_dat_do[23] reg_dat_do[24] reg_dat_do[25] reg_dat_do[26] reg_dat_do[27]
+ reg_dat_do[28] reg_dat_do[29] reg_dat_do[2] reg_dat_do[30] reg_dat_do[31] reg_dat_do[3]
+ reg_dat_do[4] reg_dat_do[5] reg_dat_do[6] reg_dat_do[7] reg_dat_do[8] reg_dat_do[9]
+ reg_dat_re reg_dat_wait reg_dat_we reg_div_di[0] reg_div_di[10] reg_div_di[11] reg_div_di[12]
+ reg_div_di[13] reg_div_di[14] reg_div_di[15] reg_div_di[16] reg_div_di[17] reg_div_di[18]
+ reg_div_di[19] reg_div_di[1] reg_div_di[20] reg_div_di[21] reg_div_di[22] reg_div_di[23]
+ reg_div_di[24] reg_div_di[25] reg_div_di[26] reg_div_di[27] reg_div_di[28] reg_div_di[29]
+ reg_div_di[2] reg_div_di[30] reg_div_di[31] reg_div_di[3] reg_div_di[4] reg_div_di[5]
+ reg_div_di[6] reg_div_di[7] reg_div_di[8] reg_div_di[9] reg_div_do[0] reg_div_do[10]
+ reg_div_do[11] reg_div_do[12] reg_div_do[13] reg_div_do[14] reg_div_do[15] reg_div_do[16]
+ reg_div_do[17] reg_div_do[18] reg_div_do[19] reg_div_do[1] reg_div_do[20] reg_div_do[21]
+ reg_div_do[22] reg_div_do[23] reg_div_do[24] reg_div_do[25] reg_div_do[26] reg_div_do[27]
+ reg_div_do[28] reg_div_do[29] reg_div_do[2] reg_div_do[30] reg_div_do[31] reg_div_do[3]
+ reg_div_do[4] reg_div_do[5] reg_div_do[6] reg_div_do[7] reg_div_do[8] reg_div_do[9]
+ reg_div_we[0] reg_div_we[1] reg_div_we[2] reg_div_we[3] resetn ser_rx ser_tx
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0965__A0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1534__A _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0956__A0 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1270_ _0408_ _0637_ _0641_ _0509_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0985_ _0381_ _0390_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0947__A0 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1606_ clknet_4_2_0_clk _0058_ VGND VGND VPWR VPWR send_divcnt\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__1354__A _0700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1537_ _0349_ _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__and2_1
X_1468_ _0146_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__1124__B1 _0514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1399_ recv_divcnt\[1\] recv_divcnt\[0\] VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1430__C _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0770_ send_dummy send_bitcnt\[3\] _0204_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__or3_1
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1322_ send_divcnt\[24\] _0677_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1253_ send_divcnt\[6\] _0625_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_88_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1184_ net87 recv_divcnt\[13\] VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
X_0968_ net95 net24 net45 VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0899_ _0299_ _0308_ _0323_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1250__C _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0822_ recv_divcnt\[6\] VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1592__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1305_ _0667_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1236_ _0513_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1167_ net104 recv_divcnt\[1\] VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1098_ send_dummy _0491_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_670 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1022__A_N net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1021_ send_divcnt\[5\] VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_818 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0805_ _0229_ recv_divcnt\[7\] VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1219_ _0600_ _0602_ _0603_ _0497_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_140_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_595 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1539__A0 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1537__A _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ clknet_4_12_0_clk _0022_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output86_A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1630__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1004_ send_divcnt\[12\] _0258_ net86 _0403_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_122_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1357__A _0700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1699_ net73 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1653__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput64 net64 VGND VGND VPWR VPWR reg_dat_do[23] sky130_fd_sc_hd__clkbuf_1
Xoutput53 net53 VGND VGND VPWR VPWR reg_dat_do[13] sky130_fd_sc_hd__clkbuf_1
Xoutput75 net75 VGND VGND VPWR VPWR reg_dat_do[4] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput97 net97 VGND VGND VPWR VPWR reg_div_do[23] sky130_fd_sc_hd__clkbuf_1
Xoutput86 net86 VGND VGND VPWR VPWR reg_div_do[13] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1622_ clknet_4_11_0_clk _0074_ VGND VGND VPWR VPWR send_divcnt\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1553_ clknet_4_7_0_clk _0005_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_120_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1484_ _0158_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1676__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_782 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1549__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0804__A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0984_ net100 net29 net46 VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1605_ clknet_4_2_0_clk _0057_ VGND VGND VPWR VPWR send_divcnt\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1536_ net108 net37 net43 VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1467_ _0144_ _0735_ _0145_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__and3b_1
XANTENNA__1124__A1 _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1398_ recv_divcnt\[1\] recv_divcnt\[0\] VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_718 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_782 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1348__D1 _0493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1321_ _0679_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1252_ send_divcnt\[6\] send_divcnt\[5\] send_divcnt\[4\] _0619_ VGND VGND VPWR VPWR
+ _0628_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_88_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1190__A net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1183_ net88 recv_divcnt\[14\] VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_746 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0967_ _0378_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0898_ _0311_ _0318_ _0322_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1519_ _0183_ _0735_ _0184_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__and3b_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0821_ net110 VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__clkinv_2
XFILLER_0_24_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1304_ _0665_ _0666_ _0616_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__and3b_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1235_ _0613_ _0611_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1166_ net107 recv_divcnt\[2\] VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__and2b_1
XFILLER_0_126_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1097_ net47 VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1020_ _0246_ send_divcnt\[6\] VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0804_ net111 VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1218_ recv_state\[1\] recv_state\[0\] _0527_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1149_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1582__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ send_divcnt\[13\] VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0807__A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1698_ net73 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput65 net65 VGND VGND VPWR VPWR reg_dat_do[24] sky130_fd_sc_hd__clkbuf_1
Xoutput54 net54 VGND VGND VPWR VPWR reg_dat_do[14] sky130_fd_sc_hd__clkbuf_1
Xoutput76 net76 VGND VGND VPWR VPWR reg_dat_do[5] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput98 net98 VGND VGND VPWR VPWR reg_div_do[24] sky130_fd_sc_hd__clkbuf_1
Xoutput87 net87 VGND VGND VPWR VPWR reg_div_do[14] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_19_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1621_ clknet_4_10_0_clk _0073_ VGND VGND VPWR VPWR send_divcnt\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1384__C1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1552_ clknet_4_5_0_clk _0004_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dfxtp_2
X_1483_ _0729_ _0156_ _0157_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1185__A_N net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_780 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0910__A net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0892__A1 _0315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0892__B2 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0983_ _0389_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1604_ clknet_4_0_0_clk _0056_ VGND VGND VPWR VPWR send_divcnt\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1535_ _0195_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1466_ _0301_ _0140_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1397_ _0730_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1643__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1098__A send_dummy VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1320_ _0677_ _0678_ _0616_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_9_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_775 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1251_ _0627_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1106__A2 _0493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1182_ _0565_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1666__CLK clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_96_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_758 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0966_ _0360_ _0377_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0897_ _0313_ recv_divcnt\[23\] recv_divcnt\[21\] _0319_ _0321_ VGND VGND VPWR VPWR
+ _0322_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1518_ recv_divcnt\[30\] _0180_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1449_ recv_divcnt\[13\] _0766_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1033__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0820_ _0231_ recv_divcnt\[5\] VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1303_ send_divcnt\[19\] _0662_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__or2_1
X_1234_ _0613_ _0611_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1165_ recv_divcnt\[1\] net104 VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__or2b_1
XFILLER_0_149_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1096_ _0492_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__nor2_4
XFILLER_0_149_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0949_ _0366_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_803 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1006__B2 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1006__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0803_ _0225_ _0227_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1217_ recv_state\[3\] _0601_ _0599_ _0217_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1148_ net98 recv_divcnt\[23\] VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1079_ net105 _0477_ _0478_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1002_ _0313_ send_divcnt\[23\] send_divcnt\[22\] _0315_ VGND VGND VPWR VPWR _0402_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1697_ net73 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0968__A0 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput66 net66 VGND VGND VPWR VPWR reg_dat_do[25] sky130_fd_sc_hd__clkbuf_1
Xoutput55 net55 VGND VGND VPWR VPWR reg_dat_do[15] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput77 net77 VGND VGND VPWR VPWR reg_dat_do[6] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput99 net99 VGND VGND VPWR VPWR reg_div_do[25] sky130_fd_sc_hd__clkbuf_1
Xoutput88 net88 VGND VGND VPWR VPWR reg_div_do[15] sky130_fd_sc_hd__clkbuf_1
XANTENNA__0908__A net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0959__A0 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1620_ clknet_4_10_0_clk _0072_ VGND VGND VPWR VPWR send_divcnt\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output91_A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1551_ clknet_4_5_0_clk _0003_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dfxtp_2
X_1482_ _0316_ _0154_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1572__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_116_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0982_ _0381_ _0388_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_143_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_662 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1595__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1603_ clknet_4_0_0_clk _0055_ VGND VGND VPWR VPWR send_divcnt\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1534_ _0349_ _0194_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__and2_1
X_1465_ _0137_ _0143_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1396_ recv_divcnt\[0\] _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1348__B1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1250_ _0625_ _0626_ _0617_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__and3b_1
XANTENNA__1471__B _0735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1181_ _0270_ recv_divcnt\[10\] recv_divcnt\[9\] _0268_ _0566_ VGND VGND VPWR VPWR
+ _0567_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_91_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_478 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0965_ net94 net23 net45 VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0896_ _0320_ recv_divcnt\[20\] VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1517_ recv_divcnt\[30\] recv_divcnt\[29\] recv_divcnt\[28\] _0174_ VGND VGND VPWR
+ VPWR _0183_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1448_ recv_divcnt\[13\] _0766_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__and2_1
XANTENNA__1610__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1379_ recv_pattern\[1\] _0219_ _0347_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1633__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1302_ send_divcnt\[19\] send_divcnt\[18\] _0661_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__and3_1
X_1233_ send_divcnt\[2\] VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1164_ _0541_ _0542_ _0547_ _0549_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__o31a_1
XFILLER_0_149_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1095_ _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0948_ _0360_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0879_ recv_divcnt\[20\] VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1656__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0802_ net103 _0220_ _0226_ net102 VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_643 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1216_ recv_state\[2\] VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1147_ net97 _0312_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1078_ _0222_ send_divcnt\[31\] VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0990__S net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1172__A1 _0246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1163__A1 _0319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ _0401_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1696_ net73 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1154__A1 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput67 net67 VGND VGND VPWR VPWR reg_dat_do[26] sky130_fd_sc_hd__clkbuf_1
Xoutput56 net56 VGND VGND VPWR VPWR reg_dat_do[16] sky130_fd_sc_hd__clkbuf_1
Xoutput78 net78 VGND VGND VPWR VPWR reg_dat_do[7] sky130_fd_sc_hd__clkbuf_1
XANTENNA__1145__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput89 net89 VGND VGND VPWR VPWR reg_div_do[16] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0924__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1458__C _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1550_ clknet_4_5_0_clk _0002_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dfxtp_4
XANTENNA_output84_A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1481_ _0316_ _0154_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1679_ net73 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0981_ net99 net28 net46 VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_674 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1602_ clknet_4_0_0_clk _0054_ VGND VGND VPWR VPWR send_divcnt\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1533_ net107 net36 net43 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__mux2_1
X_1464_ _0301_ _0302_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1395_ _0728_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__buf_4
XFILLER_0_38_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1395__A _0728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1180_ net85 recv_divcnt\[11\] VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_88_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_696 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0964_ _0376_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0895_ net94 VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_132_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1516_ _0182_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1447_ _0768_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__1381__C _0347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1378_ recv_buf_data\[0\] _0348_ _0719_ _0350_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_52_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0993__S net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1585__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0932__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_814 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_858 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1301_ _0664_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
X_1232_ _0612_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
X_1163_ _0319_ recv_divcnt\[20\] _0536_ _0535_ _0548_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1094_ net10 _0491_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_482 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0947_ net87 net16 net44 VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0878_ net90 _0301_ _0302_ net89 VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0927__A _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_747 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0801_ recv_divcnt\[28\] VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1477__B _0150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1600__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1215_ recv_state\[0\] _0527_ _0600_ _0351_ _0219_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_79_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1146_ _0313_ recv_divcnt\[22\] VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1077_ send_divcnt\[30\] VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1623__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1000_ _0381_ _0400_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1695_ net73 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_9_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1646__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1129_ send_bitcnt\[1\] send_bitcnt\[0\] send_bitcnt\[2\] VGND VGND VPWR VPWR _0518_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1090__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1090__B2 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1378__C1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_783 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput57 net57 VGND VGND VPWR VPWR reg_dat_do[17] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput68 net68 VGND VGND VPWR VPWR reg_dat_do[27] sky130_fd_sc_hd__clkbuf_1
Xoutput79 net79 VGND VGND VPWR VPWR reg_dat_do[8] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1081__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0940__A _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ _0155_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1669__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1678_ clknet_4_5_0_clk _0130_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_4
XANTENNA__1681__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0996__S net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1063__A1 _0319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1530__S net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0935__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0980_ _0387_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1601_ clknet_4_0_0_clk _0053_ VGND VGND VPWR VPWR send_divcnt\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1532_ _0193_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1463_ _0142_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1394_ _0525_ _0727_ _0702_ net47 VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__o211a_2
XFILLER_0_38_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0845__A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1379__C _0347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_723 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1289__C _0616_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_528 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0963_ _0360_ _0375_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0894_ net95 VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__clkinv_2
XFILLER_0_3_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_859 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1515_ _0180_ _0735_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__and3b_1
XFILLER_0_10_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1446_ _0766_ _0767_ _0740_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__and3b_1
X_1377_ recv_pattern\[0\] _0219_ _0347_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_74_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1009__B2 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_9 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1300_ _0662_ _0663_ _0616_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__and3b_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1231_ _0514_ _0610_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__and3_1
X_1162_ _0319_ recv_divcnt\[20\] _0537_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1093_ _0492_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0946_ _0364_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0877_ recv_divcnt\[16\] VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0931__A0 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1429_ _0261_ _0751_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1552__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0800_ net103 _0220_ _0221_ _0223_ _0224_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_862 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1214_ recv_state\[0\] _0599_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_148_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1145_ net100 _0296_ _0528_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1076_ _0283_ send_divcnt\[28\] VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_5_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0853__A net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1387__C _0347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0999__S net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_667 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1684__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0929_ _0351_ _0352_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1575__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_784 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1533__S net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0938__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1694_ net73 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1679__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1128_ _0517_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1059_ _0446_ _0447_ _0450_ _0458_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput58 net58 VGND VGND VPWR VPWR reg_dat_do[18] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput69 net69 VGND VGND VPWR VPWR reg_dat_do[28] sky130_fd_sc_hd__clkbuf_1
XANTENNA__1353__S _0702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1677_ clknet_4_5_0_clk _0129_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1613__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_13_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output108_A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_526 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1600_ clknet_4_0_0_clk _0052_ VGND VGND VPWR VPWR send_divcnt\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1636__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1531_ _0700_ _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__and2_1
X_1462_ _0729_ _0140_ _0141_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1393_ _0596_ _0598_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_121_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0861__A net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_130_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1692__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0962_ net92 net21 net45 VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0893_ net96 _0312_ _0314_ _0317_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1514_ _0220_ _0178_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1445_ recv_divcnt\[12\] _0763_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__or2_1
X_1376_ _0718_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1687__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1536__S net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1230_ send_divcnt\[1\] send_divcnt\[0\] VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__nand2_1
X_1161_ net91 _0301_ _0543_ _0544_ _0546_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__o2111a_1
X_1092_ _0465_ _0482_ _0490_ _0478_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0945_ _0360_ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0876_ recv_divcnt\[17\] VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__clkinv_2
XFILLER_0_15_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_149_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1428_ _0261_ _0751_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1359_ recv_pattern\[3\] recv_pattern\[2\] _0702_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1356__S _0702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1175__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1213_ _0596_ _0598_ _0527_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_144_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1144_ _0288_ recv_divcnt\[26\] _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1075_ _0288_ send_divcnt\[27\] VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0928_ net112 net41 net44 VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0859_ _0283_ recv_divcnt\[28\] VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1157__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1157__B2 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1693_ net73 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1127_ _0349_ _0515_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1058_ net92 _0451_ _0452_ net91 _0457_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1695__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput59 net59 VGND VGND VPWR VPWR reg_dat_do[19] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1565__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1499__B _0735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1676_ clknet_4_5_0_clk _0128_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_1_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1539__S net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1485__D _0150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1530_ net104 net33 net43 VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output82_A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1461_ recv_divcnt\[16\] _0137_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1392_ recv_buf_data\[7\] _0348_ _0726_ _0351_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1659_ clknet_4_6_0_clk _0111_ VGND VGND VPWR VPWR recv_divcnt\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_611 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1359__S _0702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0961_ _0374_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_119_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1603__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0892_ _0315_ recv_divcnt\[22\] _0316_ net95 VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1513_ recv_divcnt\[29\] recv_divcnt\[28\] _0174_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__and3_1
X_1444_ recv_divcnt\[12\] recv_divcnt\[11\] recv_divcnt\[10\] _0757_ VGND VGND VPWR
+ VPWR _0766_ sky130_fd_sc_hd__and4_1
X_1375_ _0700_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_52_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_706 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_774 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1626__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_728 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1118__A _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1160_ _0541_ _0545_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_129_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1091_ send_bitcnt\[3\] _0204_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__nor2_2
XFILLER_0_99_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1102__C1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0944_ net86 net15 net44 VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0875_ net89 VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1427_ _0753_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
X_1358_ _0706_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
X_1289_ _0654_ _0655_ _0616_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__and3b_1
XFILLER_0_78_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1698__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_886 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_864 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1212_ net106 _0336_ _0597_ recv_state\[0\] VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_144_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1143_ _0283_ recv_divcnt\[27\] VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__and2_1
X_1074_ _0473_ send_divcnt\[29\] VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0927_ _0349_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0858_ net102 VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0789_ _0214_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_89_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1692_ net73 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1126_ send_bitcnt\[1\] _0511_ _0508_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__nand3_1
XFILLER_0_79_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1057_ _0453_ send_divcnt\[18\] send_divcnt\[17\] _0454_ _0456_ VGND VGND VPWR VPWR
+ _0457_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput49 net49 VGND VGND VPWR VPWR reg_dat_do[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0774__B net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0790__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_696 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_44_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1675_ clknet_4_5_0_clk _0127_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0875__A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1109_ send_pattern\[4\] _0496_ _0504_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1460_ recv_divcnt\[16\] _0137_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__nand2_1
X_1391_ recv_pattern\[7\] _0219_ _0347_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_26_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1202__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1202__B2 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1658_ clknet_4_3_0_clk _0110_ VGND VGND VPWR VPWR recv_divcnt\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_44_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1589_ clknet_4_10_0_clk _0041_ VGND VGND VPWR VPWR recv_state\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_623 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output113_A net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0960_ _0360_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_136_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0891_ recv_divcnt\[21\] VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1512_ _0179_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1443_ _0765_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
X_1374_ net48 recv_pattern\[7\] _0702_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1578__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_786 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0934__A0 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0782__B net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1090_ net106 _0483_ _0477_ net105 _0489_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1300__C _0616_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0943_ _0362_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0874_ _0285_ _0293_ _0295_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__or4b_1
XFILLER_0_3_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1426_ _0729_ _0751_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__and3_1
X_1357_ _0700_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1044__A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1288_ send_divcnt\[14\] _0648_ send_divcnt\[15\] VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1211_ _0525_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_144_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1142_ _0283_ recv_divcnt\[27\] recv_divcnt\[26\] _0288_ VGND VGND VPWR VPWR _0528_
+ sky130_fd_sc_hd__o22a_1
X_1073_ net103 VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_615 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0926_ _0215_ _0348_ _0350_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_754 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0857_ _0256_ _0265_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0788_ recv_buf_data\[7\] net73 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1616__CLK clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1409_ _0728_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_67_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_807 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1691_ net73 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1125_ _0511_ _0508_ send_bitcnt\[1\] VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_49_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1056_ _0320_ send_divcnt\[20\] send_divcnt\[19\] _0455_ VGND VGND VPWR VPWR _0456_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_146_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0909_ net97 _0328_ _0318_ _0332_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1674_ clknet_4_5_0_clk _0126_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1108_ send_pattern\[5\] _0493_ _0495_ net4 _0500_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1039_ _0258_ send_divcnt\[12\] _0437_ _0438_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1137__A net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1390_ recv_buf_data\[6\] _0348_ _0725_ _0351_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1047__A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1657_ clknet_4_3_0_clk _0109_ VGND VGND VPWR VPWR recv_divcnt\[18\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1588_ clknet_4_10_0_clk _0040_ VGND VGND VPWR VPWR recv_state\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_668 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0796__A net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output106_A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ net96 VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__clkinv_2
XFILLER_0_55_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_808 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1511_ _0735_ _0177_ _0178_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1442_ _0763_ _0764_ _0740_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__and3b_1
X_1373_ _0716_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1187__B2 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_498 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1672__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1150__A _0315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0942_ _0360_ _0361_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0873_ net99 _0296_ _0297_ net98 VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1425_ recv_divcnt\[7\] _0748_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__or2_1
X_1356_ recv_pattern\[2\] recv_pattern\[1\] _0702_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1287_ send_divcnt\[15\] send_divcnt\[14\] _0648_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0907__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1210_ net106 _0336_ _0591_ _0594_ _0595_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_144_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1141_ _0347_ _0525_ _0526_ net48 VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__a22oi_2
XANTENNA__1568__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1072_ _0222_ send_divcnt\[31\] send_divcnt\[30\] _0335_ _0471_ VGND VGND VPWR VPWR
+ _0472_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0925_ _0349_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0856_ _0255_ _0267_ _0280_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__or3_1
XFILLER_0_140_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0787_ _0213_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1055__A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1408_ recv_divcnt\[3\] _0734_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1339_ send_divcnt\[28\] _0689_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__or2_1
XANTENNA__0894__A net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0788__B net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1690_ net73 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output98_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1124_ _0351_ _0205_ _0512_ _0514_ send_bitcnt\[0\] VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__a32o_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1055_ net92 VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0908_ net96 _0312_ _0314_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0889__A _0313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0839_ recv_divcnt\[13\] VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1526__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1606__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1673_ clknet_4_4_0_clk _0125_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_123_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1107_ send_pattern\[3\] _0496_ _0503_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1038_ net88 _0436_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1629__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_690 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1380__C1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1656_ clknet_4_3_0_clk _0108_ VGND VGND VPWR VPWR recv_divcnt\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1587_ clknet_4_11_0_clk _0039_ VGND VGND VPWR VPWR recv_state\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_622 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1510__B _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1114__C1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1701__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1148__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1510_ recv_divcnt\[28\] _0174_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1441_ _0277_ _0760_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1372_ _0700_ _0715_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_52_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1639_ clknet_4_6_0_clk _0091_ VGND VGND VPWR VPWR recv_divcnt\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1102__A2 _0493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0941_ net85 net14 net44 VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0872_ recv_divcnt\[24\] VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1424_ recv_divcnt\[7\] _0748_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__nand2_1
X_1355_ _0704_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1286_ _0653_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_786 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1426__A _0729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1140_ recv_state\[0\] _0525_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_144_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1071_ _0288_ send_divcnt\[27\] _0468_ net100 _0470_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0924_ net47 VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_836 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0855_ _0273_ _0279_ _0259_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0786_ recv_buf_data\[6\] net73 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1407_ recv_divcnt\[3\] recv_divcnt\[2\] recv_divcnt\[1\] recv_divcnt\[0\] VGND VGND
+ VPWR VPWR _0738_ sky130_fd_sc_hd__and4_2
XFILLER_0_39_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1338_ send_divcnt\[28\] send_divcnt\[27\] _0686_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1269_ send_divcnt\[8\] send_divcnt\[7\] _0628_ _0640_ VGND VGND VPWR VPWR _0641_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_78_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1662__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0825__A1 _0246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_49_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1002__B2 _0315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1002__A1 _0313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1246__A _0514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_58_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1123_ _0513_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_49_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1054_ net90 VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0907_ net95 _0316_ _0321_ _0331_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0838_ _0256_ _0259_ _0262_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__or3b_1
XFILLER_0_141_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0769_ send_bitcnt\[2\] send_bitcnt\[1\] send_bitcnt\[0\] VGND VGND VPWR VPWR _0204_
+ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_77_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_859 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_583 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1672_ clknet_4_5_0_clk _0124_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1106_ send_pattern\[4\] _0493_ _0495_ net3 _0500_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_37_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1037_ net88 _0436_ _0405_ net87 VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_672 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_615 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1132__B1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1655_ clknet_4_3_0_clk _0107_ VGND VGND VPWR VPWR recv_divcnt\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1586_ clknet_4_15_0_clk _0038_ VGND VGND VPWR VPWR send_dummy sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_634 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0937__A0 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0928__A0 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1440_ _0277_ _0760_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__nor2_1
XANTENNA_output73_A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1371_ recv_pattern\[7\] recv_pattern\[6\] _0702_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1638_ clknet_4_15_0_clk _0090_ VGND VGND VPWR VPWR recv_buf_data\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1569_ clknet_4_13_0_clk _0021_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_6_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output111_A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0940_ _0349_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0871_ recv_divcnt\[25\] VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__inv_2
XANTENNA__1159__A net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1423_ _0750_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
X_1354_ _0700_ _0703_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__and2_1
X_1285_ _0514_ _0651_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_69_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1591__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ send_divcnt\[28\] _0283_ net103 _0469_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0923_ _0219_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__nor2_4
XFILLER_0_83_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0854_ net84 _0277_ _0262_ _0272_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0785_ _0212_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1336__B _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1406_ _0737_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
X_1337_ _0691_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1268_ _0408_ _0413_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1199_ _0543_ _0549_ _0546_ _0584_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_643 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1122_ _0497_ _0508_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1053_ net91 VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0906_ net91 _0329_ _0309_ _0330_ _0306_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__o311a_1
XFILLER_0_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0837_ net113 _0260_ _0261_ net112 VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1513__C _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_595 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_554 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_727 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_532 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1671_ clknet_4_5_0_clk _0123_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1652__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1105_ send_pattern\[2\] _0496_ _0502_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_37_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1036_ send_divcnt\[15\] VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_86_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1141__A1 _0347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1141__B2 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1540__A _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1675__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1418__C _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1328__C _0616_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1654_ clknet_4_3_0_clk _0106_ VGND VGND VPWR VPWR recv_divcnt\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1585_ clknet_4_14_0_clk _0037_ VGND VGND VPWR VPWR send_bitcnt\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1344__B _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1360__A _0700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1548__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ net112 _0411_ _0412_ net111 _0418_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__o221a_1
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1519__B _0735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1238__C _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_579 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1370_ _0714_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1637_ clknet_4_15_0_clk _0089_ VGND VGND VPWR VPWR recv_buf_data\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1568_ clknet_4_12_0_clk _0020_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_6_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1499_ _0168_ _0735_ _0169_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_87_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output104_A net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ _0294_ recv_divcnt\[24\] VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1422_ _0748_ _0749_ _0740_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__and3b_1
X_1353_ recv_pattern\[1\] recv_pattern\[0\] _0702_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__mux2_1
X_1284_ send_divcnt\[14\] _0648_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_69_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0953__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0999_ net106 net35 net46 VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1609__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0922_ _0346_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0853_ net83 _0271_ recv_divcnt\[10\] VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__or3b_1
XFILLER_0_43_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0784_ recv_buf_data\[5\] net73 VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1405_ _0734_ _0735_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__and3b_1
X_1336_ _0689_ _0617_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__and3b_1
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 reg_dat_di[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_1267_ _0639_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
X_1198_ net91 _0301_ _0302_ net90 _0544_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1543__A _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1121_ _0511_ _0508_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1052_ send_divcnt\[18\] VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_124_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1581__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0905_ _0303_ _0311_ _0307_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__or3b_1
XFILLER_0_114_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0836_ recv_divcnt\[8\] VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1363__A _0700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1319_ send_divcnt\[23\] _0674_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_142_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_886 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1392__C1 _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1670_ clknet_4_12_0_clk _0122_ VGND VGND VPWR VPWR recv_divcnt\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output96_A net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1104_ send_pattern\[3\] _0493_ _0495_ net2 _0500_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1035_ _0409_ _0410_ _0419_ _0433_ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0819_ _0237_ _0242_ _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1184__A_N net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1434__C _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1653_ clknet_4_2_0_clk _0105_ VGND VGND VPWR VPWR recv_divcnt\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0810__A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1584_ clknet_4_14_0_clk _0036_ VGND VGND VPWR VPWR send_bitcnt\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1108__C1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0956__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1018_ _0414_ _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_864 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1347__C1 _0514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1254__C _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1114__A2 _0493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0873__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0873__B2 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1050__A1 _0319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_536 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1636_ clknet_4_15_0_clk _0088_ VGND VGND VPWR VPWR recv_buf_data\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1567_ clknet_4_13_0_clk _0019_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_786 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1498_ recv_divcnt\[25\] _0165_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1665__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1032__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1546__A _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1421_ recv_divcnt\[6\] _0745_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__or2_1
X_1352_ _0701_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__clkbuf_4
X_1283_ send_divcnt\[14\] _0648_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0837__A1 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0837__B2 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0998_ _0399_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1366__A _0700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1014__B2 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1014__A1 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1619_ clknet_4_10_0_clk _0071_ VGND VGND VPWR VPWR send_divcnt\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1442__C _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0921_ _0228_ _0325_ _0339_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_16_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0852_ recv_divcnt\[11\] VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0783_ _0211_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1404_ _0341_ _0732_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__nand2_1
X_1335_ send_divcnt\[27\] _0686_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__or2_1
Xinput2 reg_dat_di[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_1266_ _0514_ _0637_ _0638_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1197_ _0575_ _0580_ _0582_ _0571_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__o22a_1
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1262__C _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1120_ send_bitcnt\[0\] VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1051_ send_divcnt\[19\] VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0904_ recv_divcnt\[18\] VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0813__A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0835_ recv_divcnt\[9\] VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0959__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1318_ send_divcnt\[23\] send_divcnt\[22\] send_divcnt\[21\] _0668_ VGND VGND VPWR
+ VPWR _0677_ sky130_fd_sc_hd__and4_1
XFILLER_0_47_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1249_ _0421_ _0622_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1208__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output89_A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1135__B1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1103_ send_pattern\[1\] _0496_ _0501_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_37_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1034_ _0417_ _0414_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_37_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_8_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0818_ _0232_ recv_divcnt\[4\] recv_divcnt\[3\] _0235_ VGND VGND VPWR VPWR _0243_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__1374__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1571__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1450__C _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1652_ clknet_4_2_0_clk _0104_ VGND VGND VPWR VPWR recv_divcnt\[13\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1583_ clknet_4_11_0_clk _0035_ VGND VGND VPWR VPWR send_bitcnt\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0972__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1017_ _0415_ send_divcnt\[9\] _0409_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1369__A _0700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_504 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1594__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_640 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1174__A_N net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0821__A net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1635_ clknet_4_15_0_clk _0087_ VGND VGND VPWR VPWR recv_buf_data\[4\] sky130_fd_sc_hd__dfxtp_1
X_1566_ clknet_4_13_0_clk _0018_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1497_ recv_divcnt\[25\] recv_divcnt\[24\] recv_divcnt\[23\] _0159_ VGND VGND VPWR
+ VPWR _0168_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1420_ recv_divcnt\[6\] recv_divcnt\[5\] recv_divcnt\[4\] _0738_ VGND VGND VPWR VPWR
+ _0748_ sky130_fd_sc_hd__and4_1
XFILLER_0_121_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1351_ _0346_ _0606_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__or2_1
X_1282_ _0650_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_69_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0997_ _0381_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1618_ clknet_4_10_0_clk _0070_ VGND VGND VPWR VPWR send_divcnt\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1632__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1549_ clknet_4_5_0_clk _0001_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_69_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ _0344_ _0275_ _0324_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__nor3_1
XFILLER_0_126_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0851_ _0230_ _0251_ _0252_ _0275_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0782_ recv_buf_data\[4\] net73 VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1655__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1403_ _0728_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1334_ send_divcnt\[27\] _0686_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__and2_1
X_1265_ send_divcnt\[9\] _0634_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__or2_1
Xinput3 reg_dat_di[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_1196_ _0581_ _0574_ _0573_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_807 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1678__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1162__A1 _0319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ _0319_ send_divcnt\[21\] _0448_ _0449_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0903_ recv_divcnt\[23\] VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0834_ _0257_ recv_divcnt\[13\] recv_divcnt\[12\] _0258_ VGND VGND VPWR VPWR _0259_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_782 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0975__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1317_ _0676_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1248_ _0421_ _0622_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1179_ _0258_ recv_divcnt\[11\] recv_divcnt\[10\] _0270_ VGND VGND VPWR VPWR _0565_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_137_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1273__C _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1102_ send_pattern\[2\] _0493_ _0495_ net1 _0500_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1033_ net111 _0412_ _0420_ _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0817_ _0236_ recv_divcnt\[2\] _0240_ _0241_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_663 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1651_ clknet_4_3_0_clk _0103_ VGND VGND VPWR VPWR recv_divcnt\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1582_ clknet_4_11_0_clk _0034_ VGND VGND VPWR VPWR send_bitcnt\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1016_ net83 _0408_ _0410_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_139_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_12_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1634_ clknet_4_15_0_clk _0086_ VGND VGND VPWR VPWR recv_buf_data\[3\] sky130_fd_sc_hd__dfxtp_1
X_1565_ clknet_4_13_0_clk _0017_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1496_ _0167_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_147_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1281__C _0616_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0922__A _0346_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_836 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1350_ net47 VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__clkbuf_4
X_1281_ _0648_ _0649_ _0616_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__and3b_1
XFILLER_0_92_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1584__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0832__A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0996_ net105 net34 net46 VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1617_ clknet_4_8_0_clk _0069_ VGND VGND VPWR VPWR send_divcnt\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__0978__S net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1548_ clknet_4_15_0_clk _0000_ VGND VGND VPWR VPWR recv_buf_valid sky130_fd_sc_hd__dfxtp_1
X_1479_ _0729_ _0153_ _0154_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output102_A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1467__B _0735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0850_ _0263_ _0267_ _0272_ _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0781_ _0210_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_474 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1507__A_N _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1483__A _0729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1402_ _0341_ _0732_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__nor2_1
X_1333_ _0688_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
X_1264_ send_divcnt\[9\] _0634_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__nand2_1
Xinput4 reg_dat_di[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0827__A net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1195_ _0569_ _0570_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_703 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_0_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0979_ _0381_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1156__C1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1622__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0902_ _0293_ _0298_ _0326_ _0291_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0833_ net85 VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1386__C1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_102_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1316_ _0674_ _0675_ _0616_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__and3b_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1247_ _0624_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1178_ recv_divcnt\[7\] net112 VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__or2b_1
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_706 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_780 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1645__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1101_ send_pattern\[1\] _0493_ _0496_ net114 _0500_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1032_ net109 _0421_ _0428_ _0430_ _0431_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_37_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1071__B2 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput40 reg_div_di[7] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0816_ _0238_ recv_divcnt\[1\] VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_92_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1668__CLK clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_675 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0925__A _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0800__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1650_ clknet_4_0_0_clk _0102_ VGND VGND VPWR VPWR recv_divcnt\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1581_ clknet_4_15_0_clk _0033_ VGND VGND VPWR VPWR send_pattern\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output94_A net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1108__A2 _0493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1491__A _0729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ net113 VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0849__B2 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1633_ clknet_4_15_0_clk _0085_ VGND VGND VPWR VPWR recv_buf_data\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1564_ clknet_4_13_0_clk _0016_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_2
X_1495_ _0165_ _0166_ _0728_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__and3b_1
XFILLER_0_146_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_612 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_778 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1280_ send_divcnt\[13\] _0645_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ _0397_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1616_ clknet_4_9_0_clk _0068_ VGND VGND VPWR VPWR send_divcnt\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1547_ _0203_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
X_1478_ recv_divcnt\[20\] _0150_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_807 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0780_ recv_buf_data\[3\] net73 VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1401_ _0733_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
X_1332_ _0686_ _0687_ _0616_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__and3b_1
XANTENNA__1551__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1263_ _0636_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 reg_dat_di[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1194_ _0565_ _0566_ _0568_ _0577_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0843__A net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1377__C _0347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0978_ net98 net27 net46 VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_751 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1574__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1478__B _0150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0901_ _0289_ _0287_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__or2b_1
XFILLER_0_56_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0832_ net86 VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1138__B1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1315_ send_divcnt\[21\] _0668_ send_divcnt\[22\] VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_108_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1246_ _0514_ _0622_ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1177_ _0229_ recv_divcnt\[6\] _0560_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_72_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1100_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1031_ _0246_ send_divcnt\[6\] VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_662 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 reg_div_di[27] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput41 reg_div_di[8] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
X_0815_ _0238_ recv_divcnt\[1\] recv_divcnt\[0\] _0239_ VGND VGND VPWR VPWR _0240_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_92_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1229_ send_divcnt\[1\] send_divcnt\[0\] VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1612__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1580_ clknet_4_15_0_clk _0032_ VGND VGND VPWR VPWR send_pattern\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1475__C _0728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output87_A net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ net113 _0413_ _0411_ net112 VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_610 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_665 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1385__C _0347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1682__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1635__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_778 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1701_ net73 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1658__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1632_ clknet_4_15_0_clk _0084_ VGND VGND VPWR VPWR recv_buf_data\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1563_ clknet_4_13_0_clk _0015_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1494_ _0297_ _0163_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1396__B _0729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_79_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_782 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0994_ _0381_ _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1615_ clknet_4_8_0_clk _0067_ VGND VGND VPWR VPWR send_divcnt\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1546_ _0349_ _0202_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__and2_1
X_1477_ recv_divcnt\[20\] _0150_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_690 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1400_ _0729_ _0731_ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__and3_1
X_1331_ send_divcnt\[26\] _0683_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__or2_1
X_1262_ _0634_ _0635_ _0617_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__and3b_1
XFILLER_0_36_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput6 reg_dat_di[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1193_ _0562_ _0563_ _0564_ _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1020__A _0246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0977_ _0385_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1156__A1 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1690__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1529_ _0191_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_126_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0900_ _0276_ _0281_ _0282_ _0324_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a31o_1
XFILLER_0_113_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0831_ _0253_ recv_divcnt\[15\] _0255_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1314_ send_divcnt\[22\] send_divcnt\[21\] _0668_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_108_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1245_ send_divcnt\[4\] _0619_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_16_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1015__A net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1176_ _0557_ _0558_ _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1685__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_43_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1030_ net109 _0421_ _0429_ net108 VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0814_ net82 VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__inv_2
Xinput20 reg_div_di[18] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 reg_div_di[28] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput42 reg_div_di[9] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1228_ send_divcnt\[0\] _0509_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1564__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1159_ net94 _0305_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_590 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_60_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1587__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1013_ send_divcnt\[9\] VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_622 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_136_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_674 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1167__A_N net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1700_ net73 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1631_ clknet_4_14_0_clk _0083_ VGND VGND VPWR VPWR recv_buf_data\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1562_ clknet_4_7_0_clk _0014_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1493_ _0297_ _0163_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1602__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1693__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0772__A _0206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1110__C1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1542__S net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1625__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1101__C1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0993_ net103 net32 net46 VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_644 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1614_ clknet_4_8_0_clk _0066_ VGND VGND VPWR VPWR send_divcnt\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1545_ net111 net40 net43 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1476_ _0152_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1688__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1362__S _0702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1330_ send_divcnt\[26\] send_divcnt\[25\] send_divcnt\[24\] _0677_ VGND VGND VPWR
+ VPWR _0686_ sky130_fd_sc_hd__and4_1
X_1261_ _0411_ _0631_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 reg_dat_di[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1192_ _0568_ _0575_ _0576_ _0577_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__or4b_1
XFILLER_0_36_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_599 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0976_ _0381_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1528_ _0700_ _0190_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__and2_1
X_1459_ _0139_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_126_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1092__A1 _0465_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output100_A net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0830_ net87 _0254_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1138__A2 _0524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1313_ _0673_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__0897__B2 _0319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0897__A1 _0313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1244_ send_divcnt\[4\] _0619_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1175_ net111 _0247_ _0559_ _0560_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__a211o_1
XFILLER_0_149_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1031__A _0246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0959_ net91 net20 net45 VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_803 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1056__A1 _0320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput10 reg_dat_we VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0813_ net93 VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__inv_2
Xinput21 reg_div_di[19] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput43 reg_div_we[0] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput32 reg_div_di[29] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1227_ _0609_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__0865__A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1158_ net92 recv_divcnt\[18\] VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1089_ net105 _0477_ _0474_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_101_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1696__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1210__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1545__S net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1012_ send_divcnt\[7\] VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1365__S _0702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1630_ clknet_4_11_0_clk _0082_ VGND VGND VPWR VPWR recv_pattern\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output92_A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1561_ clknet_4_7_0_clk _0013_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_50_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1492_ _0164_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1577__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0992_ _0395_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1613_ clknet_4_8_0_clk _0065_ VGND VGND VPWR VPWR send_divcnt\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1544_ _0201_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1475_ _0150_ _0151_ _0728_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__and3b_1
XFILLER_0_10_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1260_ _0411_ _0631_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__nor2_1
Xinput8 reg_dat_di[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_1191_ _0268_ recv_divcnt\[9\] recv_divcnt\[8\] _0415_ VGND VGND VPWR VPWR _0577_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0975_ net97 net26 net45 VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1527_ net93 net22 net43 VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__mux2_1
X_1458_ _0137_ _0138_ _0740_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_126_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_143_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1389_ recv_pattern\[6\] _0219_ _0347_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__or3_1
XANTENNA__1699__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1615__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1312_ _0514_ _0671_ _0672_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1243_ _0621_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1174_ net112 recv_divcnt\[7\] VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1312__A _0514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0958_ _0372_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1638__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0889_ _0313_ recv_divcnt\[23\] VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_835 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1368__S _0702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__B net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1525__B1 _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0971__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_615 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput11 reg_div_di[0] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
Xinput22 reg_div_di[1] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
X_0812_ _0235_ recv_divcnt\[3\] recv_divcnt\[2\] _0236_ VGND VGND VPWR VPWR _0237_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput44 reg_div_we[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput33 reg_div_di[2] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1226_ _0349_ _0607_ _0608_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1157_ net91 _0301_ _0302_ net90 VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1088_ _0484_ _0476_ _0487_ _0470_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__o31a_1
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1127__A _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1011_ send_divcnt\[8\] VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1209_ _0592_ _0593_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_0_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_830 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1560_ clknet_4_7_0_clk _0012_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfxtp_4
XANTENNA_output85_A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1491_ _0729_ _0162_ _0163_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1689_ net73 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1101__B2 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ _0381_ _0394_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_57_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1612_ clknet_4_8_0_clk _0064_ VGND VGND VPWR VPWR send_divcnt\[21\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1671__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1543_ _0349_ _0200_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1474_ recv_divcnt\[19\] _0147_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0906__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1190_ net113 _0261_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__nor2_1
Xinput9 reg_dat_re VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0974_ _0383_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1526_ net43 net11 _0189_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1045__A _0320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1457_ recv_divcnt\[15\] _0134_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_143_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1388_ recv_buf_data\[5\] _0348_ _0724_ _0350_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_143_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1567__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0778__B net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1311_ send_divcnt\[21\] _0668_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1242_ _0619_ _0620_ _0617_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1173_ _0229_ recv_divcnt\[6\] recv_divcnt\[5\] _0246_ VGND VGND VPWR VPWR _0559_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_755 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0957_ _0360_ _0371_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0888_ net97 VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__clkinv_2
Xoutput110 net110 VGND VGND VPWR VPWR reg_div_do[6] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1509_ recv_divcnt\[28\] _0174_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1165__B_N net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1503__A _0729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1525__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0811_ net104 VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput12 reg_div_di[10] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_30_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput45 reg_div_we[2] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput23 reg_div_di[20] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 reg_div_di[30] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1225_ _0216_ _0604_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1156_ net94 _0305_ _0329_ net92 VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_36_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1087_ _0475_ _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1605__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ net84 send_divcnt\[11\] VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__or2b_1
XANTENNA__1628__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_699 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1208_ net103 _0226_ _0592_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__o211a_1
XANTENNA__1053__A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1139_ recv_state\[3\] recv_state\[2\] recv_state\[1\] VGND VGND VPWR VPWR _0525_
+ sky130_fd_sc_hd__or3_2
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0786__B net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_842 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1490_ recv_divcnt\[23\] _0159_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1304__C _0616_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1104__C1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1048__A _0313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1688_ net73 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_588 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1511__A _0735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1110__A2 _0493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0797__A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1180__A_N net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1405__B _0735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1101__A2 _0493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0990_ net102 net31 net46 VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1611_ clknet_4_8_0_clk _0063_ VGND VGND VPWR VPWR send_divcnt\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1542_ net110 net39 net43 VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1473_ recv_divcnt\[19\] recv_divcnt\[18\] _0137_ _0143_ VGND VGND VPWR VPWR _0150_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_614 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0842__B2 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0842__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1151__A _0315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0973_ _0381_ _0382_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1525_ net43 _0239_ _0351_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1456_ recv_divcnt\[15\] recv_divcnt\[14\] recv_divcnt\[13\] _0766_ VGND VGND VPWR
+ VPWR _0137_ sky130_fd_sc_hd__and4_1
X_1387_ recv_pattern\[5\] _0219_ _0347_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_143_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0884__B net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0824__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1661__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_550 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_723 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_94_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1146__A _0313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1310_ send_divcnt\[21\] _0668_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__nand2_1
X_1241_ send_divcnt\[3\] _0614_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ _0246_ recv_divcnt\[5\] recv_divcnt\[4\] _0231_ VGND VGND VPWR VPWR _0558_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_125_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0956_ net90 net19 net45 VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput100 net100 VGND VGND VPWR VPWR reg_div_do[26] sky130_fd_sc_hd__clkbuf_1
X_0887_ recv_divcnt\[22\] VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0990__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput111 net111 VGND VGND VPWR VPWR reg_div_do[7] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1508_ _0176_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0895__A net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1439_ _0762_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0981__A0 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0810_ net107 VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__inv_2
Xinput13 reg_div_di[11] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput46 reg_div_we[3] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_4
XFILLER_0_24_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput24 reg_div_di[21] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput35 reg_div_di[31] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0972__A0 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1224_ _0599_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1155_ _0320_ recv_divcnt\[19\] VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1086_ _0286_ send_divcnt\[26\] _0467_ _0485_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_36_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0939_ _0359_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1207_ _0335_ recv_divcnt\[29\] VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1138_ _0498_ _0524_ _0350_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1069_ send_divcnt\[29\] VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1228__B _0509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1178__B_N net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1410__C _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1320__C _0616_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1687_ net73 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_784 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1475__A_N _0150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output109_A net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1270__C1 _0509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1610_ clknet_4_2_0_clk _0062_ VGND VGND VPWR VPWR send_divcnt\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output90_A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1541_ _0199_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1472_ _0149_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_105_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_148_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_123_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_132_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_141_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0972_ net96 net25 net45 VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1524_ _0188_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1455_ _0136_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
X_1386_ recv_buf_data\[4\] _0348_ _0723_ _0350_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_143_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1240_ send_divcnt\[3\] send_divcnt\[2\] send_divcnt\[1\] send_divcnt\[0\] VGND VGND
+ VPWR VPWR _0619_ sky130_fd_sc_hd__and4_1
XFILLER_0_47_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1171_ _0554_ _0555_ _0556_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_125_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_805 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0955_ _0370_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0886_ _0309_ _0310_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput101 net101 VGND VGND VPWR VPWR reg_div_do[27] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput112 net112 VGND VGND VPWR VPWR reg_div_do[8] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1507_ _0174_ _0735_ _0175_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__and3b_1
XFILLER_0_49_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1438_ _0729_ _0760_ _0761_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__and3_1
X_1369_ _0700_ _0713_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput36 reg_div_di[3] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput14 reg_div_di[12] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 reg_div_di[22] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput47 resetn VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1223_ _0218_ _0525_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1154_ net98 _0328_ _0535_ _0538_ _0539_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1085_ _0286_ send_divcnt\[26\] send_divcnt\[25\] _0290_ _0484_ VGND VGND VPWR VPWR
+ _0485_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0938_ _0351_ _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_151_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0869_ net98 VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1651__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1198__B2 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1198__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1674__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_587 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1206_ _0335_ recv_divcnt\[29\] recv_divcnt\[28\] _0473_ VGND VGND VPWR VPWR _0592_
+ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_4_7_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1137_ net45 _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__nor2_2
XFILLER_0_149_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1350__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1068_ send_divcnt\[26\] VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1509__B _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_142_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0918__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1686_ net73 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0909__A1 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1540_ _0349_ _0198_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output83_A net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1471_ _0147_ _0735_ _0148_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__and3b_1
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1669_ clknet_4_12_0_clk _0121_ VGND VGND VPWR VPWR recv_divcnt\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1004__B1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_15_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0971_ net47 VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1523_ _0735_ _0186_ _0187_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1454_ _0134_ _0135_ _0740_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__and3b_1
X_1385_ recv_pattern\[4\] _0219_ _0347_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_143_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1608__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_582 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ _0231_ recv_divcnt\[4\] recv_divcnt\[3\] _0232_ VGND VGND VPWR VPWR _0556_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_125_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0954_ _0360_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0885_ net91 recv_divcnt\[18\] VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput102 net102 VGND VGND VPWR VPWR reg_div_do[28] sky130_fd_sc_hd__clkbuf_1
Xoutput113 net113 VGND VGND VPWR VPWR reg_div_do[9] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1506_ recv_divcnt\[26\] _0168_ recv_divcnt\[27\] VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1437_ recv_divcnt\[10\] _0757_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__or2_1
X_1368_ recv_pattern\[6\] recv_pattern\[5\] _0702_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1299_ send_divcnt\[18\] _0661_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_39_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1580__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1528__A _0700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_699 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput37 reg_div_di[4] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput15 reg_div_di[13] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 reg_div_di[23] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput48 ser_rx VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1438__A _0729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1382__C1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1222_ _0604_ _0605_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__nor2_1
X_1153_ _0294_ recv_divcnt\[23\] _0533_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__a21oi_1
X_1084_ _0288_ send_divcnt\[27\] VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_606 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0937_ net84 net13 net44 VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_3_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0868_ _0287_ _0289_ _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__or3b_1
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0799_ _0222_ recv_divcnt\[31\] VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1258__A _0514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1183__A_N net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_599 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1205_ _0531_ _0587_ _0589_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1136_ net43 send_dummy net46 net44 VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1067_ _0290_ send_divcnt\[25\] send_divcnt\[24\] _0294_ VGND VGND VPWR VPWR _0467_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__0881__B2 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0881__A1 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1104__A2 _0493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1685_ net73 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1119_ send_pattern\[8\] _0509_ _0510_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__o21a_1
XANTENNA__0854__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1664__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_11_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1470_ recv_divcnt\[18\] _0144_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1089__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1668_ clknet_4_9_0_clk _0120_ VGND VGND VPWR VPWR recv_divcnt\[29\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1599_ clknet_4_0_0_clk _0051_ VGND VGND VPWR VPWR send_divcnt\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1266__A _0514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output114_A net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0970_ _0380_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1522_ recv_divcnt\[31\] _0183_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1453_ recv_divcnt\[14\] _0131_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__or2_1
X_1384_ recv_buf_data\[3\] _0348_ _0722_ _0350_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_143_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0993__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0984__A0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_72_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0953_ net89 net18 net45 VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0975__A0 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0884_ recv_divcnt\[19\] net92 VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput103 net103 VGND VGND VPWR VPWR reg_div_do[29] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput114 net114 VGND VGND VPWR VPWR ser_tx sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1505_ recv_divcnt\[27\] recv_divcnt\[26\] _0168_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1436_ recv_divcnt\[10\] _0757_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__nand2_1
X_1367_ _0712_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1298_ send_divcnt\[18\] _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_90_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_129_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput16 reg_div_di[14] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput27 reg_div_di[24] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput38 reg_div_di[5] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1221_ recv_state\[2\] _0603_ _0351_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__o21ai_1
X_1152_ net95 _0304_ _0536_ _0537_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__a31o_1
X_1083_ send_divcnt\[31\] VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0936_ _0357_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0867_ _0286_ recv_divcnt\[26\] recv_divcnt\[25\] _0290_ _0291_ VGND VGND VPWR VPWR
+ _0292_ sky130_fd_sc_hd__o221a_1
XFILLER_0_24_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0798_ _0222_ recv_divcnt\[31\] VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1419_ _0747_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1570__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1204_ _0529_ _0528_ _0531_ _0588_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__a2bb2o_1
X_1135_ _0521_ _0522_ _0350_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_784 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1066_ send_divcnt\[25\] VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__inv_2
XANTENNA__0962__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0919_ _0233_ _0340_ _0250_ _0343_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__or4_1
XFILLER_0_141_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1593__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1684_ net73 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0811__A net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1023__A_N net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1118_ _0500_ net8 _0495_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1049_ _0315_ send_divcnt\[22\] send_divcnt\[21\] _0319_ VGND VGND VPWR VPWR _0449_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_48_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1462__A _0729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0806__A net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1667_ clknet_4_12_0_clk _0119_ VGND VGND VPWR VPWR recv_divcnt\[28\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1598_ clknet_4_1_0_clk _0050_ VGND VGND VPWR VPWR send_divcnt\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1372__A _0700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1631__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output107_A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1521_ recv_divcnt\[31\] _0183_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1452_ recv_divcnt\[14\] recv_divcnt\[13\] _0766_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__and3_1
X_1383_ recv_pattern\[3\] _0219_ _0347_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_143_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1131__S _0493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_587 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1517__D _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1654__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1161__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_532 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0952_ _0368_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0883_ _0300_ recv_divcnt\[16\] _0303_ _0306_ _0307_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1677__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput104 net104 VGND VGND VPWR VPWR reg_div_do[2] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1504_ _0173_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1435_ _0759_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1366_ _0700_ _0711_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__and2_1
XANTENNA__1152__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0965__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1297_ _0443_ _0657_ _0661_ _0509_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_148_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1097__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput17 reg_div_di[15] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 reg_div_di[25] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput39 reg_div_di[6] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1220_ recv_state\[2\] recv_state\[1\] recv_state\[0\] _0527_ VGND VGND VPWR VPWR
+ _0604_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1151_ _0315_ recv_divcnt\[21\] VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1082_ net99 _0466_ _0467_ _0472_ _0481_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_36_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0814__A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0935_ _0351_ _0356_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1070__B1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0866_ _0288_ recv_divcnt\[27\] VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0797_ net106 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_58_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1418_ _0745_ _0746_ _0740_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__and3b_1
XFILLER_0_47_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1349_ _0483_ _0698_ _0699_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output99_A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1203_ _0290_ recv_divcnt\[24\] _0588_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_53_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1134_ _0204_ _0496_ send_bitcnt\[3\] VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_0_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1065_ _0402_ _0442_ _0459_ _0464_ _0448_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__a32o_2
XFILLER_0_88_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_721 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0918_ net104 _0341_ _0342_ _0237_ _0245_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_141_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1375__A _0700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0849_ _0270_ recv_divcnt\[11\] _0261_ net112 _0273_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_73_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1285__A _0514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1683_ net73 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_146_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1117_ _0497_ _0508_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__or2_4
XFILLER_0_88_560 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1048_ _0313_ send_divcnt\[23\] VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_700 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1446__C _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_747 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_663 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1666_ clknet_4_9_0_clk _0118_ VGND VGND VPWR VPWR recv_divcnt\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0968__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1597_ clknet_4_1_0_clk _0049_ VGND VGND VPWR VPWR send_divcnt\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1583__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1520_ _0185_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1451_ _0133_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
X_1382_ recv_buf_data\[2\] _0348_ _0721_ _0350_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_143_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_780 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1649_ clknet_4_1_0_clk _0101_ VGND VGND VPWR VPWR recv_divcnt\[10\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_886 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1394__C1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1293__A _0514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0951_ _0360_ _0367_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_45_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0882_ net90 _0301_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput105 net105 VGND VGND VPWR VPWR reg_div_do[30] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_858 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1503_ _0729_ _0171_ _0172_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__and3_1
X_1434_ _0757_ _0758_ _0740_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__and3b_1
XFILLER_0_128_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1365_ recv_pattern\[5\] recv_pattern\[4\] _0702_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1296_ send_divcnt\[15\] send_divcnt\[14\] _0648_ _0660_ VGND VGND VPWR VPWR _0661_
+ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_39_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0981__S net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput18 reg_div_di[16] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput29 reg_div_di[26] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1454__C _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1150_ _0315_ recv_divcnt\[21\] VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1081_ net100 _0468_ _0474_ _0480_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a211oi_1
XANTENNA__0893__A1 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1644__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0934_ net83 net12 net44 VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0865_ net99 VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0830__A net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0796_ net105 recv_divcnt\[30\] VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_58_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_580 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1417_ recv_divcnt\[4\] _0738_ recv_divcnt\[5\] VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1348_ _0483_ _0698_ _0500_ _0495_ _0493_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__a2111oi_1
X_1279_ send_divcnt\[13\] send_divcnt\[12\] send_divcnt\[11\] _0641_ VGND VGND VPWR
+ VPWR _0648_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_864 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_672 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1667__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_730 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1202_ net100 _0296_ _0297_ net99 VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_53_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1133_ _0491_ _0508_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1064_ _0449_ _0463_ _0402_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_0_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_642 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0917_ _0229_ recv_divcnt\[7\] recv_divcnt\[0\] _0239_ _0241_ VGND VGND VPWR VPWR
+ _0342_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0848_ _0258_ recv_divcnt\[12\] VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0779_ _0209_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_723 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1682_ net73 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1116_ _0492_ _0494_ _0498_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__or3_2
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1047_ net89 send_divcnt\[16\] VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_24_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1016__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_675 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1665_ clknet_4_8_0_clk _0117_ VGND VGND VPWR VPWR recv_divcnt\[26\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1596_ clknet_4_1_0_clk _0048_ VGND VGND VPWR VPWR send_divcnt\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0984__S net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0996__A0 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0987__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1450_ _0131_ _0132_ _0740_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__and3b_1
X_1381_ recv_pattern\[2\] _0219_ _0347_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0978__A0 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0833__A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1648_ clknet_4_1_0_clk _0100_ VGND VGND VPWR VPWR recv_divcnt\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1579_ clknet_4_15_0_clk _0031_ VGND VGND VPWR VPWR send_pattern\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1550__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1277__C _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1394__B1 _0702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output112_A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0950_ net88 net17 net44 VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0881_ net94 _0304_ _0305_ net92 VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput106 net106 VGND VGND VPWR VPWR reg_div_do[31] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1573__CLK clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1502_ recv_divcnt\[26\] _0168_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1433_ recv_divcnt\[9\] _0754_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__or2_1
X_1364_ _0710_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_50_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0828__A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1295_ send_divcnt\[17\] send_divcnt\[16\] VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput19 reg_div_di[17] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_107_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1080_ _0294_ send_divcnt\[24\] _0475_ _0476_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_36_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1479__A _0729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0933_ _0355_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0864_ _0288_ recv_divcnt\[27\] VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_868 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0795_ recv_divcnt\[29\] VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1416_ recv_divcnt\[5\] recv_divcnt\[4\] _0738_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__and3_1
X_1347_ send_divcnt\[30\] _0695_ _0698_ _0514_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__o211a_1
XANTENNA__1530__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1278_ _0647_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_578 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1201_ _0540_ _0550_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_53_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1611__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1132_ _0498_ _0520_ _0350_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_0_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1063_ _0319_ send_divcnt\[21\] _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0916_ recv_divcnt\[2\] VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_835 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0847_ _0268_ recv_divcnt\[10\] _0269_ _0271_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__a211o_1
XFILLER_0_141_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0778_ recv_buf_data\[2\] net73 VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0987__S net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1634__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1681_ net73 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1115_ send_pattern\[7\] _0496_ _0507_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1046_ _0444_ _0445_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_24_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1657__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1664_ clknet_4_8_0_clk _0116_ VGND VGND VPWR VPWR recv_divcnt\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1595_ clknet_4_4_0_clk _0047_ VGND VGND VPWR VPWR send_divcnt\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1029_ send_divcnt\[4\] VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1173__B2 _0246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0923__B _0347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1380_ recv_buf_data\[1\] _0348_ _0720_ _0350_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1010__A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1647_ clknet_4_4_0_clk _0099_ VGND VGND VPWR VPWR recv_divcnt\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__1383__C _0347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1578_ clknet_4_13_0_clk _0030_ VGND VGND VPWR VPWR send_pattern\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1680__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output105_A net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ recv_divcnt\[19\] VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput107 net107 VGND VGND VPWR VPWR reg_div_do[3] sky130_fd_sc_hd__clkbuf_1
X_1501_ recv_divcnt\[26\] _0168_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1432_ recv_divcnt\[9\] recv_divcnt\[8\] recv_divcnt\[7\] _0748_ VGND VGND VPWR VPWR
+ _0757_ sky130_fd_sc_hd__and4_1
X_1363_ _0700_ _0709_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1294_ _0659_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_19_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0929__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_814 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0932_ _0351_ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0863_ net101 VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_151_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0794_ _0218_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1415_ _0744_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1346_ _0477_ _0469_ _0692_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_71_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1277_ _0645_ _0646_ _0617_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__and3b_1
XFILLER_0_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1563__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1200_ _0579_ _0583_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_148_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1131_ send_bitcnt\[2\] _0519_ _0493_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1062_ _0460_ _0457_ _0461_ _0456_ _0445_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0915_ _0240_ _0243_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0846_ _0270_ recv_divcnt\[11\] VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__nor2_1
X_0777_ _0208_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1391__C _0347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_126_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1329_ _0685_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__1586__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_144_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_622 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1680_ net73 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output97_A net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1166__A_N net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1114_ send_pattern\[8\] _0493_ _0495_ net7 _0500_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__a221o_1
X_1045_ _0320_ send_divcnt\[20\] VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_24_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0829_ recv_divcnt\[14\] VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__inv_2
XANTENNA__1683__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1601__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_152_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1487__B _0735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1663_ clknet_4_9_0_clk _0115_ VGND VGND VPWR VPWR recv_divcnt\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1594_ clknet_4_4_0_clk _0046_ VGND VGND VPWR VPWR send_divcnt\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1028_ _0425_ _0426_ _0427_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1624__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_728 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1527__S net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1647__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1388__C1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_496 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1646_ clknet_4_4_0_clk _0098_ VGND VGND VPWR VPWR recv_divcnt\[7\] sky130_fd_sc_hd__dfxtp_2
X_1577_ clknet_4_13_0_clk _0029_ VGND VGND VPWR VPWR send_pattern\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_728 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1082__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_806 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1500_ _0170_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput108 net108 VGND VGND VPWR VPWR reg_div_do[4] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1431_ _0756_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1362_ recv_pattern\[4\] recv_pattern\[3\] _0702_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__mux2_1
Xoutput90 net90 VGND VGND VPWR VPWR reg_div_do[17] sky130_fd_sc_hd__clkbuf_1
X_1293_ _0514_ _0657_ _0658_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1629_ clknet_4_11_0_clk _0081_ VGND VGND VPWR VPWR recv_pattern\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1691__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_812 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0770__A send_dummy VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1119__A2 _0509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0878__B2 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0878__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_672 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0931_ net113 net42 net44 VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0802__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0802__B2 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0862_ _0286_ recv_divcnt\[26\] VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__and2_1
X_0793_ _0216_ recv_state\[2\] _0217_ recv_state\[0\] VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1414_ _0729_ _0742_ _0743_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1345_ _0697_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1276_ send_divcnt\[12\] _0642_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1389__C _0347_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1686__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1037__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1037__B2 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_777 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1130_ _0204_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_53_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1061_ _0455_ send_divcnt\[19\] send_divcnt\[18\] _0453_ VGND VGND VPWR VPWR _0461_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0914_ _0285_ _0327_ _0334_ _0299_ _0338_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__o221a_1
XFILLER_0_50_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0845_ net84 VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0776_ recv_buf_data\[1\] net73 VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1328_ _0683_ _0684_ _0616_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__and3b_1
X_1259_ _0633_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1019__A1 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1019__B2 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0950__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_634 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0941__A0 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1113_ send_pattern\[6\] _0496_ _0506_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1044_ net90 _0443_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_870 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0828_ net88 VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0999__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1576__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1662_ clknet_4_3_0_clk _0114_ VGND VGND VPWR VPWR recv_divcnt\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1593_ clknet_4_4_0_clk _0045_ VGND VGND VPWR VPWR send_divcnt\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0863__A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1027_ _0232_ send_divcnt\[4\] send_divcnt\[3\] _0235_ VGND VGND VPWR VPWR _0427_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_81_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1694__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1599__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1024__B_N net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_615 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1645_ clknet_4_4_0_clk _0097_ VGND VGND VPWR VPWR recv_divcnt\[6\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_20_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1576_ clknet_4_13_0_clk _0028_ VGND VGND VPWR VPWR send_pattern\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__0858__A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1689__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_818 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput109 net109 VGND VGND VPWR VPWR reg_div_do[5] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1430_ _0754_ _0755_ _0740_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__and3b_1
XFILLER_0_121_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1361_ _0708_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__1614__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput80 net80 VGND VGND VPWR VPWR reg_dat_do[9] sky130_fd_sc_hd__clkbuf_1
Xoutput91 net91 VGND VGND VPWR VPWR reg_div_do[18] sky130_fd_sc_hd__clkbuf_1
XANTENNA__1542__A0 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1292_ send_divcnt\[16\] _0654_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_19_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1628_ clknet_4_14_0_clk _0080_ VGND VGND VPWR VPWR recv_pattern\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1533__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1559_ clknet_4_6_0_clk _0011_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_107_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1297__C1 _0509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_784 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1637__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output110_A net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0930_ _0353_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0861_ net100 VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0792_ recv_state\[1\] VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1495__C _0728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_637 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1413_ recv_divcnt\[4\] _0738_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1344_ _0695_ _0617_ _0696_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_71_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1275_ send_divcnt\[12\] send_divcnt\[11\] _0641_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1060_ _0300_ send_divcnt\[16\] _0444_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0913_ _0335_ _0337_ _0223_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0844_ _0268_ recv_divcnt\[10\] _0260_ net113 VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_43_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0775_ _0207_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1327_ _0466_ _0680_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__nand2_1
X_1258_ _0514_ _0631_ _0632_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_3_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1189_ _0572_ _0573_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_84_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1697__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_805 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1371__S _0702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1400__A _0729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1112_ send_pattern\[7\] _0493_ _0495_ net6 _0500_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1043_ send_divcnt\[17\] VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0827_ net110 _0247_ _0248_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_874 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_75_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1661_ clknet_4_12_0_clk _0113_ VGND VGND VPWR VPWR recv_divcnt\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1592_ clknet_4_5_0_clk _0044_ VGND VGND VPWR VPWR send_divcnt\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_93_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1026_ _0235_ send_divcnt\[3\] send_divcnt\[2\] _0236_ VGND VGND VPWR VPWR _0426_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1670__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_866 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1644_ clknet_4_4_0_clk _0096_ VGND VGND VPWR VPWR recv_divcnt\[5\] sky130_fd_sc_hd__dfxtp_2
X_1575_ clknet_4_12_0_clk _0027_ VGND VGND VPWR VPWR send_pattern\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ _0270_ send_divcnt\[11\] _0408_ net83 VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_92_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1566__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_149_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput70 net70 VGND VGND VPWR VPWR reg_dat_do[29] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1360_ _0700_ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput81 net81 VGND VGND VPWR VPWR reg_dat_wait sky130_fd_sc_hd__clkbuf_1
Xoutput92 net92 VGND VGND VPWR VPWR reg_div_do[19] sky130_fd_sc_hd__clkbuf_1
X_1291_ send_divcnt\[16\] _0654_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1627_ clknet_4_14_0_clk _0079_ VGND VGND VPWR VPWR recv_pattern\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0869__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1558_ clknet_4_7_0_clk _0010_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfxtp_4
X_1489_ recv_divcnt\[23\] _0159_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_107_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1221__B1 _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1374__S _0702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1403__A _0728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output103_A net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_699 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0860_ _0225_ _0284_ _0227_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__or3b_1
XFILLER_0_36_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0791_ recv_state\[3\] VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1412_ recv_divcnt\[4\] _0738_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1343_ send_divcnt\[29\] _0692_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_71_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1274_ _0644_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ _0393_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1604__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0912_ _0336_ _0224_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0843_ net83 VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0774_ recv_buf_data\[0\] net73 VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1326_ _0466_ _0680_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_88_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1257_ send_divcnt\[7\] _0628_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__or2_1
X_1188_ recv_divcnt\[12\] _0257_ net87 _0264_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1627__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0882__A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0776__B net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1112__C1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_122_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1111_ send_pattern\[5\] _0496_ _0505_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1042_ _0407_ _0435_ _0439_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_728 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_644 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0826_ _0234_ _0244_ _0245_ _0250_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_6_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1038__A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_886 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1309_ _0670_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1660_ clknet_4_12_0_clk _0112_ VGND VGND VPWR VPWR recv_divcnt\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output95_A net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1591_ clknet_4_5_0_clk _0043_ VGND VGND VPWR VPWR send_divcnt\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1025_ _0236_ send_divcnt\[2\] _0422_ _0423_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__o221a_1
XFILLER_0_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0809_ _0233_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_812 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1231__A _0514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1643_ clknet_4_4_0_clk _0095_ VGND VGND VPWR VPWR recv_divcnt\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1574_ clknet_4_11_0_clk _0026_ VGND VGND VPWR VPWR send_pattern\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1008_ send_divcnt\[10\] VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0890__A net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_814 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1226__A _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0784__B net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_14_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput60 net60 VGND VGND VPWR VPWR reg_dat_do[1] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput71 net71 VGND VGND VPWR VPWR reg_dat_do[2] sky130_fd_sc_hd__clkbuf_1
XANTENNA__1136__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput82 net82 VGND VGND VPWR VPWR reg_div_do[0] sky130_fd_sc_hd__clkbuf_1
Xoutput93 net93 VGND VGND VPWR VPWR reg_div_do[1] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1290_ _0656_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_19_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1058__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1660__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1058__B2 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1626_ clknet_4_14_0_clk _0078_ VGND VGND VPWR VPWR recv_pattern\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1557_ clknet_4_7_0_clk _0009_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_94_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1488_ _0161_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0885__A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1049__A1 _0315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1049__B2 _0319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_699 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0790_ net73 net9 VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1212__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1411_ _0741_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1342_ send_divcnt\[29\] _0692_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_71_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1273_ _0642_ _0643_ _0617_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__and3b_1
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0988_ _0381_ _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0962__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1609_ clknet_4_2_0_clk _0061_ VGND VGND VPWR VPWR send_divcnt\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0953__A0 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1414__A _0729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0911_ recv_divcnt\[30\] VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1579__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0842_ net87 _0254_ _0264_ net86 _0266_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0773_ recv_buf_valid VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkinv_8
XFILLER_0_113_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0944__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1325_ _0682_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__1324__A _0514_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1256_ send_divcnt\[7\] _0628_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__nand2_1
X_1187_ _0300_ recv_divcnt\[15\] _0254_ net88 VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_94_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_2_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1188__B1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_667 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1409__A _0728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0926__B1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1110_ send_pattern\[6\] _0493_ _0495_ net5 _0500_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ _0438_ _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_670 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0825_ _0246_ recv_divcnt\[6\] _0249_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1054__A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1308_ _0668_ _0669_ _0616_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__and3b_1
X_1239_ _0618_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1590_ clknet_4_10_0_clk _0042_ VGND VGND VPWR VPWR recv_state\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1617__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output88_A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1024_ send_divcnt\[1\] net93 VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__or2b_1
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0808_ _0231_ recv_divcnt\[5\] recv_divcnt\[4\] _0232_ VGND VGND VPWR VPWR _0233_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0888__A net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_10_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_2 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1642_ clknet_4_6_0_clk _0094_ VGND VGND VPWR VPWR recv_divcnt\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ clknet_4_9_0_clk _0025_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_10_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1545__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1007_ _0404_ _0406_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_122_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1536__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1527__A0 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput61 net61 VGND VGND VPWR VPWR reg_dat_do[20] sky130_fd_sc_hd__clkbuf_1
Xoutput50 net50 VGND VGND VPWR VPWR reg_dat_do[10] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput72 net72 VGND VGND VPWR VPWR reg_dat_do[30] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput94 net94 VGND VGND VPWR VPWR reg_div_do[20] sky130_fd_sc_hd__clkbuf_1
Xoutput83 net83 VGND VGND VPWR VPWR reg_div_do[10] sky130_fd_sc_hd__clkbuf_1
XANTENNA__1136__B send_dummy VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1215__C1 _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1625_ clknet_4_14_0_clk _0077_ VGND VGND VPWR VPWR recv_pattern\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_93_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1556_ clknet_4_7_0_clk _0008_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_94_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1487_ _0159_ _0735_ _0160_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_124_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1237__A _0616_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1700__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1147__A net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1410_ _0738_ _0739_ _0740_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__and3b_1
XFILLER_0_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1341_ _0694_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1272_ send_divcnt\[11\] _0641_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ net101 net30 net46 VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1608_ clknet_4_2_0_clk _0060_ VGND VGND VPWR VPWR send_divcnt\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0896__A _0320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1539_ net109 net38 net43 VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1650__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0910_ net105 VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0841_ _0265_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0772_ _0206_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1308__C _0616_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1324_ _0514_ _0680_ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1255_ _0630_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1186_ _0257_ recv_divcnt\[12\] _0569_ _0570_ _0571_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1673__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_579 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1040_ _0404_ _0406_ _0437_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_45_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_498 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0824_ net110 _0247_ _0248_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1307_ send_divcnt\[20\] _0665_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__or2_1
X_1238_ _0614_ _0615_ _0617_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__and3b_1
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1169_ _0232_ recv_divcnt\[3\] recv_divcnt\[2\] _0235_ VGND VGND VPWR VPWR _0555_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_137_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_830 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_595 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1569__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1155__A _0320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_811 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1023_ net82 send_divcnt\[0\] VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0807_ net108 VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_71_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_80_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_119_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_3 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1641_ clknet_4_6_0_clk _0093_ VGND VGND VPWR VPWR recv_divcnt\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_151_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1572_ clknet_4_13_0_clk _0024_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1316__C _0616_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1006_ net87 _0405_ _0403_ net86 VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_122_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1507__B _0735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1523__A _0735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1607__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput51 net51 VGND VGND VPWR VPWR reg_dat_do[11] sky130_fd_sc_hd__clkbuf_1
Xoutput73 net73 VGND VGND VPWR VPWR reg_dat_do[31] sky130_fd_sc_hd__clkbuf_1
Xoutput62 net62 VGND VGND VPWR VPWR reg_dat_do[21] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput84 net84 VGND VGND VPWR VPWR reg_div_do[11] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1136__C net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput95 net95 VGND VGND VPWR VPWR reg_div_do[21] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1624_ clknet_4_14_0_clk _0076_ VGND VGND VPWR VPWR recv_pattern\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_93_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1555_ clknet_4_7_0_clk _0007_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dfxtp_4
X_1486_ _0312_ _0157_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_500 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1390__C1 _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1340_ _0692_ _0617_ _0693_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__and3b_1
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1271_ send_divcnt\[11\] _0641_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ _0391_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1607_ clknet_4_2_0_clk _0059_ VGND VGND VPWR VPWR send_divcnt\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1538_ _0197_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1073__A net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1469_ recv_divcnt\[18\] _0137_ _0143_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output101_A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0840_ _0253_ recv_divcnt\[15\] VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0771_ net10 _0205_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1158__A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1323_ send_divcnt\[24\] _0677_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__or2_1
X_1254_ _0628_ _0629_ _0617_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_88_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1106__C1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1185_ net89 recv_divcnt\[15\] VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1340__B _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0969_ _0360_ _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1515__B _0735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1112__A2 _0493_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1531__A _0700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_100_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0823_ _0229_ recv_divcnt\[7\] VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1306_ send_divcnt\[20\] send_divcnt\[19\] send_divcnt\[18\] _0661_ VGND VGND VPWR
+ VPWR _0668_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1351__A _0346_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1237_ _0616_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__buf_4
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1168_ _0238_ recv_divcnt\[0\] _0551_ _0552_ _0553_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__a311o_1
XFILLER_0_35_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1099_ _0497_ _0498_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_842 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1030__B2 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1030__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0844__B2 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1022_ net93 send_divcnt\[1\] VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1663__CLK clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_806 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_812 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0806_ net109 VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1079__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_583 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1422__C _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1640_ clknet_4_6_0_clk _0092_ VGND VGND VPWR VPWR recv_divcnt\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1571_ clknet_4_13_0_clk _0023_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output93_A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1332__C _0616_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1005_ send_divcnt\[14\] VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1242__C _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput52 net52 VGND VGND VPWR VPWR reg_dat_do[12] sky130_fd_sc_hd__clkbuf_1
Xoutput63 net63 VGND VGND VPWR VPWR reg_dat_do[22] sky130_fd_sc_hd__clkbuf_1
Xoutput74 net74 VGND VGND VPWR VPWR reg_dat_do[3] sky130_fd_sc_hd__clkbuf_1
Xoutput85 net85 VGND VGND VPWR VPWR reg_div_do[12] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput96 net96 VGND VGND VPWR VPWR reg_div_do[22] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1623_ clknet_4_14_0_clk _0075_ VGND VGND VPWR VPWR recv_pattern\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_93_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1554_ clknet_4_7_0_clk _0006_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dfxtp_4
X_1485_ recv_divcnt\[22\] recv_divcnt\[21\] recv_divcnt\[20\] _0150_ VGND VGND VPWR
+ VPWR _0159_ sky130_fd_sc_hd__and4_1
.ends

