VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alphacore
  CLASS BLOCK ;
  FOREIGN alphacore ;
  ORIGIN 0.000 0.000 ;
  SIZE 486.885 BY 497.605 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 484.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 484.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 484.400 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 484.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 484.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 484.400 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 4.000 ;
    END
  END clk
  PIN cpi_insn[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 493.605 157.690 497.605 ;
    END
  END cpi_insn[0]
  PIN cpi_insn[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 493.605 176.090 497.605 ;
    END
  END cpi_insn[10]
  PIN cpi_insn[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 493.605 177.930 497.605 ;
    END
  END cpi_insn[11]
  PIN cpi_insn[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 493.605 179.770 497.605 ;
    END
  END cpi_insn[12]
  PIN cpi_insn[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 493.605 181.610 497.605 ;
    END
  END cpi_insn[13]
  PIN cpi_insn[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 493.605 183.450 497.605 ;
    END
  END cpi_insn[14]
  PIN cpi_insn[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 493.605 185.290 497.605 ;
    END
  END cpi_insn[15]
  PIN cpi_insn[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 493.605 187.130 497.605 ;
    END
  END cpi_insn[16]
  PIN cpi_insn[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 493.605 188.970 497.605 ;
    END
  END cpi_insn[17]
  PIN cpi_insn[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 493.605 190.810 497.605 ;
    END
  END cpi_insn[18]
  PIN cpi_insn[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 493.605 192.650 497.605 ;
    END
  END cpi_insn[19]
  PIN cpi_insn[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 493.605 159.530 497.605 ;
    END
  END cpi_insn[1]
  PIN cpi_insn[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 493.605 194.490 497.605 ;
    END
  END cpi_insn[20]
  PIN cpi_insn[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 493.605 196.330 497.605 ;
    END
  END cpi_insn[21]
  PIN cpi_insn[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 493.605 198.170 497.605 ;
    END
  END cpi_insn[22]
  PIN cpi_insn[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 493.605 200.010 497.605 ;
    END
  END cpi_insn[23]
  PIN cpi_insn[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 493.605 201.850 497.605 ;
    END
  END cpi_insn[24]
  PIN cpi_insn[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 493.605 203.690 497.605 ;
    END
  END cpi_insn[25]
  PIN cpi_insn[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 493.605 205.530 497.605 ;
    END
  END cpi_insn[26]
  PIN cpi_insn[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 493.605 207.370 497.605 ;
    END
  END cpi_insn[27]
  PIN cpi_insn[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 493.605 209.210 497.605 ;
    END
  END cpi_insn[28]
  PIN cpi_insn[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 493.605 211.050 497.605 ;
    END
  END cpi_insn[29]
  PIN cpi_insn[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 493.605 161.370 497.605 ;
    END
  END cpi_insn[2]
  PIN cpi_insn[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 493.605 212.890 497.605 ;
    END
  END cpi_insn[30]
  PIN cpi_insn[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 493.605 214.730 497.605 ;
    END
  END cpi_insn[31]
  PIN cpi_insn[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 493.605 163.210 497.605 ;
    END
  END cpi_insn[3]
  PIN cpi_insn[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 493.605 165.050 497.605 ;
    END
  END cpi_insn[4]
  PIN cpi_insn[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 493.605 166.890 497.605 ;
    END
  END cpi_insn[5]
  PIN cpi_insn[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 493.605 168.730 497.605 ;
    END
  END cpi_insn[6]
  PIN cpi_insn[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 493.605 170.570 497.605 ;
    END
  END cpi_insn[7]
  PIN cpi_insn[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 493.605 172.410 497.605 ;
    END
  END cpi_insn[8]
  PIN cpi_insn[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 493.605 174.250 497.605 ;
    END
  END cpi_insn[9]
  PIN cpi_rs1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 216.290 493.605 216.570 497.605 ;
    END
  END cpi_rs1[0]
  PIN cpi_rs1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 234.690 493.605 234.970 497.605 ;
    END
  END cpi_rs1[10]
  PIN cpi_rs1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 236.530 493.605 236.810 497.605 ;
    END
  END cpi_rs1[11]
  PIN cpi_rs1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 238.370 493.605 238.650 497.605 ;
    END
  END cpi_rs1[12]
  PIN cpi_rs1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 240.210 493.605 240.490 497.605 ;
    END
  END cpi_rs1[13]
  PIN cpi_rs1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 242.050 493.605 242.330 497.605 ;
    END
  END cpi_rs1[14]
  PIN cpi_rs1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 243.890 493.605 244.170 497.605 ;
    END
  END cpi_rs1[15]
  PIN cpi_rs1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 245.730 493.605 246.010 497.605 ;
    END
  END cpi_rs1[16]
  PIN cpi_rs1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 247.570 493.605 247.850 497.605 ;
    END
  END cpi_rs1[17]
  PIN cpi_rs1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 249.410 493.605 249.690 497.605 ;
    END
  END cpi_rs1[18]
  PIN cpi_rs1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 251.250 493.605 251.530 497.605 ;
    END
  END cpi_rs1[19]
  PIN cpi_rs1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 218.130 493.605 218.410 497.605 ;
    END
  END cpi_rs1[1]
  PIN cpi_rs1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 253.090 493.605 253.370 497.605 ;
    END
  END cpi_rs1[20]
  PIN cpi_rs1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 254.930 493.605 255.210 497.605 ;
    END
  END cpi_rs1[21]
  PIN cpi_rs1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 256.770 493.605 257.050 497.605 ;
    END
  END cpi_rs1[22]
  PIN cpi_rs1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 258.610 493.605 258.890 497.605 ;
    END
  END cpi_rs1[23]
  PIN cpi_rs1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 260.450 493.605 260.730 497.605 ;
    END
  END cpi_rs1[24]
  PIN cpi_rs1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 262.290 493.605 262.570 497.605 ;
    END
  END cpi_rs1[25]
  PIN cpi_rs1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 264.130 493.605 264.410 497.605 ;
    END
  END cpi_rs1[26]
  PIN cpi_rs1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 265.970 493.605 266.250 497.605 ;
    END
  END cpi_rs1[27]
  PIN cpi_rs1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 267.810 493.605 268.090 497.605 ;
    END
  END cpi_rs1[28]
  PIN cpi_rs1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 269.650 493.605 269.930 497.605 ;
    END
  END cpi_rs1[29]
  PIN cpi_rs1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 219.970 493.605 220.250 497.605 ;
    END
  END cpi_rs1[2]
  PIN cpi_rs1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 271.490 493.605 271.770 497.605 ;
    END
  END cpi_rs1[30]
  PIN cpi_rs1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 273.330 493.605 273.610 497.605 ;
    END
  END cpi_rs1[31]
  PIN cpi_rs1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 221.810 493.605 222.090 497.605 ;
    END
  END cpi_rs1[3]
  PIN cpi_rs1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 223.650 493.605 223.930 497.605 ;
    END
  END cpi_rs1[4]
  PIN cpi_rs1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 225.490 493.605 225.770 497.605 ;
    END
  END cpi_rs1[5]
  PIN cpi_rs1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 227.330 493.605 227.610 497.605 ;
    END
  END cpi_rs1[6]
  PIN cpi_rs1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 229.170 493.605 229.450 497.605 ;
    END
  END cpi_rs1[7]
  PIN cpi_rs1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 231.010 493.605 231.290 497.605 ;
    END
  END cpi_rs1[8]
  PIN cpi_rs1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 232.850 493.605 233.130 497.605 ;
    END
  END cpi_rs1[9]
  PIN cpi_rs2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 275.170 493.605 275.450 497.605 ;
    END
  END cpi_rs2[0]
  PIN cpi_rs2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 293.570 493.605 293.850 497.605 ;
    END
  END cpi_rs2[10]
  PIN cpi_rs2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 295.410 493.605 295.690 497.605 ;
    END
  END cpi_rs2[11]
  PIN cpi_rs2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 297.250 493.605 297.530 497.605 ;
    END
  END cpi_rs2[12]
  PIN cpi_rs2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 299.090 493.605 299.370 497.605 ;
    END
  END cpi_rs2[13]
  PIN cpi_rs2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 300.930 493.605 301.210 497.605 ;
    END
  END cpi_rs2[14]
  PIN cpi_rs2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 302.770 493.605 303.050 497.605 ;
    END
  END cpi_rs2[15]
  PIN cpi_rs2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 304.610 493.605 304.890 497.605 ;
    END
  END cpi_rs2[16]
  PIN cpi_rs2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 306.450 493.605 306.730 497.605 ;
    END
  END cpi_rs2[17]
  PIN cpi_rs2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 308.290 493.605 308.570 497.605 ;
    END
  END cpi_rs2[18]
  PIN cpi_rs2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 310.130 493.605 310.410 497.605 ;
    END
  END cpi_rs2[19]
  PIN cpi_rs2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 277.010 493.605 277.290 497.605 ;
    END
  END cpi_rs2[1]
  PIN cpi_rs2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 311.970 493.605 312.250 497.605 ;
    END
  END cpi_rs2[20]
  PIN cpi_rs2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 313.810 493.605 314.090 497.605 ;
    END
  END cpi_rs2[21]
  PIN cpi_rs2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 315.650 493.605 315.930 497.605 ;
    END
  END cpi_rs2[22]
  PIN cpi_rs2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 317.490 493.605 317.770 497.605 ;
    END
  END cpi_rs2[23]
  PIN cpi_rs2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 319.330 493.605 319.610 497.605 ;
    END
  END cpi_rs2[24]
  PIN cpi_rs2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 321.170 493.605 321.450 497.605 ;
    END
  END cpi_rs2[25]
  PIN cpi_rs2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 323.010 493.605 323.290 497.605 ;
    END
  END cpi_rs2[26]
  PIN cpi_rs2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 324.850 493.605 325.130 497.605 ;
    END
  END cpi_rs2[27]
  PIN cpi_rs2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 326.690 493.605 326.970 497.605 ;
    END
  END cpi_rs2[28]
  PIN cpi_rs2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 328.530 493.605 328.810 497.605 ;
    END
  END cpi_rs2[29]
  PIN cpi_rs2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 278.850 493.605 279.130 497.605 ;
    END
  END cpi_rs2[2]
  PIN cpi_rs2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 330.370 493.605 330.650 497.605 ;
    END
  END cpi_rs2[30]
  PIN cpi_rs2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 332.210 493.605 332.490 497.605 ;
    END
  END cpi_rs2[31]
  PIN cpi_rs2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 280.690 493.605 280.970 497.605 ;
    END
  END cpi_rs2[3]
  PIN cpi_rs2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 282.530 493.605 282.810 497.605 ;
    END
  END cpi_rs2[4]
  PIN cpi_rs2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 284.370 493.605 284.650 497.605 ;
    END
  END cpi_rs2[5]
  PIN cpi_rs2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 286.210 493.605 286.490 497.605 ;
    END
  END cpi_rs2[6]
  PIN cpi_rs2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 288.050 493.605 288.330 497.605 ;
    END
  END cpi_rs2[7]
  PIN cpi_rs2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 289.890 493.605 290.170 497.605 ;
    END
  END cpi_rs2[8]
  PIN cpi_rs2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 291.730 493.605 292.010 497.605 ;
    END
  END cpi_rs2[9]
  PIN cpi_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 493.605 155.850 497.605 ;
    END
  END cpi_valid
  PIN cpi_wait
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 493.605 334.330 497.605 ;
    END
  END cpi_wait
  PIN eoi[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 335.890 493.605 336.170 497.605 ;
    END
  END eoi[0]
  PIN eoi[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 354.290 493.605 354.570 497.605 ;
    END
  END eoi[10]
  PIN eoi[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 356.130 493.605 356.410 497.605 ;
    END
  END eoi[11]
  PIN eoi[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 357.970 493.605 358.250 497.605 ;
    END
  END eoi[12]
  PIN eoi[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 359.810 493.605 360.090 497.605 ;
    END
  END eoi[13]
  PIN eoi[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 361.650 493.605 361.930 497.605 ;
    END
  END eoi[14]
  PIN eoi[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 363.490 493.605 363.770 497.605 ;
    END
  END eoi[15]
  PIN eoi[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 365.330 493.605 365.610 497.605 ;
    END
  END eoi[16]
  PIN eoi[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 367.170 493.605 367.450 497.605 ;
    END
  END eoi[17]
  PIN eoi[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 369.010 493.605 369.290 497.605 ;
    END
  END eoi[18]
  PIN eoi[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 370.850 493.605 371.130 497.605 ;
    END
  END eoi[19]
  PIN eoi[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 337.730 493.605 338.010 497.605 ;
    END
  END eoi[1]
  PIN eoi[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 372.690 493.605 372.970 497.605 ;
    END
  END eoi[20]
  PIN eoi[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 374.530 493.605 374.810 497.605 ;
    END
  END eoi[21]
  PIN eoi[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 376.370 493.605 376.650 497.605 ;
    END
  END eoi[22]
  PIN eoi[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 378.210 493.605 378.490 497.605 ;
    END
  END eoi[23]
  PIN eoi[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 380.050 493.605 380.330 497.605 ;
    END
  END eoi[24]
  PIN eoi[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 381.890 493.605 382.170 497.605 ;
    END
  END eoi[25]
  PIN eoi[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 383.730 493.605 384.010 497.605 ;
    END
  END eoi[26]
  PIN eoi[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 385.570 493.605 385.850 497.605 ;
    END
  END eoi[27]
  PIN eoi[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 387.410 493.605 387.690 497.605 ;
    END
  END eoi[28]
  PIN eoi[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 389.250 493.605 389.530 497.605 ;
    END
  END eoi[29]
  PIN eoi[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 339.570 493.605 339.850 497.605 ;
    END
  END eoi[2]
  PIN eoi[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 391.090 493.605 391.370 497.605 ;
    END
  END eoi[30]
  PIN eoi[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 392.930 493.605 393.210 497.605 ;
    END
  END eoi[31]
  PIN eoi[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 341.410 493.605 341.690 497.605 ;
    END
  END eoi[3]
  PIN eoi[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 343.250 493.605 343.530 497.605 ;
    END
  END eoi[4]
  PIN eoi[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 345.090 493.605 345.370 497.605 ;
    END
  END eoi[5]
  PIN eoi[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 346.930 493.605 347.210 497.605 ;
    END
  END eoi[6]
  PIN eoi[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 348.770 493.605 349.050 497.605 ;
    END
  END eoi[7]
  PIN eoi[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 350.610 493.605 350.890 497.605 ;
    END
  END eoi[8]
  PIN eoi[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 352.450 493.605 352.730 497.605 ;
    END
  END eoi[9]
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 16.360 486.885 16.960 ;
    END
  END irq[0]
  PIN irq[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 165.960 486.885 166.560 ;
    END
  END irq[10]
  PIN irq[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 180.920 486.885 181.520 ;
    END
  END irq[11]
  PIN irq[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 195.880 486.885 196.480 ;
    END
  END irq[12]
  PIN irq[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 210.840 486.885 211.440 ;
    END
  END irq[13]
  PIN irq[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 225.800 486.885 226.400 ;
    END
  END irq[14]
  PIN irq[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 240.760 486.885 241.360 ;
    END
  END irq[15]
  PIN irq[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 255.720 486.885 256.320 ;
    END
  END irq[16]
  PIN irq[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 270.680 486.885 271.280 ;
    END
  END irq[17]
  PIN irq[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 285.640 486.885 286.240 ;
    END
  END irq[18]
  PIN irq[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 300.600 486.885 301.200 ;
    END
  END irq[19]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 31.320 486.885 31.920 ;
    END
  END irq[1]
  PIN irq[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 315.560 486.885 316.160 ;
    END
  END irq[20]
  PIN irq[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 330.520 486.885 331.120 ;
    END
  END irq[21]
  PIN irq[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 345.480 486.885 346.080 ;
    END
  END irq[22]
  PIN irq[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 360.440 486.885 361.040 ;
    END
  END irq[23]
  PIN irq[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 375.400 486.885 376.000 ;
    END
  END irq[24]
  PIN irq[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 390.360 486.885 390.960 ;
    END
  END irq[25]
  PIN irq[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 405.320 486.885 405.920 ;
    END
  END irq[26]
  PIN irq[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 482.885 420.280 486.885 420.880 ;
    END
  END irq[27]
  PIN irq[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 482.885 435.240 486.885 435.840 ;
    END
  END irq[28]
  PIN irq[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 482.885 450.200 486.885 450.800 ;
    END
  END irq[29]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 46.280 486.885 46.880 ;
    END
  END irq[2]
  PIN irq[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 465.160 486.885 465.760 ;
    END
  END irq[30]
  PIN irq[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 480.120 486.885 480.720 ;
    END
  END irq[31]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 61.240 486.885 61.840 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 76.200 486.885 76.800 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 91.160 486.885 91.760 ;
    END
  END irq[5]
  PIN irq[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 106.120 486.885 106.720 ;
    END
  END irq[6]
  PIN irq[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 121.080 486.885 121.680 ;
    END
  END irq[7]
  PIN irq[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 136.040 486.885 136.640 ;
    END
  END irq[8]
  PIN irq[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 482.885 151.000 486.885 151.600 ;
    END
  END irq[9]
  PIN mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END mem_addr[0]
  PIN mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END mem_addr[10]
  PIN mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END mem_addr[11]
  PIN mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END mem_addr[12]
  PIN mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END mem_addr[13]
  PIN mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END mem_addr[14]
  PIN mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END mem_addr[15]
  PIN mem_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END mem_addr[16]
  PIN mem_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END mem_addr[17]
  PIN mem_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END mem_addr[18]
  PIN mem_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END mem_addr[19]
  PIN mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END mem_addr[1]
  PIN mem_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END mem_addr[20]
  PIN mem_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END mem_addr[21]
  PIN mem_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END mem_addr[22]
  PIN mem_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END mem_addr[23]
  PIN mem_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END mem_addr[24]
  PIN mem_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END mem_addr[25]
  PIN mem_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END mem_addr[26]
  PIN mem_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END mem_addr[27]
  PIN mem_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END mem_addr[28]
  PIN mem_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END mem_addr[29]
  PIN mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END mem_addr[2]
  PIN mem_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END mem_addr[30]
  PIN mem_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END mem_addr[31]
  PIN mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END mem_addr[3]
  PIN mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END mem_addr[4]
  PIN mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END mem_addr[5]
  PIN mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END mem_addr[6]
  PIN mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END mem_addr[7]
  PIN mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END mem_addr[8]
  PIN mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END mem_addr[9]
  PIN mem_instr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END mem_instr
  PIN mem_la_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 493.605 89.610 497.605 ;
    END
  END mem_la_addr[0]
  PIN mem_la_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 107.730 493.605 108.010 497.605 ;
    END
  END mem_la_addr[10]
  PIN mem_la_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 109.570 493.605 109.850 497.605 ;
    END
  END mem_la_addr[11]
  PIN mem_la_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 111.410 493.605 111.690 497.605 ;
    END
  END mem_la_addr[12]
  PIN mem_la_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 113.250 493.605 113.530 497.605 ;
    END
  END mem_la_addr[13]
  PIN mem_la_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 115.090 493.605 115.370 497.605 ;
    END
  END mem_la_addr[14]
  PIN mem_la_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 116.930 493.605 117.210 497.605 ;
    END
  END mem_la_addr[15]
  PIN mem_la_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 118.770 493.605 119.050 497.605 ;
    END
  END mem_la_addr[16]
  PIN mem_la_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 120.610 493.605 120.890 497.605 ;
    END
  END mem_la_addr[17]
  PIN mem_la_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 122.450 493.605 122.730 497.605 ;
    END
  END mem_la_addr[18]
  PIN mem_la_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 124.290 493.605 124.570 497.605 ;
    END
  END mem_la_addr[19]
  PIN mem_la_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 493.605 91.450 497.605 ;
    END
  END mem_la_addr[1]
  PIN mem_la_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 126.130 493.605 126.410 497.605 ;
    END
  END mem_la_addr[20]
  PIN mem_la_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 127.970 493.605 128.250 497.605 ;
    END
  END mem_la_addr[21]
  PIN mem_la_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 129.810 493.605 130.090 497.605 ;
    END
  END mem_la_addr[22]
  PIN mem_la_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 131.650 493.605 131.930 497.605 ;
    END
  END mem_la_addr[23]
  PIN mem_la_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 133.490 493.605 133.770 497.605 ;
    END
  END mem_la_addr[24]
  PIN mem_la_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 135.330 493.605 135.610 497.605 ;
    END
  END mem_la_addr[25]
  PIN mem_la_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 137.170 493.605 137.450 497.605 ;
    END
  END mem_la_addr[26]
  PIN mem_la_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 139.010 493.605 139.290 497.605 ;
    END
  END mem_la_addr[27]
  PIN mem_la_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 140.850 493.605 141.130 497.605 ;
    END
  END mem_la_addr[28]
  PIN mem_la_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 142.690 493.605 142.970 497.605 ;
    END
  END mem_la_addr[29]
  PIN mem_la_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 93.010 493.605 93.290 497.605 ;
    END
  END mem_la_addr[2]
  PIN mem_la_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 144.530 493.605 144.810 497.605 ;
    END
  END mem_la_addr[30]
  PIN mem_la_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 146.370 493.605 146.650 497.605 ;
    END
  END mem_la_addr[31]
  PIN mem_la_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 94.850 493.605 95.130 497.605 ;
    END
  END mem_la_addr[3]
  PIN mem_la_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 96.690 493.605 96.970 497.605 ;
    END
  END mem_la_addr[4]
  PIN mem_la_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 98.530 493.605 98.810 497.605 ;
    END
  END mem_la_addr[5]
  PIN mem_la_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 100.370 493.605 100.650 497.605 ;
    END
  END mem_la_addr[6]
  PIN mem_la_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 102.210 493.605 102.490 497.605 ;
    END
  END mem_la_addr[7]
  PIN mem_la_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 104.050 493.605 104.330 497.605 ;
    END
  END mem_la_addr[8]
  PIN mem_la_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 105.890 493.605 106.170 497.605 ;
    END
  END mem_la_addr[9]
  PIN mem_la_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 26.770 493.605 27.050 497.605 ;
    END
  END mem_la_read
  PIN mem_la_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 30.450 493.605 30.730 497.605 ;
    END
  END mem_la_wdata[0]
  PIN mem_la_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 48.850 493.605 49.130 497.605 ;
    END
  END mem_la_wdata[10]
  PIN mem_la_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 50.690 493.605 50.970 497.605 ;
    END
  END mem_la_wdata[11]
  PIN mem_la_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 52.530 493.605 52.810 497.605 ;
    END
  END mem_la_wdata[12]
  PIN mem_la_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 54.370 493.605 54.650 497.605 ;
    END
  END mem_la_wdata[13]
  PIN mem_la_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 56.210 493.605 56.490 497.605 ;
    END
  END mem_la_wdata[14]
  PIN mem_la_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 58.050 493.605 58.330 497.605 ;
    END
  END mem_la_wdata[15]
  PIN mem_la_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 59.890 493.605 60.170 497.605 ;
    END
  END mem_la_wdata[16]
  PIN mem_la_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 61.730 493.605 62.010 497.605 ;
    END
  END mem_la_wdata[17]
  PIN mem_la_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 63.570 493.605 63.850 497.605 ;
    END
  END mem_la_wdata[18]
  PIN mem_la_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 65.410 493.605 65.690 497.605 ;
    END
  END mem_la_wdata[19]
  PIN mem_la_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 32.290 493.605 32.570 497.605 ;
    END
  END mem_la_wdata[1]
  PIN mem_la_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 67.250 493.605 67.530 497.605 ;
    END
  END mem_la_wdata[20]
  PIN mem_la_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 69.090 493.605 69.370 497.605 ;
    END
  END mem_la_wdata[21]
  PIN mem_la_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 70.930 493.605 71.210 497.605 ;
    END
  END mem_la_wdata[22]
  PIN mem_la_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 72.770 493.605 73.050 497.605 ;
    END
  END mem_la_wdata[23]
  PIN mem_la_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 74.610 493.605 74.890 497.605 ;
    END
  END mem_la_wdata[24]
  PIN mem_la_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 76.450 493.605 76.730 497.605 ;
    END
  END mem_la_wdata[25]
  PIN mem_la_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 78.290 493.605 78.570 497.605 ;
    END
  END mem_la_wdata[26]
  PIN mem_la_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 80.130 493.605 80.410 497.605 ;
    END
  END mem_la_wdata[27]
  PIN mem_la_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 81.970 493.605 82.250 497.605 ;
    END
  END mem_la_wdata[28]
  PIN mem_la_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 83.810 493.605 84.090 497.605 ;
    END
  END mem_la_wdata[29]
  PIN mem_la_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 34.130 493.605 34.410 497.605 ;
    END
  END mem_la_wdata[2]
  PIN mem_la_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 85.650 493.605 85.930 497.605 ;
    END
  END mem_la_wdata[30]
  PIN mem_la_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 87.490 493.605 87.770 497.605 ;
    END
  END mem_la_wdata[31]
  PIN mem_la_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 35.970 493.605 36.250 497.605 ;
    END
  END mem_la_wdata[3]
  PIN mem_la_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 37.810 493.605 38.090 497.605 ;
    END
  END mem_la_wdata[4]
  PIN mem_la_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 39.650 493.605 39.930 497.605 ;
    END
  END mem_la_wdata[5]
  PIN mem_la_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 41.490 493.605 41.770 497.605 ;
    END
  END mem_la_wdata[6]
  PIN mem_la_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 43.330 493.605 43.610 497.605 ;
    END
  END mem_la_wdata[7]
  PIN mem_la_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 45.170 493.605 45.450 497.605 ;
    END
  END mem_la_wdata[8]
  PIN mem_la_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 47.010 493.605 47.290 497.605 ;
    END
  END mem_la_wdata[9]
  PIN mem_la_write
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 28.610 493.605 28.890 497.605 ;
    END
  END mem_la_write
  PIN mem_la_wstrb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 148.210 493.605 148.490 497.605 ;
    END
  END mem_la_wstrb[0]
  PIN mem_la_wstrb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 150.050 493.605 150.330 497.605 ;
    END
  END mem_la_wstrb[1]
  PIN mem_la_wstrb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 151.890 493.605 152.170 497.605 ;
    END
  END mem_la_wstrb[2]
  PIN mem_la_wstrb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 153.730 493.605 154.010 497.605 ;
    END
  END mem_la_wstrb[3]
  PIN mem_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END mem_rdata[0]
  PIN mem_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END mem_rdata[10]
  PIN mem_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END mem_rdata[11]
  PIN mem_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END mem_rdata[12]
  PIN mem_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END mem_rdata[13]
  PIN mem_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END mem_rdata[14]
  PIN mem_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END mem_rdata[15]
  PIN mem_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END mem_rdata[16]
  PIN mem_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END mem_rdata[17]
  PIN mem_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END mem_rdata[18]
  PIN mem_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END mem_rdata[19]
  PIN mem_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END mem_rdata[1]
  PIN mem_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END mem_rdata[20]
  PIN mem_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END mem_rdata[21]
  PIN mem_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END mem_rdata[22]
  PIN mem_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END mem_rdata[23]
  PIN mem_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END mem_rdata[24]
  PIN mem_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END mem_rdata[25]
  PIN mem_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END mem_rdata[26]
  PIN mem_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END mem_rdata[27]
  PIN mem_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END mem_rdata[28]
  PIN mem_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END mem_rdata[29]
  PIN mem_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END mem_rdata[2]
  PIN mem_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END mem_rdata[30]
  PIN mem_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END mem_rdata[31]
  PIN mem_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END mem_rdata[3]
  PIN mem_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END mem_rdata[4]
  PIN mem_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END mem_rdata[5]
  PIN mem_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END mem_rdata[6]
  PIN mem_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END mem_rdata[7]
  PIN mem_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END mem_rdata[8]
  PIN mem_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END mem_rdata[9]
  PIN mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END mem_ready
  PIN mem_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END mem_valid
  PIN mem_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END mem_wdata[0]
  PIN mem_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END mem_wdata[10]
  PIN mem_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END mem_wdata[11]
  PIN mem_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END mem_wdata[12]
  PIN mem_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END mem_wdata[13]
  PIN mem_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END mem_wdata[14]
  PIN mem_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END mem_wdata[15]
  PIN mem_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END mem_wdata[16]
  PIN mem_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END mem_wdata[17]
  PIN mem_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END mem_wdata[18]
  PIN mem_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END mem_wdata[19]
  PIN mem_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END mem_wdata[1]
  PIN mem_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END mem_wdata[20]
  PIN mem_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END mem_wdata[21]
  PIN mem_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END mem_wdata[22]
  PIN mem_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END mem_wdata[23]
  PIN mem_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END mem_wdata[24]
  PIN mem_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END mem_wdata[25]
  PIN mem_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END mem_wdata[26]
  PIN mem_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END mem_wdata[27]
  PIN mem_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END mem_wdata[28]
  PIN mem_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END mem_wdata[29]
  PIN mem_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END mem_wdata[2]
  PIN mem_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END mem_wdata[30]
  PIN mem_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END mem_wdata[31]
  PIN mem_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END mem_wdata[3]
  PIN mem_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END mem_wdata[4]
  PIN mem_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END mem_wdata[5]
  PIN mem_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END mem_wdata[6]
  PIN mem_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END mem_wdata[7]
  PIN mem_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END mem_wdata[8]
  PIN mem_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END mem_wdata[9]
  PIN mem_wstrb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END mem_wstrb[0]
  PIN mem_wstrb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END mem_wstrb[1]
  PIN mem_wstrb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END mem_wstrb[2]
  PIN mem_wstrb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END mem_wstrb[3]
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END resetn
  PIN trace_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 493.605 396.890 497.605 ;
    END
  END trace_data[0]
  PIN trace_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 493.605 415.290 497.605 ;
    END
  END trace_data[10]
  PIN trace_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 493.605 417.130 497.605 ;
    END
  END trace_data[11]
  PIN trace_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 493.605 418.970 497.605 ;
    END
  END trace_data[12]
  PIN trace_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 493.605 420.810 497.605 ;
    END
  END trace_data[13]
  PIN trace_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 493.605 422.650 497.605 ;
    END
  END trace_data[14]
  PIN trace_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 493.605 424.490 497.605 ;
    END
  END trace_data[15]
  PIN trace_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 493.605 426.330 497.605 ;
    END
  END trace_data[16]
  PIN trace_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 493.605 428.170 497.605 ;
    END
  END trace_data[17]
  PIN trace_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 493.605 430.010 497.605 ;
    END
  END trace_data[18]
  PIN trace_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 493.605 431.850 497.605 ;
    END
  END trace_data[19]
  PIN trace_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 493.605 398.730 497.605 ;
    END
  END trace_data[1]
  PIN trace_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 493.605 433.690 497.605 ;
    END
  END trace_data[20]
  PIN trace_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 493.605 435.530 497.605 ;
    END
  END trace_data[21]
  PIN trace_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 493.605 437.370 497.605 ;
    END
  END trace_data[22]
  PIN trace_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 493.605 439.210 497.605 ;
    END
  END trace_data[23]
  PIN trace_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 493.605 441.050 497.605 ;
    END
  END trace_data[24]
  PIN trace_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 493.605 442.890 497.605 ;
    END
  END trace_data[25]
  PIN trace_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 493.605 444.730 497.605 ;
    END
  END trace_data[26]
  PIN trace_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 493.605 446.570 497.605 ;
    END
  END trace_data[27]
  PIN trace_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 493.605 448.410 497.605 ;
    END
  END trace_data[28]
  PIN trace_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 493.605 450.250 497.605 ;
    END
  END trace_data[29]
  PIN trace_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 493.605 400.570 497.605 ;
    END
  END trace_data[2]
  PIN trace_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 493.605 452.090 497.605 ;
    END
  END trace_data[30]
  PIN trace_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 493.605 453.930 497.605 ;
    END
  END trace_data[31]
  PIN trace_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 493.605 455.770 497.605 ;
    END
  END trace_data[32]
  PIN trace_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 493.605 457.610 497.605 ;
    END
  END trace_data[33]
  PIN trace_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 493.605 459.450 497.605 ;
    END
  END trace_data[34]
  PIN trace_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 493.605 461.290 497.605 ;
    END
  END trace_data[35]
  PIN trace_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 493.605 402.410 497.605 ;
    END
  END trace_data[3]
  PIN trace_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 493.605 404.250 497.605 ;
    END
  END trace_data[4]
  PIN trace_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 493.605 406.090 497.605 ;
    END
  END trace_data[5]
  PIN trace_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 493.605 407.930 497.605 ;
    END
  END trace_data[6]
  PIN trace_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 493.605 409.770 497.605 ;
    END
  END trace_data[7]
  PIN trace_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 493.605 411.610 497.605 ;
    END
  END trace_data[8]
  PIN trace_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 493.605 413.450 497.605 ;
    END
  END trace_data[9]
  PIN trace_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 493.605 395.050 497.605 ;
    END
  END trace_valid
  PIN trap
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 24.930 493.605 25.210 497.605 ;
    END
  END trap
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 481.160 484.245 ;
      LAYER met1 ;
        RECT 1.450 10.640 482.470 494.320 ;
      LAYER met2 ;
        RECT 1.480 493.325 24.650 494.350 ;
        RECT 25.490 493.325 26.490 494.350 ;
        RECT 27.330 493.325 28.330 494.350 ;
        RECT 29.170 493.325 30.170 494.350 ;
        RECT 31.010 493.325 32.010 494.350 ;
        RECT 32.850 493.325 33.850 494.350 ;
        RECT 34.690 493.325 35.690 494.350 ;
        RECT 36.530 493.325 37.530 494.350 ;
        RECT 38.370 493.325 39.370 494.350 ;
        RECT 40.210 493.325 41.210 494.350 ;
        RECT 42.050 493.325 43.050 494.350 ;
        RECT 43.890 493.325 44.890 494.350 ;
        RECT 45.730 493.325 46.730 494.350 ;
        RECT 47.570 493.325 48.570 494.350 ;
        RECT 49.410 493.325 50.410 494.350 ;
        RECT 51.250 493.325 52.250 494.350 ;
        RECT 53.090 493.325 54.090 494.350 ;
        RECT 54.930 493.325 55.930 494.350 ;
        RECT 56.770 493.325 57.770 494.350 ;
        RECT 58.610 493.325 59.610 494.350 ;
        RECT 60.450 493.325 61.450 494.350 ;
        RECT 62.290 493.325 63.290 494.350 ;
        RECT 64.130 493.325 65.130 494.350 ;
        RECT 65.970 493.325 66.970 494.350 ;
        RECT 67.810 493.325 68.810 494.350 ;
        RECT 69.650 493.325 70.650 494.350 ;
        RECT 71.490 493.325 72.490 494.350 ;
        RECT 73.330 493.325 74.330 494.350 ;
        RECT 75.170 493.325 76.170 494.350 ;
        RECT 77.010 493.325 78.010 494.350 ;
        RECT 78.850 493.325 79.850 494.350 ;
        RECT 80.690 493.325 81.690 494.350 ;
        RECT 82.530 493.325 83.530 494.350 ;
        RECT 84.370 493.325 85.370 494.350 ;
        RECT 86.210 493.325 87.210 494.350 ;
        RECT 88.050 493.325 89.050 494.350 ;
        RECT 89.890 493.325 90.890 494.350 ;
        RECT 91.730 493.325 92.730 494.350 ;
        RECT 93.570 493.325 94.570 494.350 ;
        RECT 95.410 493.325 96.410 494.350 ;
        RECT 97.250 493.325 98.250 494.350 ;
        RECT 99.090 493.325 100.090 494.350 ;
        RECT 100.930 493.325 101.930 494.350 ;
        RECT 102.770 493.325 103.770 494.350 ;
        RECT 104.610 493.325 105.610 494.350 ;
        RECT 106.450 493.325 107.450 494.350 ;
        RECT 108.290 493.325 109.290 494.350 ;
        RECT 110.130 493.325 111.130 494.350 ;
        RECT 111.970 493.325 112.970 494.350 ;
        RECT 113.810 493.325 114.810 494.350 ;
        RECT 115.650 493.325 116.650 494.350 ;
        RECT 117.490 493.325 118.490 494.350 ;
        RECT 119.330 493.325 120.330 494.350 ;
        RECT 121.170 493.325 122.170 494.350 ;
        RECT 123.010 493.325 124.010 494.350 ;
        RECT 124.850 493.325 125.850 494.350 ;
        RECT 126.690 493.325 127.690 494.350 ;
        RECT 128.530 493.325 129.530 494.350 ;
        RECT 130.370 493.325 131.370 494.350 ;
        RECT 132.210 493.325 133.210 494.350 ;
        RECT 134.050 493.325 135.050 494.350 ;
        RECT 135.890 493.325 136.890 494.350 ;
        RECT 137.730 493.325 138.730 494.350 ;
        RECT 139.570 493.325 140.570 494.350 ;
        RECT 141.410 493.325 142.410 494.350 ;
        RECT 143.250 493.325 144.250 494.350 ;
        RECT 145.090 493.325 146.090 494.350 ;
        RECT 146.930 493.325 147.930 494.350 ;
        RECT 148.770 493.325 149.770 494.350 ;
        RECT 150.610 493.325 151.610 494.350 ;
        RECT 152.450 493.325 153.450 494.350 ;
        RECT 154.290 493.325 155.290 494.350 ;
        RECT 156.130 493.325 157.130 494.350 ;
        RECT 157.970 493.325 158.970 494.350 ;
        RECT 159.810 493.325 160.810 494.350 ;
        RECT 161.650 493.325 162.650 494.350 ;
        RECT 163.490 493.325 164.490 494.350 ;
        RECT 165.330 493.325 166.330 494.350 ;
        RECT 167.170 493.325 168.170 494.350 ;
        RECT 169.010 493.325 170.010 494.350 ;
        RECT 170.850 493.325 171.850 494.350 ;
        RECT 172.690 493.325 173.690 494.350 ;
        RECT 174.530 493.325 175.530 494.350 ;
        RECT 176.370 493.325 177.370 494.350 ;
        RECT 178.210 493.325 179.210 494.350 ;
        RECT 180.050 493.325 181.050 494.350 ;
        RECT 181.890 493.325 182.890 494.350 ;
        RECT 183.730 493.325 184.730 494.350 ;
        RECT 185.570 493.325 186.570 494.350 ;
        RECT 187.410 493.325 188.410 494.350 ;
        RECT 189.250 493.325 190.250 494.350 ;
        RECT 191.090 493.325 192.090 494.350 ;
        RECT 192.930 493.325 193.930 494.350 ;
        RECT 194.770 493.325 195.770 494.350 ;
        RECT 196.610 493.325 197.610 494.350 ;
        RECT 198.450 493.325 199.450 494.350 ;
        RECT 200.290 493.325 201.290 494.350 ;
        RECT 202.130 493.325 203.130 494.350 ;
        RECT 203.970 493.325 204.970 494.350 ;
        RECT 205.810 493.325 206.810 494.350 ;
        RECT 207.650 493.325 208.650 494.350 ;
        RECT 209.490 493.325 210.490 494.350 ;
        RECT 211.330 493.325 212.330 494.350 ;
        RECT 213.170 493.325 214.170 494.350 ;
        RECT 215.010 493.325 216.010 494.350 ;
        RECT 216.850 493.325 217.850 494.350 ;
        RECT 218.690 493.325 219.690 494.350 ;
        RECT 220.530 493.325 221.530 494.350 ;
        RECT 222.370 493.325 223.370 494.350 ;
        RECT 224.210 493.325 225.210 494.350 ;
        RECT 226.050 493.325 227.050 494.350 ;
        RECT 227.890 493.325 228.890 494.350 ;
        RECT 229.730 493.325 230.730 494.350 ;
        RECT 231.570 493.325 232.570 494.350 ;
        RECT 233.410 493.325 234.410 494.350 ;
        RECT 235.250 493.325 236.250 494.350 ;
        RECT 237.090 493.325 238.090 494.350 ;
        RECT 238.930 493.325 239.930 494.350 ;
        RECT 240.770 493.325 241.770 494.350 ;
        RECT 242.610 493.325 243.610 494.350 ;
        RECT 244.450 493.325 245.450 494.350 ;
        RECT 246.290 493.325 247.290 494.350 ;
        RECT 248.130 493.325 249.130 494.350 ;
        RECT 249.970 493.325 250.970 494.350 ;
        RECT 251.810 493.325 252.810 494.350 ;
        RECT 253.650 493.325 254.650 494.350 ;
        RECT 255.490 493.325 256.490 494.350 ;
        RECT 257.330 493.325 258.330 494.350 ;
        RECT 259.170 493.325 260.170 494.350 ;
        RECT 261.010 493.325 262.010 494.350 ;
        RECT 262.850 493.325 263.850 494.350 ;
        RECT 264.690 493.325 265.690 494.350 ;
        RECT 266.530 493.325 267.530 494.350 ;
        RECT 268.370 493.325 269.370 494.350 ;
        RECT 270.210 493.325 271.210 494.350 ;
        RECT 272.050 493.325 273.050 494.350 ;
        RECT 273.890 493.325 274.890 494.350 ;
        RECT 275.730 493.325 276.730 494.350 ;
        RECT 277.570 493.325 278.570 494.350 ;
        RECT 279.410 493.325 280.410 494.350 ;
        RECT 281.250 493.325 282.250 494.350 ;
        RECT 283.090 493.325 284.090 494.350 ;
        RECT 284.930 493.325 285.930 494.350 ;
        RECT 286.770 493.325 287.770 494.350 ;
        RECT 288.610 493.325 289.610 494.350 ;
        RECT 290.450 493.325 291.450 494.350 ;
        RECT 292.290 493.325 293.290 494.350 ;
        RECT 294.130 493.325 295.130 494.350 ;
        RECT 295.970 493.325 296.970 494.350 ;
        RECT 297.810 493.325 298.810 494.350 ;
        RECT 299.650 493.325 300.650 494.350 ;
        RECT 301.490 493.325 302.490 494.350 ;
        RECT 303.330 493.325 304.330 494.350 ;
        RECT 305.170 493.325 306.170 494.350 ;
        RECT 307.010 493.325 308.010 494.350 ;
        RECT 308.850 493.325 309.850 494.350 ;
        RECT 310.690 493.325 311.690 494.350 ;
        RECT 312.530 493.325 313.530 494.350 ;
        RECT 314.370 493.325 315.370 494.350 ;
        RECT 316.210 493.325 317.210 494.350 ;
        RECT 318.050 493.325 319.050 494.350 ;
        RECT 319.890 493.325 320.890 494.350 ;
        RECT 321.730 493.325 322.730 494.350 ;
        RECT 323.570 493.325 324.570 494.350 ;
        RECT 325.410 493.325 326.410 494.350 ;
        RECT 327.250 493.325 328.250 494.350 ;
        RECT 329.090 493.325 330.090 494.350 ;
        RECT 330.930 493.325 331.930 494.350 ;
        RECT 332.770 493.325 333.770 494.350 ;
        RECT 334.610 493.325 335.610 494.350 ;
        RECT 336.450 493.325 337.450 494.350 ;
        RECT 338.290 493.325 339.290 494.350 ;
        RECT 340.130 493.325 341.130 494.350 ;
        RECT 341.970 493.325 342.970 494.350 ;
        RECT 343.810 493.325 344.810 494.350 ;
        RECT 345.650 493.325 346.650 494.350 ;
        RECT 347.490 493.325 348.490 494.350 ;
        RECT 349.330 493.325 350.330 494.350 ;
        RECT 351.170 493.325 352.170 494.350 ;
        RECT 353.010 493.325 354.010 494.350 ;
        RECT 354.850 493.325 355.850 494.350 ;
        RECT 356.690 493.325 357.690 494.350 ;
        RECT 358.530 493.325 359.530 494.350 ;
        RECT 360.370 493.325 361.370 494.350 ;
        RECT 362.210 493.325 363.210 494.350 ;
        RECT 364.050 493.325 365.050 494.350 ;
        RECT 365.890 493.325 366.890 494.350 ;
        RECT 367.730 493.325 368.730 494.350 ;
        RECT 369.570 493.325 370.570 494.350 ;
        RECT 371.410 493.325 372.410 494.350 ;
        RECT 373.250 493.325 374.250 494.350 ;
        RECT 375.090 493.325 376.090 494.350 ;
        RECT 376.930 493.325 377.930 494.350 ;
        RECT 378.770 493.325 379.770 494.350 ;
        RECT 380.610 493.325 381.610 494.350 ;
        RECT 382.450 493.325 383.450 494.350 ;
        RECT 384.290 493.325 385.290 494.350 ;
        RECT 386.130 493.325 387.130 494.350 ;
        RECT 387.970 493.325 388.970 494.350 ;
        RECT 389.810 493.325 390.810 494.350 ;
        RECT 391.650 493.325 392.650 494.350 ;
        RECT 393.490 493.325 394.490 494.350 ;
        RECT 395.330 493.325 396.330 494.350 ;
        RECT 397.170 493.325 398.170 494.350 ;
        RECT 399.010 493.325 400.010 494.350 ;
        RECT 400.850 493.325 401.850 494.350 ;
        RECT 402.690 493.325 403.690 494.350 ;
        RECT 404.530 493.325 405.530 494.350 ;
        RECT 406.370 493.325 407.370 494.350 ;
        RECT 408.210 493.325 409.210 494.350 ;
        RECT 410.050 493.325 411.050 494.350 ;
        RECT 411.890 493.325 412.890 494.350 ;
        RECT 413.730 493.325 414.730 494.350 ;
        RECT 415.570 493.325 416.570 494.350 ;
        RECT 417.410 493.325 418.410 494.350 ;
        RECT 419.250 493.325 420.250 494.350 ;
        RECT 421.090 493.325 422.090 494.350 ;
        RECT 422.930 493.325 423.930 494.350 ;
        RECT 424.770 493.325 425.770 494.350 ;
        RECT 426.610 493.325 427.610 494.350 ;
        RECT 428.450 493.325 429.450 494.350 ;
        RECT 430.290 493.325 431.290 494.350 ;
        RECT 432.130 493.325 433.130 494.350 ;
        RECT 433.970 493.325 434.970 494.350 ;
        RECT 435.810 493.325 436.810 494.350 ;
        RECT 437.650 493.325 438.650 494.350 ;
        RECT 439.490 493.325 440.490 494.350 ;
        RECT 441.330 493.325 442.330 494.350 ;
        RECT 443.170 493.325 444.170 494.350 ;
        RECT 445.010 493.325 446.010 494.350 ;
        RECT 446.850 493.325 447.850 494.350 ;
        RECT 448.690 493.325 449.690 494.350 ;
        RECT 450.530 493.325 451.530 494.350 ;
        RECT 452.370 493.325 453.370 494.350 ;
        RECT 454.210 493.325 455.210 494.350 ;
        RECT 456.050 493.325 457.050 494.350 ;
        RECT 457.890 493.325 458.890 494.350 ;
        RECT 459.730 493.325 460.730 494.350 ;
        RECT 461.570 493.325 482.450 494.350 ;
        RECT 1.480 4.280 482.450 493.325 ;
        RECT 1.480 4.000 121.250 4.280 ;
        RECT 122.090 4.000 364.590 4.280 ;
        RECT 365.430 4.000 482.450 4.280 ;
      LAYER met3 ;
        RECT 0.270 481.120 482.885 493.500 ;
        RECT 0.270 479.720 482.485 481.120 ;
        RECT 0.270 466.160 482.885 479.720 ;
        RECT 0.270 464.760 482.485 466.160 ;
        RECT 0.270 456.640 482.885 464.760 ;
        RECT 4.400 455.240 482.885 456.640 ;
        RECT 0.270 452.560 482.885 455.240 ;
        RECT 4.400 451.200 482.885 452.560 ;
        RECT 4.400 451.160 482.485 451.200 ;
        RECT 0.270 449.800 482.485 451.160 ;
        RECT 0.270 448.480 482.885 449.800 ;
        RECT 4.400 447.080 482.885 448.480 ;
        RECT 0.270 444.400 482.885 447.080 ;
        RECT 4.400 443.000 482.885 444.400 ;
        RECT 0.270 440.320 482.885 443.000 ;
        RECT 4.400 438.920 482.885 440.320 ;
        RECT 0.270 436.240 482.885 438.920 ;
        RECT 4.400 434.840 482.485 436.240 ;
        RECT 0.270 432.160 482.885 434.840 ;
        RECT 4.400 430.760 482.885 432.160 ;
        RECT 0.270 428.080 482.885 430.760 ;
        RECT 4.400 426.680 482.885 428.080 ;
        RECT 0.270 424.000 482.885 426.680 ;
        RECT 4.400 422.600 482.885 424.000 ;
        RECT 0.270 421.280 482.885 422.600 ;
        RECT 0.270 419.920 482.485 421.280 ;
        RECT 4.400 419.880 482.485 419.920 ;
        RECT 4.400 418.520 482.885 419.880 ;
        RECT 0.270 415.840 482.885 418.520 ;
        RECT 4.400 414.440 482.885 415.840 ;
        RECT 0.270 411.760 482.885 414.440 ;
        RECT 4.400 410.360 482.885 411.760 ;
        RECT 0.270 407.680 482.885 410.360 ;
        RECT 4.400 406.320 482.885 407.680 ;
        RECT 4.400 406.280 482.485 406.320 ;
        RECT 0.270 404.920 482.485 406.280 ;
        RECT 0.270 403.600 482.885 404.920 ;
        RECT 4.400 402.200 482.885 403.600 ;
        RECT 0.270 399.520 482.885 402.200 ;
        RECT 4.400 398.120 482.885 399.520 ;
        RECT 0.270 395.440 482.885 398.120 ;
        RECT 4.400 394.040 482.885 395.440 ;
        RECT 0.270 391.360 482.885 394.040 ;
        RECT 4.400 389.960 482.485 391.360 ;
        RECT 0.270 387.280 482.885 389.960 ;
        RECT 4.400 385.880 482.885 387.280 ;
        RECT 0.270 383.200 482.885 385.880 ;
        RECT 4.400 381.800 482.885 383.200 ;
        RECT 0.270 379.120 482.885 381.800 ;
        RECT 4.400 377.720 482.885 379.120 ;
        RECT 0.270 376.400 482.885 377.720 ;
        RECT 0.270 375.040 482.485 376.400 ;
        RECT 4.400 375.000 482.485 375.040 ;
        RECT 4.400 373.640 482.885 375.000 ;
        RECT 0.270 370.960 482.885 373.640 ;
        RECT 4.400 369.560 482.885 370.960 ;
        RECT 0.270 366.880 482.885 369.560 ;
        RECT 4.400 365.480 482.885 366.880 ;
        RECT 0.270 362.800 482.885 365.480 ;
        RECT 4.400 361.440 482.885 362.800 ;
        RECT 4.400 361.400 482.485 361.440 ;
        RECT 0.270 360.040 482.485 361.400 ;
        RECT 0.270 358.720 482.885 360.040 ;
        RECT 4.400 357.320 482.885 358.720 ;
        RECT 0.270 354.640 482.885 357.320 ;
        RECT 4.400 353.240 482.885 354.640 ;
        RECT 0.270 350.560 482.885 353.240 ;
        RECT 4.400 349.160 482.885 350.560 ;
        RECT 0.270 346.480 482.885 349.160 ;
        RECT 4.400 345.080 482.485 346.480 ;
        RECT 0.270 342.400 482.885 345.080 ;
        RECT 4.400 341.000 482.885 342.400 ;
        RECT 0.270 338.320 482.885 341.000 ;
        RECT 4.400 336.920 482.885 338.320 ;
        RECT 0.270 334.240 482.885 336.920 ;
        RECT 4.400 332.840 482.885 334.240 ;
        RECT 0.270 331.520 482.885 332.840 ;
        RECT 0.270 330.160 482.485 331.520 ;
        RECT 4.400 330.120 482.485 330.160 ;
        RECT 4.400 328.760 482.885 330.120 ;
        RECT 0.270 326.080 482.885 328.760 ;
        RECT 4.400 324.680 482.885 326.080 ;
        RECT 0.270 322.000 482.885 324.680 ;
        RECT 4.400 320.600 482.885 322.000 ;
        RECT 0.270 317.920 482.885 320.600 ;
        RECT 4.400 316.560 482.885 317.920 ;
        RECT 4.400 316.520 482.485 316.560 ;
        RECT 0.270 315.160 482.485 316.520 ;
        RECT 0.270 313.840 482.885 315.160 ;
        RECT 4.400 312.440 482.885 313.840 ;
        RECT 0.270 309.760 482.885 312.440 ;
        RECT 4.400 308.360 482.885 309.760 ;
        RECT 0.270 305.680 482.885 308.360 ;
        RECT 4.400 304.280 482.885 305.680 ;
        RECT 0.270 301.600 482.885 304.280 ;
        RECT 4.400 300.200 482.485 301.600 ;
        RECT 0.270 297.520 482.885 300.200 ;
        RECT 4.400 296.120 482.885 297.520 ;
        RECT 0.270 293.440 482.885 296.120 ;
        RECT 4.400 292.040 482.885 293.440 ;
        RECT 0.270 289.360 482.885 292.040 ;
        RECT 4.400 287.960 482.885 289.360 ;
        RECT 0.270 286.640 482.885 287.960 ;
        RECT 0.270 285.280 482.485 286.640 ;
        RECT 4.400 285.240 482.485 285.280 ;
        RECT 4.400 283.880 482.885 285.240 ;
        RECT 0.270 281.200 482.885 283.880 ;
        RECT 4.400 279.800 482.885 281.200 ;
        RECT 0.270 277.120 482.885 279.800 ;
        RECT 4.400 275.720 482.885 277.120 ;
        RECT 0.270 273.040 482.885 275.720 ;
        RECT 4.400 271.680 482.885 273.040 ;
        RECT 4.400 271.640 482.485 271.680 ;
        RECT 0.270 270.280 482.485 271.640 ;
        RECT 0.270 268.960 482.885 270.280 ;
        RECT 4.400 267.560 482.885 268.960 ;
        RECT 0.270 264.880 482.885 267.560 ;
        RECT 4.400 263.480 482.885 264.880 ;
        RECT 0.270 260.800 482.885 263.480 ;
        RECT 4.400 259.400 482.885 260.800 ;
        RECT 0.270 256.720 482.885 259.400 ;
        RECT 4.400 255.320 482.485 256.720 ;
        RECT 0.270 252.640 482.885 255.320 ;
        RECT 4.400 251.240 482.885 252.640 ;
        RECT 0.270 248.560 482.885 251.240 ;
        RECT 4.400 247.160 482.885 248.560 ;
        RECT 0.270 244.480 482.885 247.160 ;
        RECT 4.400 243.080 482.885 244.480 ;
        RECT 0.270 241.760 482.885 243.080 ;
        RECT 0.270 240.400 482.485 241.760 ;
        RECT 4.400 240.360 482.485 240.400 ;
        RECT 4.400 239.000 482.885 240.360 ;
        RECT 0.270 236.320 482.885 239.000 ;
        RECT 4.400 234.920 482.885 236.320 ;
        RECT 0.270 232.240 482.885 234.920 ;
        RECT 4.400 230.840 482.885 232.240 ;
        RECT 0.270 228.160 482.885 230.840 ;
        RECT 4.400 226.800 482.885 228.160 ;
        RECT 4.400 226.760 482.485 226.800 ;
        RECT 0.270 225.400 482.485 226.760 ;
        RECT 0.270 224.080 482.885 225.400 ;
        RECT 4.400 222.680 482.885 224.080 ;
        RECT 0.270 220.000 482.885 222.680 ;
        RECT 4.400 218.600 482.885 220.000 ;
        RECT 0.270 215.920 482.885 218.600 ;
        RECT 4.400 214.520 482.885 215.920 ;
        RECT 0.270 211.840 482.885 214.520 ;
        RECT 4.400 210.440 482.485 211.840 ;
        RECT 0.270 207.760 482.885 210.440 ;
        RECT 4.400 206.360 482.885 207.760 ;
        RECT 0.270 203.680 482.885 206.360 ;
        RECT 4.400 202.280 482.885 203.680 ;
        RECT 0.270 199.600 482.885 202.280 ;
        RECT 4.400 198.200 482.885 199.600 ;
        RECT 0.270 196.880 482.885 198.200 ;
        RECT 0.270 195.520 482.485 196.880 ;
        RECT 4.400 195.480 482.485 195.520 ;
        RECT 4.400 194.120 482.885 195.480 ;
        RECT 0.270 191.440 482.885 194.120 ;
        RECT 4.400 190.040 482.885 191.440 ;
        RECT 0.270 187.360 482.885 190.040 ;
        RECT 4.400 185.960 482.885 187.360 ;
        RECT 0.270 183.280 482.885 185.960 ;
        RECT 4.400 181.920 482.885 183.280 ;
        RECT 4.400 181.880 482.485 181.920 ;
        RECT 0.270 180.520 482.485 181.880 ;
        RECT 0.270 179.200 482.885 180.520 ;
        RECT 4.400 177.800 482.885 179.200 ;
        RECT 0.270 175.120 482.885 177.800 ;
        RECT 4.400 173.720 482.885 175.120 ;
        RECT 0.270 171.040 482.885 173.720 ;
        RECT 4.400 169.640 482.885 171.040 ;
        RECT 0.270 166.960 482.885 169.640 ;
        RECT 4.400 165.560 482.485 166.960 ;
        RECT 0.270 162.880 482.885 165.560 ;
        RECT 4.400 161.480 482.885 162.880 ;
        RECT 0.270 158.800 482.885 161.480 ;
        RECT 4.400 157.400 482.885 158.800 ;
        RECT 0.270 154.720 482.885 157.400 ;
        RECT 4.400 153.320 482.885 154.720 ;
        RECT 0.270 152.000 482.885 153.320 ;
        RECT 0.270 150.640 482.485 152.000 ;
        RECT 4.400 150.600 482.485 150.640 ;
        RECT 4.400 149.240 482.885 150.600 ;
        RECT 0.270 146.560 482.885 149.240 ;
        RECT 4.400 145.160 482.885 146.560 ;
        RECT 0.270 142.480 482.885 145.160 ;
        RECT 4.400 141.080 482.885 142.480 ;
        RECT 0.270 138.400 482.885 141.080 ;
        RECT 4.400 137.040 482.885 138.400 ;
        RECT 4.400 137.000 482.485 137.040 ;
        RECT 0.270 135.640 482.485 137.000 ;
        RECT 0.270 134.320 482.885 135.640 ;
        RECT 4.400 132.920 482.885 134.320 ;
        RECT 0.270 130.240 482.885 132.920 ;
        RECT 4.400 128.840 482.885 130.240 ;
        RECT 0.270 126.160 482.885 128.840 ;
        RECT 4.400 124.760 482.885 126.160 ;
        RECT 0.270 122.080 482.885 124.760 ;
        RECT 4.400 120.680 482.485 122.080 ;
        RECT 0.270 118.000 482.885 120.680 ;
        RECT 4.400 116.600 482.885 118.000 ;
        RECT 0.270 113.920 482.885 116.600 ;
        RECT 4.400 112.520 482.885 113.920 ;
        RECT 0.270 109.840 482.885 112.520 ;
        RECT 4.400 108.440 482.885 109.840 ;
        RECT 0.270 107.120 482.885 108.440 ;
        RECT 0.270 105.760 482.485 107.120 ;
        RECT 4.400 105.720 482.485 105.760 ;
        RECT 4.400 104.360 482.885 105.720 ;
        RECT 0.270 101.680 482.885 104.360 ;
        RECT 4.400 100.280 482.885 101.680 ;
        RECT 0.270 97.600 482.885 100.280 ;
        RECT 4.400 96.200 482.885 97.600 ;
        RECT 0.270 93.520 482.885 96.200 ;
        RECT 4.400 92.160 482.885 93.520 ;
        RECT 4.400 92.120 482.485 92.160 ;
        RECT 0.270 90.760 482.485 92.120 ;
        RECT 0.270 89.440 482.885 90.760 ;
        RECT 4.400 88.040 482.885 89.440 ;
        RECT 0.270 85.360 482.885 88.040 ;
        RECT 4.400 83.960 482.885 85.360 ;
        RECT 0.270 81.280 482.885 83.960 ;
        RECT 4.400 79.880 482.885 81.280 ;
        RECT 0.270 77.200 482.885 79.880 ;
        RECT 4.400 75.800 482.485 77.200 ;
        RECT 0.270 73.120 482.885 75.800 ;
        RECT 4.400 71.720 482.885 73.120 ;
        RECT 0.270 69.040 482.885 71.720 ;
        RECT 4.400 67.640 482.885 69.040 ;
        RECT 0.270 64.960 482.885 67.640 ;
        RECT 4.400 63.560 482.885 64.960 ;
        RECT 0.270 62.240 482.885 63.560 ;
        RECT 0.270 60.880 482.485 62.240 ;
        RECT 4.400 60.840 482.485 60.880 ;
        RECT 4.400 59.480 482.885 60.840 ;
        RECT 0.270 56.800 482.885 59.480 ;
        RECT 4.400 55.400 482.885 56.800 ;
        RECT 0.270 52.720 482.885 55.400 ;
        RECT 4.400 51.320 482.885 52.720 ;
        RECT 0.270 48.640 482.885 51.320 ;
        RECT 4.400 47.280 482.885 48.640 ;
        RECT 4.400 47.240 482.485 47.280 ;
        RECT 0.270 45.880 482.485 47.240 ;
        RECT 0.270 44.560 482.885 45.880 ;
        RECT 4.400 43.160 482.885 44.560 ;
        RECT 0.270 40.480 482.885 43.160 ;
        RECT 4.400 39.080 482.885 40.480 ;
        RECT 0.270 32.320 482.885 39.080 ;
        RECT 0.270 30.920 482.485 32.320 ;
        RECT 0.270 17.360 482.885 30.920 ;
        RECT 0.270 15.960 482.485 17.360 ;
        RECT 0.270 10.715 482.885 15.960 ;
      LAYER met4 ;
        RECT 0.295 484.800 462.465 493.505 ;
        RECT 0.295 13.095 20.640 484.800 ;
        RECT 23.040 13.095 97.440 484.800 ;
        RECT 99.840 13.095 174.240 484.800 ;
        RECT 176.640 13.095 251.040 484.800 ;
        RECT 253.440 13.095 327.840 484.800 ;
        RECT 330.240 13.095 404.640 484.800 ;
        RECT 407.040 13.095 462.465 484.800 ;
      LAYER met5 ;
        RECT 1.500 106.300 432.740 481.900 ;
  END
END alphacore
END LIBRARY

