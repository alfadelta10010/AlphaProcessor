* NGSPICE file created from spimemio.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

.subckt spimemio VGND VPWR addr[0] addr[10] addr[11] addr[12] addr[13] addr[14] addr[15]
+ addr[16] addr[17] addr[18] addr[19] addr[1] addr[20] addr[21] addr[22] addr[23]
+ addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] cfgreg_di[0] cfgreg_di[10]
+ cfgreg_di[11] cfgreg_di[12] cfgreg_di[13] cfgreg_di[14] cfgreg_di[15] cfgreg_di[16]
+ cfgreg_di[17] cfgreg_di[18] cfgreg_di[19] cfgreg_di[1] cfgreg_di[20] cfgreg_di[21]
+ cfgreg_di[22] cfgreg_di[23] cfgreg_di[24] cfgreg_di[25] cfgreg_di[26] cfgreg_di[27]
+ cfgreg_di[28] cfgreg_di[29] cfgreg_di[2] cfgreg_di[30] cfgreg_di[31] cfgreg_di[3]
+ cfgreg_di[4] cfgreg_di[5] cfgreg_di[6] cfgreg_di[7] cfgreg_di[8] cfgreg_di[9] cfgreg_do[0]
+ cfgreg_do[10] cfgreg_do[11] cfgreg_do[12] cfgreg_do[13] cfgreg_do[14] cfgreg_do[16]
+ cfgreg_do[17] cfgreg_do[18] cfgreg_do[19] cfgreg_do[1] cfgreg_do[20] cfgreg_do[21]
+ cfgreg_do[22] cfgreg_do[23] cfgreg_do[24] cfgreg_do[25] cfgreg_do[26] cfgreg_do[27]
+ cfgreg_do[28] cfgreg_do[29] cfgreg_do[2] cfgreg_do[31] cfgreg_do[3] cfgreg_do[4]
+ cfgreg_do[5] cfgreg_do[6] cfgreg_do[7] cfgreg_do[8] cfgreg_do[9] cfgreg_we[0] cfgreg_we[1]
+ cfgreg_we[2] cfgreg_we[3] clk flash_clk flash_csb flash_io0_di flash_io0_do flash_io0_oe
+ flash_io1_di flash_io1_do flash_io1_oe flash_io2_di flash_io2_do flash_io2_oe flash_io3_di
+ flash_io3_do flash_io3_oe rdata[0] rdata[10] rdata[11] rdata[12] rdata[13] rdata[14]
+ rdata[15] rdata[16] rdata[17] rdata[18] rdata[19] rdata[1] rdata[20] rdata[21] rdata[22]
+ rdata[23] rdata[24] rdata[25] rdata[26] rdata[27] rdata[28] rdata[29] rdata[2] rdata[30]
+ rdata[31] rdata[3] rdata[4] rdata[5] rdata[6] rdata[7] rdata[8] rdata[9] ready resetn
+ valid cfgreg_do[30] cfgreg_do[15]
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1295__2_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_778 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_934 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1518__B _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1390__B1 _0669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0956__B1 _0497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1381__B1 xfer.dout_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1270_ buffer\[0\] xfer.dout_data\[0\] _0715_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output56_A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0985_ config_qspi _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_898 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1606_ clknet_4_4_0_clk _0076_ VGND VGND VPWR VPWR xfer.din_valid sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1537_ rd_addr\[22\] _0306_ _0267_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1468_ _0376_ _0367_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_26_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1399_ _0201_ _0202_ _0620_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__o21a_1
XANTENNA__1124__B1 _0438_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_935 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1439__A rd_inc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0770_ rd_addr\[6\] net21 VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__xor2_2
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1322_ _0745_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1253_ xfer.din_data\[6\] _0703_ _0674_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__mux2_1
X_1184_ xfer.dout_data\[0\] net97 _0645_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_924 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_895 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
X_0968_ net2 VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0899_ xfer.dummy_count\[3\] xfer.dummy_count\[2\] xfer.dummy_count\[1\] xfer.dummy_count\[0\]
+ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__or4_4
XFILLER_0_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1259__A _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0822_ rd_addr\[10\] rd_addr\[11\] rd_addr\[12\] VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1592__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_166_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1305_ config_qspi net34 net45 VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1236_ xfer.din_data\[2\] _0674_ _0690_ _0673_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_526 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1167_ _0635_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__buf_4
XFILLER_0_66_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1098_ _0541_ xfer.obuffer\[1\] _0535_ xfer.obuffer\[4\] VGND VGND VPWR VPWR _0597_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1021_ _0547_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1088__A2 _0535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0805_ rd_addr\[8\] net23 VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1219_ net56 _0487_ state\[4\] _0499_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__a211o_1
XANTENNA__1079__A2 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1242__A2 _0503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1447__A rd_inc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1570_ clknet_4_1_0_clk _0040_ VGND VGND VPWR VPWR xfer.obuffer\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output86_A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1630__CLK clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1004_ _0535_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__buf_4
XANTENNA__0808__A2 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1466__C1 _0249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1481__A2 _0233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1233__A2 _0522_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1699_ clknet_4_2_0_clk _0148_ VGND VGND VPWR VPWR rd_addr\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1092__A _0585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0983__B2 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0983__A1 _0503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1653__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput75 net75 VGND VGND VPWR VPWR flash_io1_do sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput64 net64 VGND VGND VPWR VPWR cfgreg_do[2] sky130_fd_sc_hd__clkbuf_1
Xoutput53 net53 VGND VGND VPWR VPWR cfgreg_do[0] sky130_fd_sc_hd__clkbuf_1
Xoutput97 net97 VGND VGND VPWR VPWR rdata[24] sky130_fd_sc_hd__clkbuf_1
Xoutput86 net86 VGND VGND VPWR VPWR rdata[14] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1622_ clknet_4_13_0_clk _0092_ VGND VGND VPWR VPWR buffer\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__0974__B2 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1553_ clknet_4_14_0_clk _0023_ VGND VGND VPWR VPWR buffer\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1484_ net2 _0265_ _0237_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1676__CLK clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1390__B2 _0542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0956__A1 _0436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1381__A1 _0542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1381__B2 _0535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1549__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1699__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0984_ config_ddr VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__buf_4
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1605_ clknet_4_5_0_clk _0075_ VGND VGND VPWR VPWR xfer.resetn sky130_fd_sc_hd__dfxtp_1
X_1536_ net15 _0305_ rd_inc VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1354__B net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1467_ rd_addr\[6\] _0249_ _0252_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__a21bo_1
X_1398_ xfer.din_rd xfer.din_data\[1\] _0483_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1060__B1 _0571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_754 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1545__A _0669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1363__A1 xfer.dout_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1321_ _0361_ _0744_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__or2_1
X_1252_ _0686_ _0702_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1183_ _0653_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1290__B1 _0636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0967_ _0338_ net14 _0331_ _0340_ _0353_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1042__A0 xfer.dout_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0898_ xfer.xfer_dspi xfer.xfer_qspi VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__nor2_2
XFILLER_0_112_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1714__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1519_ net10 _0292_ rd_inc VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_805 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1259__B _0497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1441__C _0232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0821_ rd_addr\[8\] rd_addr\[9\] VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0801__B net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_166_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1304_ _0733_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1235_ net17 _0675_ _0689_ _0679_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__a211o_1
X_1166_ _0644_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_144_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1097_ _0596_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1034__S _0522_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1020_ config_do\[0\] _0546_ config_en VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__mux2_4
XFILLER_0_163_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0804_ rd_addr\[4\] VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_71_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1218_ state\[12\] _0455_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__and2_2
XANTENNA__1484__A0 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1149_ _0634_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1029__S _0522_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_532 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_666 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1582__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_119_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_963 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ _0534_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__buf_4
XFILLER_0_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0807__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1233__A3 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_808 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1698_ clknet_4_2_0_clk _0147_ VGND VGND VPWR VPWR rd_addr\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_12_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput65 net65 VGND VGND VPWR VPWR cfgreg_do[31] sky130_fd_sc_hd__clkbuf_1
Xoutput54 net54 VGND VGND VPWR VPWR cfgreg_do[10] sky130_fd_sc_hd__clkbuf_1
Xoutput76 net76 VGND VGND VPWR VPWR flash_io1_oe sky130_fd_sc_hd__clkbuf_1
Xoutput98 net98 VGND VGND VPWR VPWR rdata[25] sky130_fd_sc_hd__clkbuf_1
Xoutput87 net87 VGND VGND VPWR VPWR rdata[15] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1448__A0 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1621_ clknet_4_13_0_clk _0091_ VGND VGND VPWR VPWR buffer\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__0974__A2 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1552_ clknet_4_11_0_clk _0022_ VGND VGND VPWR VPWR buffer\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1483_ _0419_ _0264_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_145_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_154_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1390__A2 _0526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_163_Left_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1042__S _0559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1620__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1381__A2 xfer.dout_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1741__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0983_ _0503_ _0481_ _0485_ _0499_ _0521_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1604_ clknet_4_14_0_clk _0074_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1535_ _0382_ _0304_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1466_ _0726_ _0250_ _0251_ _0249_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__a211o_1
X_1397_ _0199_ _0200_ _0483_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1124__A2 _0454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1643__CLK clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1736__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1320_ net59 net31 net45 VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1251_ net6 _0528_ _0675_ net21 _0701_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__a221o_1
X_1182_ buffer\[23\] net96 _0645_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__mux2_1
XANTENNA__1666__CLK clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0966_ _0318_ _0347_ _0348_ _0504_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__nor4_1
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0897_ _0440_ _0441_ _0442_ _0443_ xfer.count\[3\] VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1518_ rd_addr\[18\] _0373_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1449_ rd_addr\[2\] _0238_ _0629_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_528 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1320__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1689__CLK clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1441__D _0479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1272__A1 xfer.dout_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0820_ rd_addr\[6\] rd_addr\[7\] VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_951 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1303_ _0731_ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__and2_1
X_1234_ _0687_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__or2_1
X_1165_ buffer\[15\] net87 _0636_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1096_ _0595_ xfer.obuffer\[4\] _0571_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1140__S _0629_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0949_ _0434_ rd_wait VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_861 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1050__S _0559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1190__A0 xfer.dout_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1704__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1297__4 clknet_4_1_0_clk VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__inv_2
XFILLER_0_38_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0803_ _0347_ _0348_ _0349_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1135__S _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1217_ state\[0\] _0671_ _0673_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1148_ _0363_ xfer.dout_tag\[1\] xfer.dout_tag\[2\] _0557_ VGND VGND VPWR VPWR _0634_
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_88_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1079_ xfer.obuffer\[0\] _0536_ _0482_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_622 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1475__A1 _0232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_840 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1744__A net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1463__B _0363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0910__B1 _0363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1002_ _0465_ _0445_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__and2_2
XFILLER_0_88_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1466__A1 _0726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0823__A _0366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1697_ clknet_4_13_0_clk _0146_ VGND VGND VPWR VPWR rd_addr\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_954 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput55 net55 VGND VGND VPWR VPWR cfgreg_do[11] sky130_fd_sc_hd__clkbuf_1
Xoutput66 net66 VGND VGND VPWR VPWR cfgreg_do[3] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput99 net99 VGND VGND VPWR VPWR rdata[26] sky130_fd_sc_hd__clkbuf_1
Xoutput88 net88 VGND VGND VPWR VPWR rdata[16] sky130_fd_sc_hd__clkbuf_1
Xoutput77 net77 VGND VGND VPWR VPWR flash_io2_do sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1503__S _0267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0908__A _0438_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_670 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1739__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1620_ clknet_4_4_0_clk _0090_ VGND VGND VPWR VPWR din_ddr sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_786 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1551_ clknet_4_14_0_clk _0021_ VGND VGND VPWR VPWR buffer\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1482_ rd_addr\[10\] _0402_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1572__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_165_Right_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0982_ _0436_ _0520_ _0497_ _0500_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_119_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1595__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1603_ clknet_4_15_0_clk _0073_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dfxtp_1
XANTENNA__1357__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1534_ rd_addr\[22\] _0430_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1465_ _0726_ net21 VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1396_ _0448_ xfer.dummy_count\[1\] xfer.dummy_count\[0\] VGND VGND VPWR VPWR _0200_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_96_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1060__A2 _0526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_924 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1289__A rd_inc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1250_ config_qspi _0499_ _0503_ net15 VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__a22o_1
X_1181_ _0652_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1290__A2 _0363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0965_ _0319_ _0320_ _0323_ _0358_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0896_ xfer.xfer_dspi xfer.count\[1\] VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1517_ _0291_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_149_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1448_ net17 _0236_ _0237_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1502__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1610__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1379_ _0188_ xfer.dout_data\[5\] _0174_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1048__S _0559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0916__A xfer.count\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_963 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1482__A rd_addr\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1302_ _0522_ net35 net45 VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__mux2_1
X_1233_ config_qspi _0522_ _0499_ _0528_ net2 VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_144_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1164_ _0643_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1095_ xfer.din_data\[4\] _0594_ _0455_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0948_ state\[7\] _0437_ _0491_ _0481_ state\[4\] VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__a32o_1
XFILLER_0_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1420__C1 _0585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0879_ _0396_ _0398_ _0417_ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1392__A _0526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1656__CLK clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0802_ rd_addr\[18\] net10 VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_146_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1216_ _0670_ _0672_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__or2_2
X_1147_ _0633_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1151__S _0636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1078_ _0581_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1679__CLK clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0995__B2 _0530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1475__A2 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_634 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1163__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ xfer.dummy_count\[3\] xfer.dummy_count\[2\] xfer.dummy_count\[1\] xfer.dummy_count\[0\]
+ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__nor4_4
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1696_ clknet_4_13_0_clk _0145_ VGND VGND VPWR VPWR rd_addr\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_38_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1146__S _0629_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput56 net56 VGND VGND VPWR VPWR cfgreg_do[16] sky130_fd_sc_hd__clkbuf_1
Xoutput67 net67 VGND VGND VPWR VPWR cfgreg_do[4] sky130_fd_sc_hd__clkbuf_1
Xoutput89 net89 VGND VGND VPWR VPWR rdata[17] sky130_fd_sc_hd__clkbuf_1
Xoutput78 net78 VGND VGND VPWR VPWR flash_io2_oe sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0908__B _0454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_922 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1550_ clknet_4_14_0_clk _0020_ VGND VGND VPWR VPWR buffer\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output84_A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1481_ net24 _0233_ _0263_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_59_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1375__A1 xfer.dout_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1717__CLK clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_640 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1748_ config_en VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1679_ clknet_4_9_0_clk xfer.xfer_tag\[1\] VGND VGND VPWR VPWR xfer.dout_tag\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_77_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_696 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1366__A1 xfer.dout_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_95_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0981_ state\[9\] _0519_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1054__A0 xfer.dout_data\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_754 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1602_ clknet_4_15_0_clk _0072_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1357__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1533_ _0303_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1464_ rd_addr\[6\] _0376_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0829__A _0366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1395_ _0448_ xfer.dummy_count\[0\] xfer.dummy_count\[1\] VGND VGND VPWR VPWR _0199_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0859__B1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_581 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1180_ buffer\[22\] net95 _0645_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__mux2_1
XANTENNA__1511__A1 _0726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1562__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0964_ state\[9\] VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0895_ xfer.count\[0\] xfer.xfer_dspi VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_41_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1516_ rd_addr\[17\] _0290_ _0267_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1447_ rd_inc VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__buf_4
XFILLER_0_156_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1378_ xfer.dout_data\[3\] _0592_ _0187_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1585__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1257__B1 _0698_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1301_ net51 VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__clkbuf_2
X_1232_ net58 _0487_ _0503_ net10 VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_144_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1163_ buffer\[14\] net86 _0636_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1094_ xfer.obuffer\[2\] _0592_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1003__A _0534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0947_ _0489_ _0490_ _0457_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_42_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0878_ _0420_ _0421_ _0422_ _0423_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_3_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_699 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_917 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_894 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0801_ rd_addr\[22\] net15 VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1600__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1402__B1 _0456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1215_ _0487_ state\[12\] state\[9\] _0663_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__nor4_1
XFILLER_0_46_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1146_ net110 buffer\[7\] _0629_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1077_ buffer\[23\] xfer.dout_data\[7\] _0573_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_861 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1623__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0910__A2 _0437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1000_ _0532_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_141_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1695_ clknet_4_4_0_clk _0144_ VGND VGND VPWR VPWR xfer.flash_csb sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_38_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_9_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1646__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1129_ xfer.dout_tag\[1\] xfer.dout_tag\[2\] _0479_ _0557_ VGND VGND VPWR VPWR _0623_
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_95_639 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput57 net57 VGND VGND VPWR VPWR cfgreg_do[17] sky130_fd_sc_hd__clkbuf_1
Xoutput79 net79 VGND VGND VPWR VPWR flash_io3_do sky130_fd_sc_hd__clkbuf_1
Xoutput68 net68 VGND VGND VPWR VPWR cfgreg_do[5] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0924__B xfer.count\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ _0262_ rd_addr\[9\] _0249_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1669__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0850__A _0333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1157__S _0636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1747_ config_ddr VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1678_ clknet_4_12_0_clk xfer.xfer_tag\[0\] VGND VGND VPWR VPWR xfer.dout_tag\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1063__A1 xfer.dout_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1067__S _0573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1366__A2 _0592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0980_ _0505_ _0510_ _0518_ _0434_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1601_ clknet_4_15_0_clk _0071_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1532_ rd_addr\[21\] _0302_ _0267_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1463_ xfer.dout_tag\[1\] _0363_ _0724_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__or3_4
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1109__A2 _0535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1394_ _0197_ _0198_ _0620_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0845__A _0333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1293__A1 _0726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1293__B2 _0363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1284__A1 xfer.dout_data\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1511__A2 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1707__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1296__3_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0963_ state\[10\] _0437_ _0502_ _0485_ state\[4\] VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0894_ xfer.xfer_qspi xfer.flash_clk VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1515_ net9 _0289_ _0237_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1446_ rd_addr\[2\] VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__inv_1
XFILLER_0_156_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1377_ _0542_ xfer.dout_data\[1\] xfer.dout_data\[4\] _0536_ VGND VGND VPWR VPWR
+ _0187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1170__S _0645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1009__A1 config_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1300_ _0730_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1231_ _0670_ _0684_ _0686_ _0674_ xfer.din_data\[1\] VGND VGND VPWR VPWR _0081_
+ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_144_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1162_ _0642_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1093_ _0541_ xfer.obuffer\[0\] xfer.obuffer\[3\] _0534_ VGND VGND VPWR VPWR _0593_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1248__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0946_ xfer.last_fetch xfer.xfer_ddr_q xfer.fetch VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_71_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1420__A1 _0534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0877_ _0321_ _0399_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__xnor2_1
XANTENNA__1225__B1_N _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1165__S _0636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1184__A0 xfer.dout_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1429_ state\[8\] state\[11\] _0226_ _0227_ _0500_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_71_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1239__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1075__S _0573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1552__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0800_ rd_addr\[12\] net4 VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__xor2_2
XFILLER_0_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1214_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1145_ _0632_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1076_ _0580_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_5_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0999__S config_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_160_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0929_ _0451_ _0461_ _0474_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1575__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_670 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0910__A3 _0456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1320__A0 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_934 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1598__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1694_ clknet_4_4_0_clk _0143_ VGND VGND VPWR VPWR xfer.flash_clk sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0848__A _0333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1311__A0 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1128_ _0622_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1059_ _0454_ _0569_ _0570_ _0438_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_76_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_606 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput58 net58 VGND VGND VPWR VPWR cfgreg_do[18] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput69 net69 VGND VGND VPWR VPWR cfgreg_do[8] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1302__A0 _0522_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1369__B1 xfer.dout_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1528__S _0267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1541__B1 _0636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1746_ config_qspi VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1677_ clknet_4_10_0_clk _0129_ VGND VGND VPWR VPWR xfer.dout_data\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1613__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1523__B1 _0232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_13_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1600_ clknet_4_14_0_clk _0070_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1258__S _0530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1531_ _0232_ net14 _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__a21o_1
XANTENNA__1636__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1462_ _0248_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1393_ xfer.din_rd xfer.din_data\[0\] _0483_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1293__A2 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1022__A _0538_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1168__S _0645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_724 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1659__CLK clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_142_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0962_ _0491_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0893_ xfer.count\[0\] xfer.count\[1\] VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1514_ rd_addr\[17\] _0383_ _0373_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_160_Left_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1445_ _0235_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1376_ _0186_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1451__S _0237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_724 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0766__A rd_addr\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1009__A2 _0533_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1536__S rd_inc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1230_ _0685_ _0487_ _0455_ _0672_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__a31o_1
X_1161_ buffer\[13\] net85 _0636_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1092_ _0585_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__buf_4
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0945_ _0444_ _0447_ _0452_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0876_ net23 _0399_ _0400_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1428_ xfer.din_tag\[0\] _0226_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1359_ _0438_ _0569_ _0173_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__nand3_4
XFILLER_0_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1239__A2 _0487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1411__A2 _0459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1213_ _0363_ _0520_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_53_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1144_ net109 buffer\[6\] _0629_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1075_ buffer\[22\] xfer.dout_data\[6\] _0573_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_930 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0928_ _0448_ _0451_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__nand2_1
XANTENNA__1176__S _0645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0859_ _0404_ _0405_ net19 VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1086__S _0571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0938__B _0483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_946 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1084__B1 _0585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1387__A1 xfer.dout_data\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1693_ clknet_4_4_0_clk _0142_ VGND VGND VPWR VPWR xfer.xfer_dspi sky130_fd_sc_hd__dfxtp_2
XFILLER_0_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_29_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1127_ _0465_ _0457_ xfer.fetch VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__or3_1
XFILLER_0_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1058_ xfer.xfer_ddr _0464_ _0568_ _0459_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__a211o_1
XFILLER_0_165_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1398__C _0483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1378__A1 xfer.dout_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1692__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput59 net59 VGND VGND VPWR VPWR cfgreg_do[19] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1369__A1 _0542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1369__B2 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1541__A1 _0726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1565__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1745_ config_cont VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1676_ clknet_4_10_0_clk _0128_ VGND VGND VPWR VPWR xfer.dout_data\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_68_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1048__A0 xfer.dout_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1588__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1211__B1 _0669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output82_A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1530_ _0232_ _0428_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_73_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1461_ rd_addr\[5\] _0247_ _0629_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1392_ _0526_ _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1303__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0861__B _0345_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1449__S _0629_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1184__S _0645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1659_ clknet_4_7_0_clk _0008_ VGND VGND VPWR VPWR state\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1213__A _0363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0771__B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0962__A _0491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0961_ state\[11\] _0481_ _0485_ state\[5\] VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1603__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0892_ xfer.din_valid VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__clkinv_2
XFILLER_0_140_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1513_ _0288_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_149_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1444_ rd_addr\[1\] net12 _0233_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1375_ _0185_ xfer.dout_data\[4\] _0174_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0766__B net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1626__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1009__A3 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1089__S _0456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1160_ _0641_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_144_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1091_ _0591_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1248__A3 _0456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0944_ xfer.fetch xfer.xfer_ddr_q VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0875_ _0319_ _0419_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1427_ state\[3\] _0492_ _0520_ _0225_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_10_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1649__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1358_ xfer.xfer_ddr _0464_ _0448_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__a21o_1
X_1289_ rd_inc VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1239__A3 _0483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_833 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0777__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_864 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1120__B _0533_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1212_ xfer.din_tag\[2\] _0526_ _0669_ xfer.xfer_tag\[2\] VGND VGND VPWR VPWR _0079_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_53_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1143_ _0631_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
X_1074_ _0579_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0927_ xfer.count\[3\] _0472_ _0459_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0858_ rd_addr\[2\] rd_addr\[3\] rd_addr\[4\] VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0789_ rd_addr\[3\] VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_914 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1093__B2 _0534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1093__A1 _0541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1367__S _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0938__C _0479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0954__B _0491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1692_ clknet_4_4_0_clk _0141_ VGND VGND VPWR VPWR xfer.xfer_ddr sky130_fd_sc_hd__dfxtp_2
XFILLER_0_151_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1306__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1126_ xfer.count\[3\] _0544_ _0609_ _0621_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__o31a_1
XFILLER_0_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1057_ _0447_ _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__nor2_4
XANTENNA__1075__A1 xfer.dout_data\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_914 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1378__A2 _0592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0889__A1 _0427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1369__A2 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1744_ net80 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1675_ clknet_4_10_0_clk _0127_ VGND VGND VPWR VPWR xfer.dout_data\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_110_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1036__A _0556_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ xfer.obuffer\[6\] _0535_ _0482_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1202__C state\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1220__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0934__A_N _0436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1220__B2 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_623 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_950 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1460_ _0726_ net20 _0246_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__o21a_1
XANTENNA_output75_A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1391_ _0459_ xfer.dummy_count\[0\] VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1278__A1 xfer.dout_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1682__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1658_ clknet_4_7_0_clk _0007_ VGND VGND VPWR VPWR state\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1589_ clknet_4_15_0_clk _0059_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1375__S _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_931 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1555__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output113_A net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0960_ _0363_ _0498_ _0501_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_7_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0891_ xfer.resetn VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1196__A0 xfer.dout_data\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1512_ rd_addr\[16\] _0287_ _0267_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1443_ _0234_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_149_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1374_ xfer.dout_data\[2\] _0592_ _0184_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__a21o_1
XANTENNA__1499__A1 _0333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_612 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1578__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_783 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1350__A0 config_do\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1090_ _0590_ xfer.obuffer\[3\] _0571_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1720__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0943_ state\[12\] _0485_ _0486_ _0481_ _0487_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_924 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0874_ rd_addr\[11\] _0348_ _0419_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_840 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1309__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1426_ _0667_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__inv_2
X_1357_ net47 net48 _0536_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1341__A0 config_do\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1288_ rd_valid _0725_ _0437_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_526 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xspimemio_120 VGND VGND VPWR VPWR spimemio_120/HI cfgreg_do[23] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_161_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_139_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_867 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0968__A net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1211_ xfer.din_tag\[1\] _0526_ _0669_ xfer.xfer_tag\[1\] VGND VGND VPWR VPWR _0078_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_53_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1142_ net108 buffer\[5\] _0629_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1073_ buffer\[21\] xfer.dout_data\[5\] _0573_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_148_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0926_ _0470_ _0458_ _0471_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_157_Left_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0857_ rd_addr\[2\] rd_addr\[3\] rd_addr\[4\] VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0788_ net18 VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1616__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1409_ xfer.count\[1\] VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__inv_1
XANTENNA__1314__A0 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_166_Left_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_926 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1514__B1_N _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1383__S _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0788__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1305__A0 config_qspi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1084__A2 _0535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0990__A_N _0436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1691_ clknet_4_6_0_clk _0140_ VGND VGND VPWR VPWR xfer.din_tag\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__1639__CLK clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1125_ _0438_ _0619_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1056_ _0440_ _0458_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__nor2_2
XFILLER_0_146_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_926 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0909_ _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_14 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1743_ net78 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1674_ clknet_4_10_0_clk _0126_ VGND VGND VPWR VPWR xfer.dout_data\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_124_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0973__D1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1108_ _0541_ xfer.obuffer\[3\] _0585_ xfer.obuffer\[5\] VGND VGND VPWR VPWR _0605_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1039_ _0557_ _0558_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_101_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1220__A2 _0503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1523__A3 _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1211__A2 _0526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_112_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0970__B2 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1390_ xfer.din_qspi _0526_ _0669_ _0542_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_130_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1657_ clknet_4_3_0_clk _0006_ VGND VGND VPWR VPWR state\[3\] sky130_fd_sc_hd__dfxtp_1
X_1588_ clknet_4_14_0_clk _0058_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_718 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_941 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ _0363_ _0436_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__nor2_4
XFILLER_0_83_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1432__A2 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1511_ _0726_ net8 _0286_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1442_ rd_addr\[0\] net1 _0233_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__mux2_1
XANTENNA__0943__B2 _0487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1373_ _0542_ xfer.dout_data\[0\] xfer.dout_data\[3\] _0536_ VGND VGND VPWR VPWR
+ _0184_ sky130_fd_sc_hd__a22o_1
XANTENNA__1499__A2 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1330__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1476__S _0629_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1709_ clknet_4_9_0_clk _0158_ VGND VGND VPWR VPWR rd_addr\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1672__CLK clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1415__A _0438_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0942_ state\[1\] VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0873_ rd_addr\[11\] _0419_ _0348_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_97_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1425_ _0224_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1356_ _0438_ _0453_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__nand2_1
X_1287_ xfer.dout_tag\[1\] _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1695__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xspimemio_121 VGND VGND VPWR VPWR spimemio_121/HI cfgreg_do[24] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_161_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0843__B1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_843 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1020__A0 config_do\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1210_ xfer.din_tag\[0\] _0526_ _0669_ xfer.xfer_tag\[0\] VGND VGND VPWR VPWR _0077_
+ sky130_fd_sc_hd__a22o_1
X_1141_ _0630_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1568__CLK clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1072_ _0578_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0834__B1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0925_ _0451_ xfer.count\[3\] VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0856_ _0314_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0787_ rd_addr\[20\] _0332_ _0333_ _0334_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_23_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1408_ _0209_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1339_ net51 _0756_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1250__B1 _0503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0792__A_N net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1710__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_696 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1690_ clknet_4_3_0_clk _0139_ VGND VGND VPWR VPWR xfer.din_tag\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1544__A1 _0459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1124_ _0446_ _0454_ _0438_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__o21a_1
X_1055_ _0567_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1232__B1 _0503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0908_ _0438_ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__nand2_4
XFILLER_0_31_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0839_ _0316_ _0382_ _0384_ _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__1484__S _0237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0774__D _0321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0982__C1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_26 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0981__B _0519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1606__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1742_ net76 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1673_ clknet_4_10_0_clk _0125_ VGND VGND VPWR VPWR xfer.dout_data\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1333__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1107_ _0604_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1038_ xfer.dout_tag\[2\] _0479_ xfer.dout_tag\[1\] VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__and3b_1
XFILLER_0_165_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_894 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1508__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1629__CLK clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1435__B1 _0669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1656_ clknet_4_6_0_clk _0005_ VGND VGND VPWR VPWR state\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1587_ clknet_4_14_0_clk _0057_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_498 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1148__A _0363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1510_ _0285_ _0383_ _0237_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output80_A net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1441_ _0724_ xfer.dout_tag\[1\] _0232_ _0479_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_49_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1372_ _0183_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_945 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_730 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1708_ clknet_4_8_0_clk _0157_ VGND VGND VPWR VPWR rd_addr\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1639_ clknet_4_7_0_clk _0105_ VGND VGND VPWR VPWR config_cont sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1415__B _0478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0941_ config_qspi config_ddr VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0872_ _0418_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_97_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_899 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1424_ _0438_ _0478_ _0223_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1355_ _0171_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1286_ xfer.dout_tag\[2\] _0557_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__nand2_1
XANTENNA__0883__C _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xspimemio_122 VGND VGND VPWR VPWR spimemio_122/HI cfgreg_do[25] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_161_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1297__4_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1129__C _0479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1140_ net107 buffer\[4\] _0629_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1071_ buffer\[20\] xfer.dout_data\[4\] _0573_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_775 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1100__S _0455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0924_ xfer.count\[0\] xfer.count\[1\] VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0855_ _0376_ _0367_ _0368_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0786_ net5 VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1336__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1407_ _0620_ _0208_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1338_ config_clk net39 net43 VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1269_ _0714_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1662__CLK clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_723 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1250__B2 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1250__A1 config_qspi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_89_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_98_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1069__A1 xfer.dout_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_164_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1544__A2 _0533_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1685__CLK clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1123_ xfer.count\[3\] _0614_ _0615_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__a211o_1
X_1054_ xfer.dout_data\[7\] buffer\[15\] _0559_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1232__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0907_ _0439_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__nor2_8
XFILLER_0_114_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1232__B2 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0838_ _0327_ _0383_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0769_ _0315_ _0316_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0844__S _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1471__A1 _0726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_870 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1558__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0799__B net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0982__B1 _0497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1741_ net74 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1672_ clknet_4_10_0_clk _0124_ VGND VGND VPWR VPWR xfer.dout_data\[2\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1106_ _0603_ xfer.obuffer\[6\] _0571_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1037_ xfer.dout_tag\[0\] _0491_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_859 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1700__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1495__S _0267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_614 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1508__A2 _0233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1524__A _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0955__B1 config_cont VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1655_ clknet_4_7_0_clk _0004_ VGND VGND VPWR VPWR state\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1586_ clknet_4_11_0_clk _0056_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1362__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1440_ _0231_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1371_ _0182_ xfer.dout_data\[3\] _0174_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1339__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1707_ clknet_4_8_0_clk _0156_ VGND VGND VPWR VPWR rd_addr\[11\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_113_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1619__CLK clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1638_ clknet_4_7_0_clk _0104_ VGND VGND VPWR VPWR config_qspi sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ clknet_4_0_0_clk _0039_ VGND VGND VPWR VPWR xfer.obuffer\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__1344__A0 config_do\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_637 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0940_ state\[5\] _0481_ _0485_ state\[8\] VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0871_ rd_addr\[10\] _0366_ _0367_ _0368_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_97_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_640 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1423_ _0569_ _0613_ _0221_ _0222_ _0451_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_118_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1354_ _0537_ net46 _0361_ _0170_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__or4_1
X_1285_ _0723_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_127_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_550 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1591__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1317__A0 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xspimemio_123 VGND VGND VPWR VPWR spimemio_123/HI cfgreg_do[26] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_143_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1308__A0 config_cont VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1070_ _0577_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0923_ _0465_ xfer.xfer_qspi VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0854_ _0399_ _0400_ net23 VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0785_ rd_addr\[13\] VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1406_ xfer.din_rd xfer.din_data\[3\] _0483_ _0478_ _0207_ VGND VGND VPWR VPWR _0208_
+ sky130_fd_sc_hd__a32o_1
X_1337_ _0755_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1268_ xfer.dout_tag\[0\] _0479_ _0491_ _0713_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1199_ _0661_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1250__A2 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_144_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1262__A _0437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_153_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1226__C1 state\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1544__A3 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1122_ _0465_ _0541_ _0473_ _0616_ _0617_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__a311o_1
X_1053_ _0566_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1111__S _0571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1232__A2 _0487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0906_ _0444_ _0447_ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__or3_2
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0837_ _0327_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0768_ rd_addr\[23\] net16 VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0982__A1 _0436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_727 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_863 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1740_ net72 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1671_ clknet_4_10_0_clk _0123_ VGND VGND VPWR VPWR xfer.dout_data\[1\] sky130_fd_sc_hd__dfxtp_4
XANTENNA__0973__A1 _0333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_963 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1652__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1106__S _0571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1105_ xfer.din_data\[6\] _0602_ _0455_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1036_ _0556_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1429__C1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1675__CLK clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0955__A1 _0427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1295__2 clknet_4_0_0_clk VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__inv_2
X_1654_ clknet_4_3_0_clk _0000_ VGND VGND VPWR VPWR state\[0\] sky130_fd_sc_hd__dfxtp_1
X_1585_ clknet_4_14_0_clk _0055_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1371__A1 xfer.dout_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1548__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_635 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ xfer.flash_io0_do xfer_io0_90 _0522_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1698__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1362__A1 xfer.dout_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1050__A0 xfer.dout_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1370_ xfer.dout_data\[1\] _0592_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1706_ clknet_4_8_0_clk _0155_ VGND VGND VPWR VPWR rd_addr\[10\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1637_ clknet_4_7_0_clk _0103_ VGND VGND VPWR VPWR config_ddr sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1568_ clknet_4_1_0_clk _0038_ VGND VGND VPWR VPWR xfer.obuffer\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1499_ _0333_ _0624_ _0277_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1265__A _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1713__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0870_ _0401_ _0403_ _0408_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__and4_1
XFILLER_0_82_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1422_ _0542_ _0536_ _0462_ _0569_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_3_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1353_ net43 net44 net45 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__or3_1
X_1284_ buffer\[7\] xfer.dout_data\[7\] _0715_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0999_ config_clk _0459_ config_en VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_779 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xspimemio_124 VGND VGND VPWR VPWR spimemio_124/HI cfgreg_do[27] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_143_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1024__S _0522_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1609__CLK clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0922_ xfer.count\[0\] _0463_ _0464_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__o31a_1
XFILLER_0_43_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0853_ _0376_ _0367_ rd_addr\[8\] VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0784_ net13 VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1405_ xfer.dummy_count\[3\] _0203_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__xor2_1
X_1336_ net51 _0754_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_108_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 addr[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_160_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1267_ xfer.dout_tag\[1\] xfer.dout_tag\[2\] VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1198_ xfer.dout_data\[7\] net105 _0635_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1019__S _0522_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1121_ _0612_ xfer.count\[3\] _0585_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__nor3b_1
X_1052_ xfer.dout_data\[6\] buffer\[14\] _0559_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1581__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_700 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0905_ _0448_ _0449_ _0450_ _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0976__C1 _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0836_ _0333_ rd_addr\[16\] _0365_ _0371_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__and4_1
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0991__A2 _0437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0767_ rd_addr\[19\] net11 VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1319_ _0743_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_123_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_614 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1302__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_941 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1670_ clknet_4_10_0_clk _0122_ VGND VGND VPWR VPWR xfer.dout_data\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output96_A net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1104_ xfer.obuffer\[4\] _0592_ _0601_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1035_ config_do\[3\] _0555_ config_en VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__mux2_4
XFILLER_0_146_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0819_ rd_addr\[2\] rd_addr\[3\] rd_addr\[4\] rd_addr\[5\] VGND VGND VPWR VPWR _0366_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_13_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1435__A3 _0526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1653_ clknet_4_5_0_clk _0119_ VGND VGND VPWR VPWR config_do\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1584_ clknet_4_14_0_clk _0054_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1018_ xfer.obuffer\[7\] _0466_ _0545_ VGND VGND VPWR VPWR xfer.flash_io0_do sky130_fd_sc_hd__o21a_1
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1642__CLK clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output59_A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1705_ clknet_4_8_0_clk _0154_ VGND VGND VPWR VPWR rd_addr\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_53_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1636_ clknet_4_5_0_clk _0102_ VGND VGND VPWR VPWR config_en sky130_fd_sc_hd__dfxtp_4
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1567_ clknet_4_0_0_clk _0037_ VGND VGND VPWR VPWR xfer.obuffer\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1498_ _0624_ _0276_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_506 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1665__CLK clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0803__C_N _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1280__A1 xfer.dout_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1265__B _0497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1421_ _0465_ _0541_ _0475_ _0220_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a31o_1
X_1352_ _0765_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
X_1283_ _0722_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__1688__CLK clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_149_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0998_ _0531_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_6
XFILLER_0_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1619_ clknet_4_6_0_clk _0089_ VGND VGND VPWR VPWR xfer.din_rd sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_165_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1305__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xspimemio_125 VGND VGND VPWR VPWR spimemio_125/HI cfgreg_do[28] sky130_fd_sc_hd__conb_1
Xspimemio_114 VGND VGND VPWR VPWR spimemio_114/HI cfgreg_do[6] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_143_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1040__S _0559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1253__A1 _0703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1244__A1 _0696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0921_ xfer.count\[0\] _0448_ xfer.count\[1\] _0466_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0852_ rd_addr\[8\] _0366_ _0367_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0802__B net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0783_ net13 rd_addr\[20\] VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_77_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1404_ _0205_ _0206_ _0620_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1335_ config_csb net40 net43 VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 addr[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_160_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1266_ _0712_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
X_1197_ _0660_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1235__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1703__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1035__S config_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1226__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1226__B2 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1120_ xfer.xfer_ddr _0533_ _0445_ _0460_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__and4_1
XFILLER_0_88_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1051_ _0565_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0904_ xfer.count\[2\] VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__buf_2
XFILLER_0_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0835_ rd_addr\[21\] rd_addr\[22\] _0375_ _0373_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_12_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0766_ rd_addr\[10\] net2 VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_94_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0991__A3 _0526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1318_ _0731_ _0742_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1249_ xfer.din_data\[5\] _0674_ _0698_ _0700_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__o22a_1
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1103_ _0541_ xfer.obuffer\[2\] _0535_ xfer.obuffer\[5\] VGND VGND VPWR VPWR _0601_
+ sky130_fd_sc_hd__a22o_1
X_1034_ xfer.flash_io3_do xfer_io3_90 _0522_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_8_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0818_ rd_addr\[14\] rd_addr\[15\] VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_133_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_924 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1268__B _0479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1365__B1 xfer.dout_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1571__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1652_ clknet_4_5_0_clk _0118_ VGND VGND VPWR VPWR config_do\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1583_ clknet_4_11_0_clk _0053_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0810__B net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1108__B1 _0585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1133__S _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1017_ _0449_ xfer.obuffer\[4\] _0464_ xfer.obuffer\[6\] _0544_ VGND VGND VPWR VPWR
+ _0545_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1594__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1308__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1347__A0 config_do\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_31_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1742__A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1510__B1 _0237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0805__B net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0821__A rd_addr\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1704_ clknet_4_8_0_clk _0153_ VGND VGND VPWR VPWR rd_addr\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1635_ net131 xfer.flash_io3_do VGND VGND VPWR VPWR xfer_io3_90 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1566_ clknet_4_0_0_clk _0036_ VGND VGND VPWR VPWR xfer.obuffer\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1497_ _0334_ _0388_ _0726_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_724 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0791__B2 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1099__A2 _0592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1737__A net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1420_ _0534_ _0218_ _0219_ _0460_ _0585_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a221o_1
XANTENNA_output71_A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1351_ net51 _0764_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__and2_1
X_1282_ buffer\[6\] xfer.dout_data\[6\] _0715_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0997_ config_csb xfer.flash_csb config_en VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1618_ clknet_4_5_0_clk _0088_ VGND VGND VPWR VPWR xfer.din_qspi sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1549_ clknet_4_11_0_clk _0019_ VGND VGND VPWR VPWR buffer\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_105_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xspimemio_126 VGND VGND VPWR VPWR spimemio_126/HI cfgreg_do[29] sky130_fd_sc_hd__conb_1
Xspimemio_115 VGND VGND VPWR VPWR spimemio_115/HI cfgreg_do[7] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_2_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_805 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1292__A _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_123_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0920_ _0465_ _0445_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__nand2_2
XFILLER_0_166_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0851_ _0328_ _0397_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0782_ _0314_ _0317_ _0322_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_77_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1655__CLK clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1403_ xfer.din_rd xfer.din_data\[2\] _0483_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1334_ _0753_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1265_ _0500_ _0497_ _0711_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_160_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 addr[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_4
X_1196_ xfer.dout_data\[6\] net104 _0635_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1226__A2 _0503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1678__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_941 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1050_ xfer.dout_data\[5\] buffer\[13\] _0559_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_830 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0903_ xfer.xfer_ddr xfer.xfer_qspi VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0834_ _0374_ _0379_ net13 VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_4_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1317_ net58 net30 net45 VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1248_ net20 state\[12\] _0456_ _0699_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1121__C_N _0585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1179_ _0651_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1046__S _0559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1745__A config_cont VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1383__A1 xfer.dout_data\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1102_ _0600_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1033_ _0554_ VGND VGND VPWR VPWR xfer.flash_io3_do sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1438__A2 _0478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0817_ rd_addr\[16\] rd_addr\[17\] VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput50 flash_io3_di VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_133_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1374__A1 xfer.dout_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1268__C _0491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1716__CLK clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1365__B2 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1365__A1 _0542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0909__A _0455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1720_ clknet_4_4_0_clk _0169_ VGND VGND VPWR VPWR xfer.count\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1651_ clknet_4_5_0_clk _0117_ VGND VGND VPWR VPWR config_do\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1582_ clknet_4_12_0_clk _0052_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1108__A1 _0541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1016_ xfer.xfer_ddr _0445_ _0446_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1044__A0 xfer.dout_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1035__A0 config_do\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_12_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1703_ clknet_4_2_0_clk _0152_ VGND VGND VPWR VPWR rd_addr\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1634_ net130 xfer.flash_io2_do VGND VGND VPWR VPWR xfer_io2_90 sky130_fd_sc_hd__dfxtp_1
X_1565_ clknet_4_0_0_clk _0035_ VGND VGND VPWR VPWR xfer.obuffer\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _0275_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1144__S _0629_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1561__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0791__A2 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1054__S _0559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1205__C_N _0519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1350_ config_do\[3\] net38 net43 VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__mux2_1
X_1281_ _0721_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1584__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0996_ state\[12\] _0481_ _0485_ _0528_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1617_ clknet_4_3_0_clk _0087_ VGND VGND VPWR VPWR xfer.din_data\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_165_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1548_ clknet_4_11_0_clk _0018_ VGND VGND VPWR VPWR buffer\[9\] sky130_fd_sc_hd__dfxtp_1
X_1479_ rd_addr\[9\] _0399_ _0261_ _0726_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__o211a_1
Xspimemio_127 VGND VGND VPWR VPWR spimemio_127/HI cfgreg_do[30] sky130_fd_sc_hd__conb_1
Xspimemio_116 VGND VGND VPWR VPWR spimemio_116/HI cfgreg_do[12] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_2_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1486__A0 rd_addr\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1292__B _0436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1512__S _0267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1748__A config_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ _0333_ _0371_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0781_ _0323_ _0324_ _0327_ _0328_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_77_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1402_ _0203_ _0204_ _0456_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1333_ _0731_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__and2_1
X_1264_ din_ddr _0522_ _0530_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 addr[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1195_ _0659_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_0_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0979_ _0512_ _0513_ _0515_ _0517_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1459__B1 _0237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_780 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1507__S _0249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_842 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1622__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0902_ xfer.xfer_qspi VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__clkinv_2
XFILLER_0_43_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0833_ net13 _0374_ _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__and3_1
XANTENNA__0976__A2 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1316_ _0741_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1247_ net14 _0503_ _0528_ net5 VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__a22o_1
X_1178_ buffer\[21\] net94 _0645_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0967__A2 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1645__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_155_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1101_ _0599_ xfer.obuffer\[5\] _0571_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1032_ _0541_ xfer.obuffer\[7\] _0533_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__and3_1
XFILLER_0_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1071__A1 xfer.dout_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_141_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput40 cfgreg_di[5] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0816_ _0362_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__clkbuf_4
Xinput51 resetn VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1374__A2 _0592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_150_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1668__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1365__A2 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1520__S _0267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_672 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1650_ clknet_4_5_0_clk _0116_ VGND VGND VPWR VPWR config_do\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1581_ clknet_4_11_0_clk _0051_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1015_ config_oe\[3\] _0537_ _0543_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__a21o_4
XFILLER_0_44_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1515__S _0237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1274__A1 xfer.dout_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1702_ clknet_4_2_0_clk _0151_ VGND VGND VPWR VPWR rd_addr\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1633_ net129 xfer.flash_io1_do VGND VGND VPWR VPWR xfer_io1_90 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1564_ clknet_4_2_0_clk _0034_ VGND VGND VPWR VPWR xfer.obuffer\[1\] sky130_fd_sc_hd__dfxtp_1
X_1495_ rd_addr\[12\] _0274_ _0267_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1706__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1396__A _0448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1256__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1192__A0 xfer.dout_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1280_ buffer\[5\] xfer.dout_data\[5\] _0715_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__mux2_1
XANTENNA_output57_A net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1247__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1247__B2 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ _0528_ _0481_ _0485_ _0530_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1616_ clknet_4_2_0_clk _0086_ VGND VGND VPWR VPWR xfer.din_data\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1155__S _0636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1547_ clknet_4_11_0_clk _0017_ VGND VGND VPWR VPWR buffer\[8\] sky130_fd_sc_hd__dfxtp_1
X_1478_ _0402_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__inv_2
Xspimemio_117 VGND VGND VPWR VPWR spimemio_117/HI cfgreg_do[13] sky130_fd_sc_hd__conb_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1238__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1238__B2 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_894 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1065__S _0573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0921__B1 xfer.count\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0780_ rd_addr\[14\] net6 VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_77_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1401_ xfer.dummy_count\[2\] _0200_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1551__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1332_ config_oe\[3\] net27 net44 VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__mux2_1
X_1263_ _0710_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_160_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput5 addr[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
XFILLER_0_36_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1194_ xfer.dout_data\[5\] net102 _0635_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1004__A _0535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0978_ _0516_ _0321_ _0324_ _0315_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1574__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0928__A _0448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0901_ xfer.flash_clk VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0832_ _0375_ _0364_ _0365_ _0378_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__nand4_2
XFILLER_0_98_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1315_ _0731_ _0740_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_140_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1246_ _0499_ _0486_ _0673_ state\[4\] _0679_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__a2111o_1
X_1177_ _0650_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1597__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1377__B1 xfer.dout_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0914__C xfer.count\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1080__A2 _0456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_1100_ xfer.din_data\[5\] _0598_ _0455_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1031_ _0553_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 cfgreg_di[18] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0840__B _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0815_ _0361_ softreset VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput52 valid VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_4
Xinput41 cfgreg_di[8] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_133_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1163__S _0636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1229_ config_cont VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1073__S _0573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1612__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_721 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0941__A config_qspi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1580_ clknet_4_11_0_clk _0050_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output87_A net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ config_oe\[2\] _0537_ _0543_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__a21o_4
XFILLER_0_158_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_640 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1012__A _0541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1201__C1 _0437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0997__S config_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0936__A _0438_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_941 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1701_ clknet_4_2_0_clk _0150_ VGND VGND VPWR VPWR rd_addr\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__1431__C1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1658__CLK clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1632_ net128 xfer.flash_io0_do VGND VGND VPWR VPWR xfer_io0_90 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1563_ clknet_4_14_0_clk _0033_ VGND VGND VPWR VPWR buffer\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1494_ _0232_ net4 _0272_ _0273_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_930 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_759 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1247__A2 _0503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0994_ _0529_ _0519_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__nor2_2
XFILLER_0_70_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1615_ clknet_4_3_0_clk _0085_ VGND VGND VPWR VPWR xfer.din_data\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1546_ _0313_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_165_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1477_ _0260_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
Xspimemio_118 VGND VGND VPWR VPWR spimemio_118/HI cfgreg_do[14] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_2_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1238__A2 _0503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1081__S _0571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1400_ xfer.dummy_count\[2\] _0200_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__nor2_1
XANTENNA__1165__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1331_ _0751_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
X_1262_ _0437_ _0709_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_160_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 addr[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_160_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1193_ _0658_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_125_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0977_ rd_addr\[23\] net16 VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1393__C _0483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1529_ _0300_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_145_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1719__CLK clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1395__A1 _0448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ xfer.xfer_ddr _0445_ _0446_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0831_ _0376_ _0367_ _0368_ _0377_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1386__A1 xfer.dout_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1314_ net57 net29 net45 VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__mux2_1
X_1245_ _0697_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
X_1176_ buffer\[20\] net93 _0645_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1377__B2 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1377__A1 _0542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1691__CLK clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1030_ config_do\[2\] _0552_ config_en VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__mux2_4
XFILLER_0_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput20 addr[5] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
XFILLER_0_72_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0814_ net51 VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__clkinv_2
Xinput31 cfgreg_di[19] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput42 cfgreg_di[9] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1444__S _0233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1531__A1 _0232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1228_ net57 _0487_ _0483_ _0683_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1159_ buffer\[12\] net84 _0636_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__mux2_1
XANTENNA__1564__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1522__A1 _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_644 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1210__B1 _0669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1264__S _0530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1587__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1013_ xfer.xfer_rd config_en _0533_ _0542_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_157_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_919 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1174__S _0645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_836 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0936__B _0454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0952__A _0437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1700_ clknet_4_2_0_clk _0149_ VGND VGND VPWR VPWR rd_addr\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1631_ clknet_4_12_0_clk _0101_ VGND VGND VPWR VPWR rd_inc sky130_fd_sc_hd__dfxtp_2
XFILLER_0_2_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1562_ clknet_4_15_0_clk _0032_ VGND VGND VPWR VPWR buffer\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_894 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1493_ rd_addr\[11\] _0419_ rd_addr\[12\] VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1602__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_147_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1489__A0 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_156_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1256__A3 _0456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_165_Left_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1625__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0993_ _0503_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_833 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1614_ clknet_4_2_0_clk _0084_ VGND VGND VPWR VPWR xfer.din_data\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1545_ _0669_ _0311_ _0312_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_165_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_163_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1476_ rd_addr\[8\] _0259_ _0629_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1452__S _0629_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xspimemio_119 VGND VGND VPWR VPWR spimemio_119/HI cfgreg_do[15] sky130_fd_sc_hd__conb_1
XFILLER_0_66_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_588 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0921__A2 _0448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1362__S _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1648__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_728 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1537__S _0267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1330_ _0731_ _0750_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__and2_1
X_1261_ _0438_ _0487_ _0454_ xfer.din_rd VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__a31o_1
X_1192_ xfer.dout_data\[4\] net101 _0635_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 addr[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
XFILLER_0_79_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1301__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0976_ _0514_ net2 _0328_ _0349_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_693 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1528_ rd_addr\[20\] _0299_ _0267_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1182__S _0645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1459_ _0376_ _0245_ _0237_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_52_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1357__S _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0830_ rd_addr\[10\] rd_addr\[11\] rd_addr\[12\] _0333_ VGND VGND VPWR VPWR _0377_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_25_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1386__A2 _0592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_102_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1313_ _0739_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
X_1244_ xfer.din_data\[4\] _0696_ _0674_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1175_ _0649_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1031__A _0553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_111_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1377__A2 xfer.dout_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0959_ _0436_ _0456_ _0499_ _0500_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__and4b_1
XFILLER_0_43_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_120_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1065__A1 xfer.dout_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput10 addr[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 addr[6] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
X_0813_ _0330_ _0346_ _0360_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__nor3_2
XFILLER_0_4_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput43 cfgreg_we[0] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
XFILLER_0_25_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput32 cfgreg_di[1] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1531__A2 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1026__A _0550_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1227_ net12 _0675_ _0681_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1158_ _0640_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__1709__CLK clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1089_ xfer.din_data\[3\] _0589_ _0456_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_870 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_867 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1012_ _0541_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0835__D _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_728 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1455__S _0237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1681__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1630_ clknet_4_9_0_clk _0100_ VGND VGND VPWR VPWR rd_wait sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1561_ clknet_4_15_0_clk _0031_ VGND VGND VPWR VPWR buffer\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1554__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1492_ _0232_ _0371_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1007__C _0538_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1422__A1 _0542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1186__A0 xfer.dout_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_750 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0772__B net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1413__B2 _0535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1577__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1095__S _0455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0992_ state\[6\] VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1613_ clknet_4_3_0_clk _0083_ VGND VGND VPWR VPWR xfer.din_data\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1544_ _0459_ _0533_ _0536_ _0460_ xfer.count\[0\] VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_165_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1475_ _0232_ net23 _0258_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0767__B net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0958__A _0479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1260_ _0708_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
X_1191_ _0657_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
Xinput8 addr[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_160_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0975_ rd_addr\[10\] VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1389__B1 _0669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1527_ _0232_ net13 _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__a21o_1
X_1458_ rd_addr\[5\] _0404_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_52_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1389_ xfer.din_rd _0526_ _0669_ xfer.xfer_rd VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1615__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_924 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1312_ _0731_ _0738_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1243_ net19 _0675_ _0686_ _0695_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_140_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1174_ buffer\[19\] net91 _0645_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1312__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1059__C1 _0438_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0958_ _0479_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0889_ _0427_ _0433_ _0435_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_70_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1638__CLK clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1222__A _0487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0780__B net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1116__B xfer.count\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0971__A _0345_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput11 addr[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
XFILLER_0_108_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput22 addr[7] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
X_0812_ _0351_ _0357_ _0358_ _0359_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__or4b_1
XFILLER_0_71_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput33 cfgreg_di[20] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput44 cfgreg_we[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1226_ net9 _0503_ _0528_ net24 state\[4\] VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1157_ buffer\[11\] net83 _0636_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1088_ xfer.obuffer\[2\] _0535_ _0585_ xfer.obuffer\[1\] VGND VGND VPWR VPWR _0589_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_723 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0775__B net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1210__A2 _0526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1011_ xfer.xfer_qspi VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0960__A1 _0363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0876__A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1209_ _0457_ _0454_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__nor2_4
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0786__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1560_ clknet_4_15_0_clk _0030_ VGND VGND VPWR VPWR buffer\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_718 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output85_A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1491_ _0271_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_810 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1422__A2 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1689_ clknet_4_6_0_clk _0138_ VGND VGND VPWR VPWR xfer.din_tag\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_148_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1413__A2 _0585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ state\[0\] _0437_ _0526_ _0527_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1612_ clknet_4_3_0_clk _0082_ VGND VGND VPWR VPWR xfer.din_data\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1671__CLK clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1543_ _0211_ _0446_ _0466_ _0461_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_165_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1474_ _0231_ _0399_ _0400_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1315__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1159__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1209__B _0454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0783__B rd_addr\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1694__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1119__B _0542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1190_ xfer.dout_data\[3\] net100 _0635_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 addr[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XFILLER_0_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0974_ _0337_ net18 _0354_ net5 _0350_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1526_ rd_inc _0374_ _0379_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1457_ _0244_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
X_1388_ _0195_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0884__A _0349_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1567__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_777 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1311_ net56 net28 net45 VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__mux2_1
X_1242_ net13 _0503_ _0528_ net4 _0694_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_14 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1173_ _0648_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_858 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0957_ state\[2\] VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput110 net110 VGND VGND VPWR VPWR rdata[7] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0888_ _0434_ net113 rd_valid VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__or3b_2
XFILLER_0_88_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1509_ rd_addr\[16\] _0395_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1298__A0 config_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1222__B _0455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1525__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput12 addr[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
X_0811_ _0352_ net19 net52 rd_valid VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput23 addr[8] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
XFILLER_0_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput34 cfgreg_di[21] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput45 cfgreg_we[2] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1225_ config_qspi _0522_ _0499_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_79_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1156_ _0639_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1087_ _0588_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1605__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1379__S _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_51_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1010_ config_oe\[1\] _0537_ _0539_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__a21bo_4
XANTENNA__1628__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_931 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_874 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1318__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1037__B _0491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1208_ _0668_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1139_ _0623_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_727 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0951__A2 _0483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_920 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1490_ rd_addr\[11\] _0270_ _0267_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output78_A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1688_ clknet_4_1_0_clk _0137_ VGND VGND VPWR VPWR xfer.count\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0887__A net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1110__A2 _0456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_134_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_143_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0990_ _0436_ _0502_ state\[7\] _0500_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__and4b_1
XFILLER_0_39_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1611_ clknet_4_3_0_clk _0081_ VGND VGND VPWR VPWR xfer.din_data\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1542_ rd_addr\[23\] _0624_ _0308_ _0310_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1473_ _0257_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_143_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1387__S _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_917 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0973_ _0333_ _0334_ _0511_ rd_valid net52 VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_70_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1389__A2 _0526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1525_ net11 _0233_ _0295_ _0297_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1456_ rd_addr\[4\] _0243_ _0629_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__mux2_1
X_1387_ _0194_ xfer.dout_data\[7\] _0174_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1077__A1 xfer.dout_data\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1661__CLK clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_723 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_970 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1310_ _0737_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
X_1241_ config_qspi _0522_ _0499_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__and3b_1
XANTENNA__0985__A config_qspi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ buffer\[18\] net90 _0645_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1059__A1 _0454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0956_ _0436_ _0496_ _0497_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput100 net100 VGND VGND VPWR VPWR rdata[27] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0887_ net52 VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput111 net111 VGND VGND VPWR VPWR rdata[8] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1508_ net7 _0233_ _0284_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1490__S _0267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1439_ rd_inc VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__inv_2
XANTENNA__1241__A_N config_qspi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1684__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0959__A_N _0436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1525__A2 _0233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput13 addr[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
X_0810_ rd_addr\[16\] net8 VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__xor2_2
XFILLER_0_71_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput24 addr[9] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput35 cfgreg_di[22] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput46 cfgreg_we[3] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_141_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1557__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1224_ xfer.din_data\[0\] _0674_ _0680_ _0673_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1155_ buffer\[10\] net82 _0636_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1086_ _0587_ xfer.obuffer\[2\] _0571_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0939_ _0484_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1424__A _0438_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1198__A0 xfer.dout_data\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1207_ _0500_ _0456_ _0666_ _0667_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_49_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1138_ _0628_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1069_ buffer\[19\] xfer.dout_data\[3\] _0573_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0977__B net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0993__A _0503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_840 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_867 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1687_ clknet_4_0_0_clk _0136_ VGND VGND VPWR VPWR xfer.count\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1618__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_935 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1149__A _0634_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1610_ clknet_4_3_0_clk _0080_ VGND VGND VPWR VPWR xfer.din_data\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1541_ _0726_ _0432_ _0309_ _0636_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__a31o_1
X_1472_ rd_addr\[7\] _0256_ _0629_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0927__S _0459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1739_ net71 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1241__B _0522_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1590__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0972_ rd_addr\[4\] net19 VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1524_ _0624_ _0296_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1455_ net19 _0242_ _0237_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1386_ xfer.dout_data\[5\] _0592_ _0193_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_52_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1342__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1061__B _0491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_162_Left_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1252__A _0686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1240__A2 _0686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1528__A0 rd_addr\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1240_ _0670_ _0686_ _0693_ _0674_ xfer.din_data\[3\] VGND VGND VPWR VPWR _0083_
+ sky130_fd_sc_hd__o32a_1
XANTENNA__0985__B _0522_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1171_ _0647_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1101__S _0571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0955_ _0427_ _0433_ config_cont _0435_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__a211o_2
XFILLER_0_55_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0886_ _0316_ _0382_ _0429_ _0431_ _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput101 net101 VGND VGND VPWR VPWR rdata[28] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1519__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput112 net112 VGND VGND VPWR VPWR rdata[9] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1507_ _0283_ rd_addr\[15\] _0249_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1438_ xfer.flash_csb _0478_ _0457_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__a21o_1
X_1369_ _0542_ net50 xfer.dout_data\[2\] _0536_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput14 addr[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput25 cfgreg_di[0] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 cfgreg_di[2] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput47 flash_io0_di VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_149_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1223_ net1 _0675_ _0678_ _0679_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__a211o_1
XFILLER_0_165_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1154_ _0638_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1085_ xfer.din_data\[2\] _0586_ _0456_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0938_ _0436_ _0483_ _0479_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__and3b_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0869_ _0409_ _0410_ _0413_ _0414_ _0415_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__o2111a_1
XANTENNA__0963__B2 state\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1651__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1530__A _0232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1424__B _0478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1674__CLK clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1370__A1 xfer.dout_data\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1206_ state\[3\] state\[9\] _0665_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_4_7_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1137_ net106 buffer\[3\] _0624_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1068_ _0576_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1547__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1697__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1040__A0 xfer.dout_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1686_ clknet_4_1_0_clk _0135_ VGND VGND VPWR VPWR xfer.dummy_count\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1345__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0854__B1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1098__B1 _0535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1540_ rd_addr\[23\] _0382_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1471_ _0726_ _0253_ _0254_ _0255_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1712__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1738_ net50 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1669_ clknet_4_4_0_clk _0121_ VGND VGND VPWR VPWR xfer.fetch sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_595 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0827__B1 rd_addr\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1241__C _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_93_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_15_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0971_ _0345_ _0506_ _0508_ _0509_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1243__B1 _0686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1523_ rd_addr\[18\] rd_addr\[19\] _0373_ _0232_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1454_ _0404_ _0405_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1385_ _0542_ xfer.dout_data\[3\] xfer.dout_data\[6\] _0535_ VGND VGND VPWR VPWR
+ _0193_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1608__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_758 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ buffer\[17\] net89 _0645_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0954_ state\[10\] _0491_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0885_ rd_addr\[23\] _0382_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__nand2_1
XANTENNA__1231__A3 _0686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput102 net102 VGND VGND VPWR VPWR rdata[29] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput113 net113 VGND VGND VPWR VPWR ready sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1506_ rd_addr\[15\] _0392_ _0282_ _0237_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1437_ _0448_ _0609_ _0669_ _0230_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__o211a_1
X_1368_ _0180_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1299_ _0361_ _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_69_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1455__A0 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1580__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_896 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_963 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput15 addr[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
XFILLER_0_107_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput37 cfgreg_di[31] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput26 cfgreg_di[10] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput48 flash_io1_di VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_133_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1222_ _0487_ _0455_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__and2_1
X_1153_ buffer\[9\] net112 _0636_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__mux2_1
X_1084_ xfer.obuffer\[1\] _0535_ _0585_ xfer.obuffer\[0\] VGND VGND VPWR VPWR _0586_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1437__B1 _0669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0937_ _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_3_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1348__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0868_ _0318_ _0376_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__xnor2_1
XANTENNA__0963__A2 _0437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0799_ rd_addr\[5\] net20 VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__xor2_2
XFILLER_0_61_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1083__A _0541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1370__A2 _0592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1205_ _0665_ _0524_ _0519_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1136_ _0627_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1122__A2 _0541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1067_ buffer\[18\] xfer.dout_data\[2\] _0573_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_945 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_113_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1104__A2 _0592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1641__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1685_ clknet_4_1_0_clk _0134_ VGND VGND VPWR VPWR xfer.dummy_count\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1119_ xfer.xfer_ddr _0542_ _0472_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__and3_1
XFILLER_0_165_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1098__A1 _0541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1664__CLK clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_11_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1270__A1 xfer.dout_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1470_ _0232_ net22 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output76_A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1261__A1 _0438_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1737_ net49 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
XANTENNA__1356__A _0438_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1668_ clknet_4_4_0_clk xfer.xfer_ddr VGND VGND VPWR VPWR xfer.xfer_ddr_q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1599_ clknet_4_15_0_clk _0069_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1687__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1030__S config_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_125_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0990__D _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0970_ rd_addr\[3\] _0336_ _0338_ net14 _0325_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1243__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1522_ _0500_ _0387_ _0725_ rd_addr\[19\] VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1453_ _0241_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1384_ _0192_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1025__S config_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1225__A1 config_qspi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1702__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0953_ _0495_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0884_ _0349_ _0430_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput103 net103 VGND VGND VPWR VPWR rdata[2] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1505_ _0395_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1436_ xfer.flash_csb _0609_ _0448_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__o21ai_1
X_1367_ _0179_ xfer.dout_data\[2\] _0174_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1298_ config_en net37 net46 VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput16 addr[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
XFILLER_0_108_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput27 cfgreg_di[11] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput49 flash_io2_di VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_8
Xinput38 cfgreg_di[3] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_133_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1221_ _0676_ _0677_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__or2_1
X_1152_ _0637_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1083_ _0541_ _0534_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__nor2_4
XANTENNA__1437__A1 _0448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0936_ _0438_ _0454_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0867_ _0336_ _0412_ _0347_ _0411_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_3_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0798_ _0331_ _0335_ _0341_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__or4b_1
XFILLER_0_3_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1373__B1 xfer.dout_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1083__B _0534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1419_ _0451_ _0450_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_818 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_159_Left_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1539__A _0232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0800__B net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1570__CLK clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1204_ state\[0\] state\[1\] _0663_ _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__or4_1
X_1135_ net103 buffer\[2\] _0624_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1066_ _0575_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1359__A _0438_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0919_ xfer.xfer_ddr VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__clkinv_2
XFILLER_0_141_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_637 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1593__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1296__3 clknet_4_0_0_clk VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__inv_2
XFILLER_0_53_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_870 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1684_ clknet_4_4_0_clk _0133_ VGND VGND VPWR VPWR xfer.dummy_count\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1118_ _0466_ _0611_ _0613_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1049_ _0564_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1246__C1 state\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_584 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1261__A2 _0487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1736_ net48 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1667_ clknet_4_5_0_clk _0120_ VGND VGND VPWR VPWR softreset sky130_fd_sc_hd__dfxtp_1
X_1598_ clknet_4_15_0_clk _0068_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1237__C1 state\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1311__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1631__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1521_ _0294_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1452_ rd_addr\[3\] _0240_ _0629_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1383_ _0191_ xfer.dout_data\[6\] _0174_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0809__A2 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1131__S _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1219__C1 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1719_ clknet_4_9_0_clk _0168_ VGND VGND VPWR VPWR rd_addr\[23\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__1654__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_140_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1225__A2 _0522_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1161__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1740__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0952_ _0437_ _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1677__CLK clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0883_ rd_addr\[21\] _0375_ _0373_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput104 net104 VGND VGND VPWR VPWR rdata[30] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1504_ _0281_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1435_ _0229_ din_ddr _0526_ _0669_ xfer.xfer_dspi VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__a32o_1
X_1366_ xfer.dout_data\[0\] _0592_ _0178_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1353__C net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 addr[2] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_0_91_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput28 cfgreg_di[16] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput39 cfgreg_di[4] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1735__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1382__A1 xfer.dout_data\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1220_ net8 _0503_ _0528_ net23 VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1151_ buffer\[8\] net111 _0636_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__mux2_1
XANTENNA__1470__A _0232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1082_ _0584_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0814__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0935_ _0480_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0866_ _0347_ _0411_ _0412_ _0336_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__0948__B2 state\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0797_ _0342_ _0343_ _0344_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1373__A1 _0542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1373__B2 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1418_ _0451_ _0217_ _0611_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1125__A1 _0438_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1349_ _0763_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1539__B net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1052__A0 xfer.dout_data\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1465__A _0726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1715__CLK clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1203_ state\[8\] state\[12\] state\[11\] VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1134_ _0626_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_49_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1065_ buffer\[17\] xfer.dout_data\[1\] _0573_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0918_ xfer.xfer_dspi _0449_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__nand2_2
XFILLER_0_141_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0849_ _0358_ _0395_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1314__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_162_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_693 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_838 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1025__A0 config_do\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1683_ clknet_4_4_0_clk _0132_ VGND VGND VPWR VPWR xfer.dummy_count\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1117_ _0592_ _0612_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__nand2_1
X_1048_ xfer.dout_data\[4\] buffer\[12\] _0559_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1044__S _0559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1560__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1743__A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1261__A3 _0454_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0822__A rd_addr\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1735_ net47 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1666_ clknet_4_7_0_clk _0003_ VGND VGND VPWR VPWR state\[12\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_57_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1597_ clknet_4_15_0_clk _0067_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_53_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0827__A3 _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_700 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1583__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1502__S _0237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1476__A0 rd_addr\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_703 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0987__C1 _0487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1738__A net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1520_ rd_addr\[18\] _0293_ _0267_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1451_ net18 _0412_ _0237_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux2_1
X_1382_ xfer.dout_data\[4\] _0592_ _0190_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_52_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1219__B1 state\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1718_ clknet_4_10_0_clk _0167_ VGND VGND VPWR VPWR rd_addr\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1649_ clknet_4_5_0_clk _0115_ VGND VGND VPWR VPWR config_clk sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_703 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0951_ state\[11\] _0483_ _0493_ state\[3\] VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0882_ _0355_ _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput105 net105 VGND VGND VPWR VPWR rdata[31] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1503_ rd_addr\[14\] _0280_ _0267_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1434_ xfer.din_qspi VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1365_ _0542_ net49 xfer.dout_data\[1\] _0536_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1142__S _0629_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1621__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_706 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1317__S net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1052__S _0559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput18 addr[3] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
XFILLER_0_65_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput29 cfgreg_di[17] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1382__A2 _0592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1150_ _0635_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1470__B net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1081_ _0583_ xfer.obuffer\[1\] _0571_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1644__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0934_ _0436_ _0478_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__and3b_1
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0865_ rd_addr\[2\] rd_addr\[3\] VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0948__A2 _0437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0830__A rd_addr\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0796_ rd_addr\[1\] net12 VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1373__A2 xfer.dout_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1137__S _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1417_ _0459_ _0470_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1348_ net51 _0762_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__and2_1
X_1279_ _0720_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1667__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0915__A _0459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1746__A config_qspi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1465__B net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1202_ state\[5\] state\[2\] state\[4\] state\[6\] VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1133_ net92 buffer\[1\] _0624_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1064_ _0574_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_66_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0825__A _0333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1291__A1 _0726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0917_ _0448_ xfer.count\[1\] _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0848_ _0333_ _0365_ _0371_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0779_ _0325_ _0326_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1391__A _0459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1282__A1 xfer.dout_data\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1682_ clknet_4_4_0_clk _0131_ VGND VGND VPWR VPWR xfer.xfer_qspi sky130_fd_sc_hd__dfxtp_2
XFILLER_0_151_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1116_ _0451_ xfer.count\[1\] _0461_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1047_ _0563_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1264__A1 _0522_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1255__B2 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1255__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1705__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1494__A1 _0232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1246__A1 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_759 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1665_ clknet_4_6_0_clk _0002_ VGND VGND VPWR VPWR state\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1596_ clknet_4_14_0_clk _0066_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_931 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1237__A1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1237__B2 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1228__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_759 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1450_ _0239_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
X_1381_ _0542_ xfer.dout_data\[2\] xfer.dout_data\[5\] _0535_ VGND VGND VPWR VPWR
+ _0190_ sky130_fd_sc_hd__a22o_1
XANTENNA_output74_A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1219__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0833__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1717_ clknet_4_10_0_clk _0166_ VGND VGND VPWR VPWR rd_addr\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1648_ clknet_4_5_0_clk _0114_ VGND VGND VPWR VPWR config_csb sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1579_ clknet_4_13_0_clk _0049_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1550__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0969__B1 rd_addr\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_637 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0950_ _0455_ _0492_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0881_ _0338_ _0379_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1385__B1 xfer.dout_data\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput106 net106 VGND VGND VPWR VPWR rdata[3] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1502_ net6 _0279_ _0237_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__mux2_1
XANTENNA__1573__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1433_ xfer.din_qspi din_ddr _0526_ _0669_ xfer.xfer_ddr VGND VGND VPWR VPWR _0141_
+ sky130_fd_sc_hd__a32o_1
X_1364_ _0177_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_129_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput19 addr[4] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1596__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1080_ xfer.din_data\[1\] _0456_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0933_ _0361_ softreset VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__nor2_4
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0864_ rd_addr\[2\] rd_addr\[3\] rd_addr\[4\] VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__nand3_1
XFILLER_0_71_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0948__A3 _0491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0795_ rd_addr\[0\] net1 VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1358__B1 _0448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1416_ _0216_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
X_1347_ config_do\[2\] net36 net43 VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__mux2_1
XANTENNA__1153__S _0636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1278_ buffer\[4\] xfer.dout_data\[4\] _0715_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_137_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1063__S _0573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_146_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_155_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1201_ _0662_ _0502_ _0496_ _0437_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__o211a_1
XANTENNA__1611__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1132_ _0625_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1063_ buffer\[16\] xfer.dout_data\[0\] _0573_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_164_Left_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0841__A _0333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0916_ xfer.count\[1\] _0461_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0847_ _0315_ _0387_ _0389_ _0391_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0778_ rd_addr\[17\] net9 VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0798__D_N _0345_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_868 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1681_ clknet_4_4_0_clk _0130_ VGND VGND VPWR VPWR xfer.xfer_rd sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1492__A _0232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0836__A _0333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1115_ _0451_ _0610_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1046_ xfer.dout_data\[3\] buffer\[11\] _0559_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1657__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1255__A2 _0503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1516__S _0267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1479__C1 _0726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1494__A2 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1664_ clknet_4_7_0_clk _0001_ VGND VGND VPWR VPWR state\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1595_ clknet_4_15_0_clk _0065_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1182__A1 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1161__S _0636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1029_ xfer.flash_io2_do xfer_io2_90 _0522_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1071__S _0573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1228__A2 _0487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1380_ _0189_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1467__A2 _0249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1219__A2 _0487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1716_ clknet_4_9_0_clk _0165_ VGND VGND VPWR VPWR rd_addr\[20\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1647_ clknet_4_5_0_clk _0113_ VGND VGND VPWR VPWR config_oe\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1155__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1578_ clknet_4_13_0_clk _0048_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0969__A1 rd_addr\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0880_ _0380_ _0381_ _0386_ _0394_ _0426_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__o2111a_2
XFILLER_0_103_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1385__A1 _0542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput107 net107 VGND VGND VPWR VPWR rdata[4] sky130_fd_sc_hd__clkbuf_1
XANTENNA__1718__CLK clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1385__B2 _0535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1501_ _0392_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1432_ xfer.din_tag\[2\] _0500_ _0226_ _0671_ _0524_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_71_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1363_ _0176_ xfer.dout_data\[1\] _0174_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1005__A config_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0811__B1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1367__A1 xfer.dout_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0932_ _0439_ _0457_ _0446_ _0477_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__or4_4
XFILLER_0_43_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0863_ rd_addr\[6\] _0376_ _0320_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_858 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0794_ rd_addr\[0\] net1 VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1690__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1415_ _0438_ _0478_ _0215_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__and3_1
X_1346_ _0761_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
X_1277_ _0719_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_84_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1046__A0 xfer.dout_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1563__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1519__S rd_inc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1200_ state\[7\] VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1131_ net81 buffer\[0\] _0624_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1062_ _0572_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1291__A3 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0915_ _0459_ _0460_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_836 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0846_ _0323_ _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0777_ net9 rd_addr\[17\] VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__or2b_1
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1329_ config_oe\[2\] net26 net44 VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__mux2_1
XANTENNA__1586__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1680_ clknet_4_12_0_clk xfer.xfer_tag\[2\] VGND VGND VPWR VPWR xfer.dout_tag\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1114_ _0459_ _0470_ _0458_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__and3_1
XANTENNA__1249__B1 _0698_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_152_10 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1045_ _0562_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0852__A rd_addr\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1159__S _0636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0829_ _0366_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_23_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1601__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1069__S _0573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1532__S _0267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1663_ clknet_4_6_0_clk _0012_ VGND VGND VPWR VPWR state\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1594_ clknet_4_15_0_clk _0064_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1442__S _0233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_861 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1028_ _0551_ VGND VGND VPWR VPWR xfer.flash_io2_do sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1624__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1228__A3 _0483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_780 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1647__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1498__A _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1715_ clknet_4_9_0_clk _0164_ VGND VGND VPWR VPWR rd_addr\[19\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_53_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1646_ clknet_4_5_0_clk _0112_ VGND VGND VPWR VPWR config_oe\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1577_ clknet_4_13_0_clk _0047_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1172__S _0645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0803__D_N _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0934__B _0478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0950__A _0455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1385__A2 xfer.dout_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput108 net108 VGND VGND VPWR VPWR rdata[5] sky130_fd_sc_hd__clkbuf_1
X_1500_ rd_addr\[14\] _0378_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1431_ state\[5\] state\[11\] _0226_ _0228_ _0500_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__o311a_1
XFILLER_0_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput90 net90 VGND VGND VPWR VPWR rdata[18] sky130_fd_sc_hd__clkbuf_1
X_1362_ net48 xfer.dout_data\[0\] _0536_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__mux2_1
XANTENNA__0828__C rd_addr\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1293_ _0726_ _0624_ _0728_ _0363_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1021__A _0547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1073__A1 xfer.dout_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0860__A net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_948 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1629_ clknet_4_9_0_clk _0099_ VGND VGND VPWR VPWR rd_valid sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0787__A1_N rd_addr\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1077__S _0573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_150_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ _0458_ _0468_ _0476_ _0440_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0862_ rd_addr\[6\] _0320_ _0376_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0793_ rd_addr\[3\] _0336_ _0339_ _0340_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0830__D _0333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1414_ _0210_ _0213_ _0569_ _0214_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_48_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1345_ net51 _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1276_ buffer\[3\] xfer.dout_data\[3\] _0715_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1506__C1 _0237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1360__S _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1708__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1130_ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_69_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1061_ xfer.dout_tag\[0\] _0491_ _0558_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1276__A1 xfer.dout_data\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0914_ xfer.count\[0\] xfer.count\[2\] xfer.count\[1\] xfer.count\[3\] VGND VGND
+ VPWR VPWR _0460_ sky130_fd_sc_hd__or4_2
XFILLER_0_28_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0845_ _0333_ rd_addr\[14\] _0371_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__and3_1
XANTENNA__0787__B1 _0333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0776_ net17 rd_addr\[2\] VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__xor2_2
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_87_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1328_ _0749_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__1180__S _0645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1259_ _0500_ _0497_ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_96_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1090__S _0571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1258__A1 config_qspi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1680__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0805__A_N rd_addr\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1194__A0 xfer.dout_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1113_ _0446_ _0460_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__nor2_1
X_1044_ xfer.dout_data\[2\] buffer\[10\] _0559_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1013__B config_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0852__B _0366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0828_ rd_addr\[18\] rd_addr\[19\] rd_addr\[20\] VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1553__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1412__A1 _0459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1085__S _0456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1114__A _0459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1576__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1662_ clknet_4_7_0_clk _0011_ VGND VGND VPWR VPWR state\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1593_ clknet_4_15_0_clk _0063_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1027_ _0541_ xfer.obuffer\[6\] _0533_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__and3_1
XFILLER_0_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_164_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1294__1_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1599__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1397__B1 _0483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1714_ clknet_4_12_0_clk _0163_ VGND VGND VPWR VPWR rd_addr\[18\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_81_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1645_ clknet_4_5_0_clk _0111_ VGND VGND VPWR VPWR config_oe\[1\] sky130_fd_sc_hd__dfxtp_1
X_1576_ clknet_4_12_0_clk _0046_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1363__S _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0934__C _0479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput109 net109 VGND VGND VPWR VPWR rdata[6] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1430_ xfer.din_tag\[1\] _0226_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__or2b_1
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output72_A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1361_ _0175_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1614__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput91 net91 VGND VGND VPWR VPWR rdata[19] sky130_fd_sc_hd__clkbuf_1
Xoutput80 net80 VGND VGND VPWR VPWR flash_io3_oe sky130_fd_sc_hd__clkbuf_1
X_1292_ _0499_ _0436_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_50_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1058__C1 _0459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1448__S _0237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1628_ clknet_4_11_0_clk _0098_ VGND VGND VPWR VPWR buffer\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1559_ clknet_4_14_0_clk _0029_ VGND VGND VPWR VPWR buffer\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0811__A2 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0770__B net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1637__CLK clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_107_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0930_ _0469_ _0473_ _0475_ _0450_ xfer.count\[3\] VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__o32a_1
XFILLER_0_166_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0861_ _0324_ _0345_ _0406_ _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__and4_1
XFILLER_0_83_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0792_ net23 rd_addr\[8\] VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1515__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1413_ _0462_ _0585_ _0610_ _0535_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a22o_1
X_1344_ config_do\[1\] net32 net43 VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__mux2_1
X_1275_ _0718_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1032__A _0541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0871__A rd_addr\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1178__S _0645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1207__A _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_919 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1117__A _0592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ xfer.din_data\[0\] _0526_ _0571_ xfer.obuffer\[0\] VGND VGND VPWR VPWR _0025_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0913_ xfer.flash_clk VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__buf_4
XFILLER_0_28_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_133_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0844_ _0350_ _0390_ _0373_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0775_ rd_addr\[15\] net7 VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__xor2_2
XFILLER_0_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1027__A _0541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1461__S _0629_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1327_ _0731_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__and2_1
X_1258_ xfer.din_qspi config_qspi _0530_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__mux2_1
X_1189_ _0656_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_166_Right_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1371__S _0174_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0776__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1112_ _0608_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1043_ _0561_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1013__C _0533_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1421__A2 _0541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0827_ rd_addr\[18\] rd_addr\[19\] _0373_ rd_addr\[20\] VGND VGND VPWR VPWR _0374_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1456__S _0629_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0999__A1 _0459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_164_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_941 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_840 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1412__A2 _0535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_14 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1661_ clknet_4_6_0_clk _0010_ VGND VGND VPWR VPWR state\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1592_ clknet_4_14_0_clk _0062_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1026_ _0550_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_146_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1186__S _0645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1670__CLK clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0905__A1 _0448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1215__A _0487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0773__B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_927 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1096__S _0571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_693 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_774 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1713_ clknet_4_8_0_clk _0162_ VGND VGND VPWR VPWR rd_addr\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1693__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1644_ clknet_4_5_0_clk _0110_ VGND VGND VPWR VPWR config_oe\[0\] sky130_fd_sc_hd__dfxtp_1
X_1575_ clknet_4_13_0_clk _0045_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_619 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ config_en _0533_ _0536_ _0540_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__a31o_4
XFILLER_0_92_836 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1379__A1 xfer.dout_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_777 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0768__B net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0784__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1566__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1360_ _0172_ xfer.dout_data\[0\] _0174_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput70 net70 VGND VGND VPWR VPWR cfgreg_do[9] sky130_fd_sc_hd__clkbuf_1
Xoutput92 net92 VGND VGND VPWR VPWR rdata[1] sky130_fd_sc_hd__clkbuf_1
Xoutput81 net81 VGND VGND VPWR VPWR rdata[0] sky130_fd_sc_hd__clkbuf_1
XANTENNA_output65_A net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1291_ _0726_ _0434_ _0624_ _0727_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__a31o_1
XFILLER_0_156_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1627_ clknet_4_13_0_clk _0097_ VGND VGND VPWR VPWR buffer\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1558_ clknet_4_15_0_clk _0028_ VGND VGND VPWR VPWR buffer\[18\] sky130_fd_sc_hd__dfxtp_1
X_1489_ net3 _0269_ _0237_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__mux2_1
XANTENNA__1589__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_746 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1288__B1 _0437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0860_ net19 _0404_ _0405_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0791_ _0337_ net18 _0338_ net14 VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1212__B1 _0669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1412_ _0459_ _0535_ _0569_ _0212_ _0449_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_139_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1343_ _0759_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
X_1274_ buffer\[2\] xfer.dout_data\[2\] _0715_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0871__B _0366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1451__A0 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ _0483_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1207__B _0456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1604__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0912_ _0451_ xfer.count\[3\] VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__or2_2
XANTENNA__1433__B1 _0669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0843_ rd_addr\[18\] _0315_ _0350_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0774_ _0318_ _0319_ _0320_ _0321_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1326_ config_oe\[1\] net42 net44 VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__mux2_1
X_1257_ xfer.din_data\[7\] _0674_ _0698_ _0706_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__o22a_1
X_1188_ xfer.dout_data\[2\] net99 _0635_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__mux2_1
XANTENNA__1627__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1111_ _0607_ xfer.obuffer\[7\] _0571_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__mux2_1
X_1042_ xfer.dout_data\[1\] buffer\[9\] _0559_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1013__D _0542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1406__B1 _0478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0826_ _0372_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_6_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0877__A _0321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1472__S _0629_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1309_ _0731_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_127_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_152_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_26 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_161_Left_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_945 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1660_ clknet_4_6_0_clk _0009_ VGND VGND VPWR VPWR state\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1591_ clknet_4_15_0_clk _0061_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1025_ config_do\[1\] _0549_ config_en VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__mux2_2
XFILLER_0_159_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_750 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0809_ _0352_ net19 _0353_ _0356_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1712_ clknet_4_8_0_clk _0161_ VGND VGND VPWR VPWR rd_addr\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_786 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1643_ clknet_4_7_0_clk _0109_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1574_ clknet_4_13_0_clk _0044_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1008_ config_oe\[0\] _0537_ _0539_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_146_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0890__A _0363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1067__A1 xfer.dout_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_14_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0959__B _0456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput60 net60 VGND VGND VPWR VPWR cfgreg_do[1] sky130_fd_sc_hd__clkbuf_1
Xoutput71 net71 VGND VGND VPWR VPWR flash_clk sky130_fd_sc_hd__clkbuf_1
Xoutput93 net93 VGND VGND VPWR VPWR rdata[20] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput82 net82 VGND VGND VPWR VPWR rdata[10] sky130_fd_sc_hd__clkbuf_1
XANTENNA__1542__A2 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1290_ _0434_ _0363_ _0636_ rd_wait VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__o211a_1
XANTENNA_output58_A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0975__A rd_addr\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1660__CLK clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1626_ clknet_4_12_0_clk _0096_ VGND VGND VPWR VPWR buffer\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1557_ clknet_4_15_0_clk _0027_ VGND VGND VPWR VPWR buffer\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1488_ rd_addr\[11\] _0419_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1480__S _0249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_758 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1683__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1460__A1 _0726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0790_ rd_addr\[21\] VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1411_ _0211_ _0459_ _0466_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1342_ net51 _0758_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__and2_1
X_1273_ _0717_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1032__C _0533_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0988_ state\[8\] _0481_ _0485_ _0525_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1556__CLK clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1609_ clknet_4_6_0_clk _0079_ VGND VGND VPWR VPWR xfer.xfer_tag\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0972__B net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0911_ xfer.resetn VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1579__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0842_ _0334_ _0388_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0773_ rd_addr\[9\] net24 VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__xor2_4
XFILLER_0_4_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1027__C _0533_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1325_ _0747_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__1324__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1256_ net22 state\[12\] _0456_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__a31o_1
X_1187_ _0655_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_56_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_2_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1188__A0 xfer.dout_data\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1218__B _0455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_74_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0792__B rd_addr\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1409__A xfer.count\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1110_ xfer.din_data\[7\] _0456_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ _0560_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__1103__B1 _0535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0825_ _0333_ _0364_ _0365_ _0371_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__and4_1
XFILLER_0_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_670 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1038__B _0479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1308_ config_cont net33 net45 VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1239_ net59 _0487_ _0483_ _0692_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1229__A config_cont VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_754 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1590_ clknet_4_15_0_clk _0060_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1617__CLK clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1024_ xfer.flash_io1_do xfer_io1_90 _0522_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0808_ _0354_ net5 rd_addr\[21\] _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1094__A2 _0592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_959 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_10_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1711_ clknet_4_8_0_clk _0160_ VGND VGND VPWR VPWR rd_addr\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_584 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1642_ clknet_4_7_0_clk _0108_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1573_ clknet_4_13_0_clk _0043_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1007_ xfer.xfer_rd _0537_ _0538_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0890__B _0436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1536__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0959__C _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1417__A _0459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput61 net61 VGND VGND VPWR VPWR cfgreg_do[20] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput72 net72 VGND VGND VPWR VPWR flash_csb sky130_fd_sc_hd__clkbuf_1
Xoutput94 net94 VGND VGND VPWR VPWR rdata[21] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput83 net83 VGND VGND VPWR VPWR rdata[11] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1298__S net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1230__A2 _0487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1625_ clknet_4_13_0_clk _0095_ VGND VGND VPWR VPWR buffer\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1327__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1556_ clknet_4_15_0_clk _0026_ VGND VGND VPWR VPWR buffer\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1487_ _0268_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1403__C _0483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1460__A2 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0778__B_N net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1212__A2 _0526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1410_ xfer.count\[0\] VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1341_ config_do\[0\] net25 net43 VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__mux2_1
X_1272_ buffer\[1\] xfer.dout_data\[1\] _0715_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_103_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ state\[12\] _0523_ _0524_ _0487_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1608_ clknet_4_3_0_clk _0078_ VGND VGND VPWR VPWR xfer.xfer_tag\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1539_ _0232_ net16 VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_874 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1650__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0910_ state\[0\] _0437_ _0456_ _0363_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_32_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0841_ _0333_ _0371_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0772_ rd_addr\[7\] net22 VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__xor2_2
XFILLER_0_4_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1324_ _0731_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__and2_1
X_1255_ net16 _0503_ _0528_ net7 VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1186_ xfer.dout_data\[1\] net98 _0645_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1486__S _0267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1673__CLK clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1360__A1 xfer.dout_data\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1040_ xfer.dout_data\[0\] buffer\[8\] _0559_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1103__A1 _0541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1696__CLK clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0824_ _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0917__A1 _0448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1307_ _0735_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_127_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1238_ net11 _0503_ _0675_ net18 _0691_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__a221o_1
XANTENNA__0893__B xfer.count\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1169_ _0646_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0853__B1 rd_addr\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1030__A0 config_do\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1569__CLK clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0844__A0 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_730 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0978__B _0321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1088__B1 _0585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1023_ _0449_ xfer.obuffer\[5\] _0464_ xfer.obuffer\[7\] _0548_ VGND VGND VPWR VPWR
+ xfer.flash_io1_do sky130_fd_sc_hd__o221a_1
XFILLER_0_163_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0807_ net14 VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0888__B net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1711__CLK clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_662 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1710_ clknet_4_8_0_clk _0159_ VGND VGND VPWR VPWR rd_addr\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0989__A _0483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1641_ clknet_4_5_0_clk _0107_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_950 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1572_ clknet_4_4_0_clk _0042_ VGND VGND VPWR VPWR xfer.last_fetch sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1006_ _0446_ _0445_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1607__CLK clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_149_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1527__A1 _0232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0959__D _0500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput84 net84 VGND VGND VPWR VPWR rdata[12] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput73 net73 VGND VGND VPWR VPWR flash_io0_do sky130_fd_sc_hd__clkbuf_1
Xoutput62 net62 VGND VGND VPWR VPWR cfgreg_do[21] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_158_Left_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput95 net95 VGND VGND VPWR VPWR rdata[22] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_746 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0974__C1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1230__A3 _0455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1624_ clknet_4_12_0_clk _0094_ VGND VGND VPWR VPWR buffer\[3\] sky130_fd_sc_hd__dfxtp_1
X_1294__1 clknet_4_0_0_clk VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__inv_2
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1555_ clknet_4_3_0_clk _0025_ VGND VGND VPWR VPWR xfer.obuffer\[0\] sky130_fd_sc_hd__dfxtp_1
X_1486_ rd_addr\[10\] _0266_ _0267_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1489__S _0237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1340_ _0757_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1271_ _0716_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1436__B1 _0448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ _0492_ state\[3\] VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1607_ clknet_4_12_0_clk _0077_ VGND VGND VPWR VPWR xfer.xfer_tag\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1538_ _0307_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__0896__B xfer.count\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1469_ rd_addr\[6\] _0376_ rd_addr\[7\] VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_923 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1433__A3 _0526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0840_ rd_addr\[18\] _0373_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0771_ rd_addr\[11\] net3 VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__xor2_2
XFILLER_0_3_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_730 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_774 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1323_ config_oe\[0\] net41 net44 VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1254_ _0704_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1185_ _0654_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_866 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0969_ rd_addr\[10\] _0507_ rd_addr\[20\] _0332_ _0326_ VGND VGND VPWR VPWR _0508_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_691 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_858 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1406__A3 _0483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0823_ _0366_ _0367_ _0368_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__and4_1
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_691 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0917__A2 xfer.count\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1306_ _0731_ _0734_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_4_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1237_ net3 _0528_ _0486_ _0499_ state\[4\] VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1351__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1168_ buffer\[16\] net88 _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1099_ xfer.obuffer\[3\] _0592_ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1497__S _0726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1640__CLK clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_582 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_700 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1526__A rd_inc VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0994__B _0519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1022_ _0538_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1663__CLK clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__0938__A_N _0436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0806_ rd_addr\[13\] VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_146_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_674 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1251__A1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1020__S config_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_161_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1251__B2 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1686__CLK clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1242__B2 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1242__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1640_ clknet_4_5_0_clk _0106_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1571_ clknet_4_4_0_clk _0041_ VGND VGND VPWR VPWR xfer.count\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_158_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1105__S _0455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1005_ config_en VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__clkinv_2
XFILLER_0_159_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1481__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1233__A1 config_qspi VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1233__B2 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1559__CLK clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_892 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_636 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1527__A2 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput85 net85 VGND VGND VPWR VPWR rdata[13] sky130_fd_sc_hd__clkbuf_1
Xoutput63 net63 VGND VGND VPWR VPWR cfgreg_do[22] sky130_fd_sc_hd__clkbuf_1
Xoutput74 net74 VGND VGND VPWR VPWR flash_io0_oe sky130_fd_sc_hd__clkbuf_1
Xoutput96 net96 VGND VGND VPWR VPWR rdata[23] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0783__A_N net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_758 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_870 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1701__CLK clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1623_ clknet_4_12_0_clk _0093_ VGND VGND VPWR VPWR buffer\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1554_ clknet_4_11_0_clk _0024_ VGND VGND VPWR VPWR buffer\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1485_ _0623_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__buf_4
.ends

