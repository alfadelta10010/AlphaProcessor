magic
tech sky130A
magscale 1 2
timestamp 1701598694
<< obsli1 >>
rect 1104 2159 91908 93041
<< obsm1 >>
rect 934 2048 92078 93072
<< metal2 >>
rect 23202 0 23258 800
rect 69754 0 69810 800
<< obsm2 >>
rect 938 856 92074 93061
rect 938 800 23146 856
rect 23314 800 69698 856
rect 69866 800 92074 856
<< metal3 >>
rect 0 91672 800 91792
rect 0 84872 800 84992
rect 92303 81336 93103 81456
rect 92303 80792 93103 80912
rect 92303 80248 93103 80368
rect 92303 79704 93103 79824
rect 92303 79160 93103 79280
rect 92303 78616 93103 78736
rect 0 78072 800 78192
rect 92303 78072 93103 78192
rect 92303 77528 93103 77648
rect 92303 76984 93103 77104
rect 92303 76440 93103 76560
rect 92303 75896 93103 76016
rect 92303 75352 93103 75472
rect 92303 74808 93103 74928
rect 92303 74264 93103 74384
rect 92303 73720 93103 73840
rect 92303 73176 93103 73296
rect 92303 72632 93103 72752
rect 92303 72088 93103 72208
rect 92303 71544 93103 71664
rect 0 71272 800 71392
rect 92303 71000 93103 71120
rect 92303 70456 93103 70576
rect 92303 69912 93103 70032
rect 92303 69368 93103 69488
rect 92303 68824 93103 68944
rect 92303 68280 93103 68400
rect 92303 67736 93103 67856
rect 92303 67192 93103 67312
rect 92303 66648 93103 66768
rect 92303 66104 93103 66224
rect 92303 65560 93103 65680
rect 92303 65016 93103 65136
rect 0 64472 800 64592
rect 92303 64472 93103 64592
rect 92303 63928 93103 64048
rect 92303 63384 93103 63504
rect 92303 62840 93103 62960
rect 92303 62296 93103 62416
rect 92303 61752 93103 61872
rect 92303 61208 93103 61328
rect 92303 60664 93103 60784
rect 92303 60120 93103 60240
rect 92303 59576 93103 59696
rect 92303 59032 93103 59152
rect 92303 58488 93103 58608
rect 92303 57944 93103 58064
rect 0 57672 800 57792
rect 92303 57400 93103 57520
rect 92303 56856 93103 56976
rect 92303 56312 93103 56432
rect 92303 55768 93103 55888
rect 92303 55224 93103 55344
rect 92303 54680 93103 54800
rect 92303 54136 93103 54256
rect 92303 53592 93103 53712
rect 92303 53048 93103 53168
rect 92303 52504 93103 52624
rect 92303 51960 93103 52080
rect 92303 51416 93103 51536
rect 0 50872 800 50992
rect 92303 50872 93103 50992
rect 92303 50328 93103 50448
rect 92303 49784 93103 49904
rect 92303 49240 93103 49360
rect 92303 48696 93103 48816
rect 92303 48152 93103 48272
rect 92303 47608 93103 47728
rect 92303 47064 93103 47184
rect 92303 46520 93103 46640
rect 92303 45976 93103 46096
rect 92303 45432 93103 45552
rect 92303 44888 93103 45008
rect 92303 44344 93103 44464
rect 0 44072 800 44192
rect 92303 43800 93103 43920
rect 92303 43256 93103 43376
rect 92303 42712 93103 42832
rect 92303 42168 93103 42288
rect 92303 41624 93103 41744
rect 92303 41080 93103 41200
rect 92303 40536 93103 40656
rect 92303 39992 93103 40112
rect 92303 39448 93103 39568
rect 92303 38904 93103 39024
rect 92303 38360 93103 38480
rect 92303 37816 93103 37936
rect 0 37272 800 37392
rect 92303 37272 93103 37392
rect 92303 36728 93103 36848
rect 92303 36184 93103 36304
rect 92303 35640 93103 35760
rect 92303 35096 93103 35216
rect 92303 34552 93103 34672
rect 92303 34008 93103 34128
rect 92303 33464 93103 33584
rect 92303 32920 93103 33040
rect 92303 32376 93103 32496
rect 92303 31832 93103 31952
rect 92303 31288 93103 31408
rect 92303 30744 93103 30864
rect 0 30472 800 30592
rect 92303 30200 93103 30320
rect 92303 29656 93103 29776
rect 92303 29112 93103 29232
rect 92303 28568 93103 28688
rect 92303 28024 93103 28144
rect 92303 27480 93103 27600
rect 92303 26936 93103 27056
rect 92303 26392 93103 26512
rect 92303 25848 93103 25968
rect 92303 25304 93103 25424
rect 92303 24760 93103 24880
rect 92303 24216 93103 24336
rect 0 23672 800 23792
rect 92303 23672 93103 23792
rect 92303 23128 93103 23248
rect 92303 22584 93103 22704
rect 92303 22040 93103 22160
rect 92303 21496 93103 21616
rect 92303 20952 93103 21072
rect 92303 20408 93103 20528
rect 92303 19864 93103 19984
rect 92303 19320 93103 19440
rect 92303 18776 93103 18896
rect 92303 18232 93103 18352
rect 92303 17688 93103 17808
rect 92303 17144 93103 17264
rect 0 16872 800 16992
rect 92303 16600 93103 16720
rect 92303 16056 93103 16176
rect 92303 15512 93103 15632
rect 92303 14968 93103 15088
rect 92303 14424 93103 14544
rect 92303 13880 93103 14000
rect 92303 13336 93103 13456
rect 0 10072 800 10192
rect 0 3272 800 3392
<< obsm3 >>
rect 798 91872 92303 93057
rect 880 91592 92303 91872
rect 798 85072 92303 91592
rect 880 84792 92303 85072
rect 798 81536 92303 84792
rect 798 81256 92223 81536
rect 798 80992 92303 81256
rect 798 80712 92223 80992
rect 798 80448 92303 80712
rect 798 80168 92223 80448
rect 798 79904 92303 80168
rect 798 79624 92223 79904
rect 798 79360 92303 79624
rect 798 79080 92223 79360
rect 798 78816 92303 79080
rect 798 78536 92223 78816
rect 798 78272 92303 78536
rect 880 77992 92223 78272
rect 798 77728 92303 77992
rect 798 77448 92223 77728
rect 798 77184 92303 77448
rect 798 76904 92223 77184
rect 798 76640 92303 76904
rect 798 76360 92223 76640
rect 798 76096 92303 76360
rect 798 75816 92223 76096
rect 798 75552 92303 75816
rect 798 75272 92223 75552
rect 798 75008 92303 75272
rect 798 74728 92223 75008
rect 798 74464 92303 74728
rect 798 74184 92223 74464
rect 798 73920 92303 74184
rect 798 73640 92223 73920
rect 798 73376 92303 73640
rect 798 73096 92223 73376
rect 798 72832 92303 73096
rect 798 72552 92223 72832
rect 798 72288 92303 72552
rect 798 72008 92223 72288
rect 798 71744 92303 72008
rect 798 71472 92223 71744
rect 880 71464 92223 71472
rect 880 71200 92303 71464
rect 880 71192 92223 71200
rect 798 70920 92223 71192
rect 798 70656 92303 70920
rect 798 70376 92223 70656
rect 798 70112 92303 70376
rect 798 69832 92223 70112
rect 798 69568 92303 69832
rect 798 69288 92223 69568
rect 798 69024 92303 69288
rect 798 68744 92223 69024
rect 798 68480 92303 68744
rect 798 68200 92223 68480
rect 798 67936 92303 68200
rect 798 67656 92223 67936
rect 798 67392 92303 67656
rect 798 67112 92223 67392
rect 798 66848 92303 67112
rect 798 66568 92223 66848
rect 798 66304 92303 66568
rect 798 66024 92223 66304
rect 798 65760 92303 66024
rect 798 65480 92223 65760
rect 798 65216 92303 65480
rect 798 64936 92223 65216
rect 798 64672 92303 64936
rect 880 64392 92223 64672
rect 798 64128 92303 64392
rect 798 63848 92223 64128
rect 798 63584 92303 63848
rect 798 63304 92223 63584
rect 798 63040 92303 63304
rect 798 62760 92223 63040
rect 798 62496 92303 62760
rect 798 62216 92223 62496
rect 798 61952 92303 62216
rect 798 61672 92223 61952
rect 798 61408 92303 61672
rect 798 61128 92223 61408
rect 798 60864 92303 61128
rect 798 60584 92223 60864
rect 798 60320 92303 60584
rect 798 60040 92223 60320
rect 798 59776 92303 60040
rect 798 59496 92223 59776
rect 798 59232 92303 59496
rect 798 58952 92223 59232
rect 798 58688 92303 58952
rect 798 58408 92223 58688
rect 798 58144 92303 58408
rect 798 57872 92223 58144
rect 880 57864 92223 57872
rect 880 57600 92303 57864
rect 880 57592 92223 57600
rect 798 57320 92223 57592
rect 798 57056 92303 57320
rect 798 56776 92223 57056
rect 798 56512 92303 56776
rect 798 56232 92223 56512
rect 798 55968 92303 56232
rect 798 55688 92223 55968
rect 798 55424 92303 55688
rect 798 55144 92223 55424
rect 798 54880 92303 55144
rect 798 54600 92223 54880
rect 798 54336 92303 54600
rect 798 54056 92223 54336
rect 798 53792 92303 54056
rect 798 53512 92223 53792
rect 798 53248 92303 53512
rect 798 52968 92223 53248
rect 798 52704 92303 52968
rect 798 52424 92223 52704
rect 798 52160 92303 52424
rect 798 51880 92223 52160
rect 798 51616 92303 51880
rect 798 51336 92223 51616
rect 798 51072 92303 51336
rect 880 50792 92223 51072
rect 798 50528 92303 50792
rect 798 50248 92223 50528
rect 798 49984 92303 50248
rect 798 49704 92223 49984
rect 798 49440 92303 49704
rect 798 49160 92223 49440
rect 798 48896 92303 49160
rect 798 48616 92223 48896
rect 798 48352 92303 48616
rect 798 48072 92223 48352
rect 798 47808 92303 48072
rect 798 47528 92223 47808
rect 798 47264 92303 47528
rect 798 46984 92223 47264
rect 798 46720 92303 46984
rect 798 46440 92223 46720
rect 798 46176 92303 46440
rect 798 45896 92223 46176
rect 798 45632 92303 45896
rect 798 45352 92223 45632
rect 798 45088 92303 45352
rect 798 44808 92223 45088
rect 798 44544 92303 44808
rect 798 44272 92223 44544
rect 880 44264 92223 44272
rect 880 44000 92303 44264
rect 880 43992 92223 44000
rect 798 43720 92223 43992
rect 798 43456 92303 43720
rect 798 43176 92223 43456
rect 798 42912 92303 43176
rect 798 42632 92223 42912
rect 798 42368 92303 42632
rect 798 42088 92223 42368
rect 798 41824 92303 42088
rect 798 41544 92223 41824
rect 798 41280 92303 41544
rect 798 41000 92223 41280
rect 798 40736 92303 41000
rect 798 40456 92223 40736
rect 798 40192 92303 40456
rect 798 39912 92223 40192
rect 798 39648 92303 39912
rect 798 39368 92223 39648
rect 798 39104 92303 39368
rect 798 38824 92223 39104
rect 798 38560 92303 38824
rect 798 38280 92223 38560
rect 798 38016 92303 38280
rect 798 37736 92223 38016
rect 798 37472 92303 37736
rect 880 37192 92223 37472
rect 798 36928 92303 37192
rect 798 36648 92223 36928
rect 798 36384 92303 36648
rect 798 36104 92223 36384
rect 798 35840 92303 36104
rect 798 35560 92223 35840
rect 798 35296 92303 35560
rect 798 35016 92223 35296
rect 798 34752 92303 35016
rect 798 34472 92223 34752
rect 798 34208 92303 34472
rect 798 33928 92223 34208
rect 798 33664 92303 33928
rect 798 33384 92223 33664
rect 798 33120 92303 33384
rect 798 32840 92223 33120
rect 798 32576 92303 32840
rect 798 32296 92223 32576
rect 798 32032 92303 32296
rect 798 31752 92223 32032
rect 798 31488 92303 31752
rect 798 31208 92223 31488
rect 798 30944 92303 31208
rect 798 30672 92223 30944
rect 880 30664 92223 30672
rect 880 30400 92303 30664
rect 880 30392 92223 30400
rect 798 30120 92223 30392
rect 798 29856 92303 30120
rect 798 29576 92223 29856
rect 798 29312 92303 29576
rect 798 29032 92223 29312
rect 798 28768 92303 29032
rect 798 28488 92223 28768
rect 798 28224 92303 28488
rect 798 27944 92223 28224
rect 798 27680 92303 27944
rect 798 27400 92223 27680
rect 798 27136 92303 27400
rect 798 26856 92223 27136
rect 798 26592 92303 26856
rect 798 26312 92223 26592
rect 798 26048 92303 26312
rect 798 25768 92223 26048
rect 798 25504 92303 25768
rect 798 25224 92223 25504
rect 798 24960 92303 25224
rect 798 24680 92223 24960
rect 798 24416 92303 24680
rect 798 24136 92223 24416
rect 798 23872 92303 24136
rect 880 23592 92223 23872
rect 798 23328 92303 23592
rect 798 23048 92223 23328
rect 798 22784 92303 23048
rect 798 22504 92223 22784
rect 798 22240 92303 22504
rect 798 21960 92223 22240
rect 798 21696 92303 21960
rect 798 21416 92223 21696
rect 798 21152 92303 21416
rect 798 20872 92223 21152
rect 798 20608 92303 20872
rect 798 20328 92223 20608
rect 798 20064 92303 20328
rect 798 19784 92223 20064
rect 798 19520 92303 19784
rect 798 19240 92223 19520
rect 798 18976 92303 19240
rect 798 18696 92223 18976
rect 798 18432 92303 18696
rect 798 18152 92223 18432
rect 798 17888 92303 18152
rect 798 17608 92223 17888
rect 798 17344 92303 17608
rect 798 17072 92223 17344
rect 880 17064 92223 17072
rect 880 16800 92303 17064
rect 880 16792 92223 16800
rect 798 16520 92223 16792
rect 798 16256 92303 16520
rect 798 15976 92223 16256
rect 798 15712 92303 15976
rect 798 15432 92223 15712
rect 798 15168 92303 15432
rect 798 14888 92223 15168
rect 798 14624 92303 14888
rect 798 14344 92223 14624
rect 798 14080 92303 14344
rect 798 13800 92223 14080
rect 798 13536 92303 13800
rect 798 13256 92223 13536
rect 798 10272 92303 13256
rect 880 9992 92303 10272
rect 798 3472 92303 9992
rect 880 3192 92303 3472
rect 798 2143 92303 3192
<< metal4 >>
rect 4208 2128 4528 93072
rect 19568 2128 19888 93072
rect 34928 2128 35248 93072
rect 50288 2128 50608 93072
rect 65648 2128 65968 93072
rect 81008 2128 81328 93072
<< obsm4 >>
rect 63539 17171 65568 69053
rect 66048 17171 66549 69053
<< labels >>
rlabel metal4 s 19568 2128 19888 93072 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 93072 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 93072 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 93072 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 93072 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 93072 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 92303 51416 93103 51536 6 addr[0]
port 3 nsew signal input
rlabel metal3 s 92303 56856 93103 56976 6 addr[10]
port 4 nsew signal input
rlabel metal3 s 92303 57400 93103 57520 6 addr[11]
port 5 nsew signal input
rlabel metal3 s 92303 57944 93103 58064 6 addr[12]
port 6 nsew signal input
rlabel metal3 s 92303 58488 93103 58608 6 addr[13]
port 7 nsew signal input
rlabel metal3 s 92303 59032 93103 59152 6 addr[14]
port 8 nsew signal input
rlabel metal3 s 92303 59576 93103 59696 6 addr[15]
port 9 nsew signal input
rlabel metal3 s 92303 60120 93103 60240 6 addr[16]
port 10 nsew signal input
rlabel metal3 s 92303 60664 93103 60784 6 addr[17]
port 11 nsew signal input
rlabel metal3 s 92303 61208 93103 61328 6 addr[18]
port 12 nsew signal input
rlabel metal3 s 92303 61752 93103 61872 6 addr[19]
port 13 nsew signal input
rlabel metal3 s 92303 51960 93103 52080 6 addr[1]
port 14 nsew signal input
rlabel metal3 s 92303 62296 93103 62416 6 addr[20]
port 15 nsew signal input
rlabel metal3 s 92303 62840 93103 62960 6 addr[21]
port 16 nsew signal input
rlabel metal3 s 92303 63384 93103 63504 6 addr[22]
port 17 nsew signal input
rlabel metal3 s 92303 63928 93103 64048 6 addr[23]
port 18 nsew signal input
rlabel metal3 s 92303 52504 93103 52624 6 addr[2]
port 19 nsew signal input
rlabel metal3 s 92303 53048 93103 53168 6 addr[3]
port 20 nsew signal input
rlabel metal3 s 92303 53592 93103 53712 6 addr[4]
port 21 nsew signal input
rlabel metal3 s 92303 54136 93103 54256 6 addr[5]
port 22 nsew signal input
rlabel metal3 s 92303 54680 93103 54800 6 addr[6]
port 23 nsew signal input
rlabel metal3 s 92303 55224 93103 55344 6 addr[7]
port 24 nsew signal input
rlabel metal3 s 92303 55768 93103 55888 6 addr[8]
port 25 nsew signal input
rlabel metal3 s 92303 56312 93103 56432 6 addr[9]
port 26 nsew signal input
rlabel metal3 s 92303 16056 93103 16176 6 cfgreg_di[0]
port 27 nsew signal input
rlabel metal3 s 92303 21496 93103 21616 6 cfgreg_di[10]
port 28 nsew signal input
rlabel metal3 s 92303 22040 93103 22160 6 cfgreg_di[11]
port 29 nsew signal input
rlabel metal3 s 92303 22584 93103 22704 6 cfgreg_di[12]
port 30 nsew signal input
rlabel metal3 s 92303 23128 93103 23248 6 cfgreg_di[13]
port 31 nsew signal input
rlabel metal3 s 92303 23672 93103 23792 6 cfgreg_di[14]
port 32 nsew signal input
rlabel metal3 s 92303 24216 93103 24336 6 cfgreg_di[15]
port 33 nsew signal input
rlabel metal3 s 92303 24760 93103 24880 6 cfgreg_di[16]
port 34 nsew signal input
rlabel metal3 s 92303 25304 93103 25424 6 cfgreg_di[17]
port 35 nsew signal input
rlabel metal3 s 92303 25848 93103 25968 6 cfgreg_di[18]
port 36 nsew signal input
rlabel metal3 s 92303 26392 93103 26512 6 cfgreg_di[19]
port 37 nsew signal input
rlabel metal3 s 92303 16600 93103 16720 6 cfgreg_di[1]
port 38 nsew signal input
rlabel metal3 s 92303 26936 93103 27056 6 cfgreg_di[20]
port 39 nsew signal input
rlabel metal3 s 92303 27480 93103 27600 6 cfgreg_di[21]
port 40 nsew signal input
rlabel metal3 s 92303 28024 93103 28144 6 cfgreg_di[22]
port 41 nsew signal input
rlabel metal3 s 92303 28568 93103 28688 6 cfgreg_di[23]
port 42 nsew signal input
rlabel metal3 s 92303 29112 93103 29232 6 cfgreg_di[24]
port 43 nsew signal input
rlabel metal3 s 92303 29656 93103 29776 6 cfgreg_di[25]
port 44 nsew signal input
rlabel metal3 s 92303 30200 93103 30320 6 cfgreg_di[26]
port 45 nsew signal input
rlabel metal3 s 92303 30744 93103 30864 6 cfgreg_di[27]
port 46 nsew signal input
rlabel metal3 s 92303 31288 93103 31408 6 cfgreg_di[28]
port 47 nsew signal input
rlabel metal3 s 92303 31832 93103 31952 6 cfgreg_di[29]
port 48 nsew signal input
rlabel metal3 s 92303 17144 93103 17264 6 cfgreg_di[2]
port 49 nsew signal input
rlabel metal3 s 92303 32376 93103 32496 6 cfgreg_di[30]
port 50 nsew signal input
rlabel metal3 s 92303 32920 93103 33040 6 cfgreg_di[31]
port 51 nsew signal input
rlabel metal3 s 92303 17688 93103 17808 6 cfgreg_di[3]
port 52 nsew signal input
rlabel metal3 s 92303 18232 93103 18352 6 cfgreg_di[4]
port 53 nsew signal input
rlabel metal3 s 92303 18776 93103 18896 6 cfgreg_di[5]
port 54 nsew signal input
rlabel metal3 s 92303 19320 93103 19440 6 cfgreg_di[6]
port 55 nsew signal input
rlabel metal3 s 92303 19864 93103 19984 6 cfgreg_di[7]
port 56 nsew signal input
rlabel metal3 s 92303 20408 93103 20528 6 cfgreg_di[8]
port 57 nsew signal input
rlabel metal3 s 92303 20952 93103 21072 6 cfgreg_di[9]
port 58 nsew signal input
rlabel metal3 s 92303 33464 93103 33584 6 cfgreg_do[0]
port 59 nsew signal output
rlabel metal3 s 92303 38904 93103 39024 6 cfgreg_do[10]
port 60 nsew signal output
rlabel metal3 s 92303 39448 93103 39568 6 cfgreg_do[11]
port 61 nsew signal output
rlabel metal3 s 92303 39992 93103 40112 6 cfgreg_do[12]
port 62 nsew signal output
rlabel metal3 s 92303 40536 93103 40656 6 cfgreg_do[13]
port 63 nsew signal output
rlabel metal3 s 92303 41080 93103 41200 6 cfgreg_do[14]
port 64 nsew signal output
rlabel metal3 s 92303 41624 93103 41744 6 cfgreg_do[15]
port 65 nsew signal output
rlabel metal3 s 92303 42168 93103 42288 6 cfgreg_do[16]
port 66 nsew signal output
rlabel metal3 s 92303 42712 93103 42832 6 cfgreg_do[17]
port 67 nsew signal output
rlabel metal3 s 92303 43256 93103 43376 6 cfgreg_do[18]
port 68 nsew signal output
rlabel metal3 s 92303 43800 93103 43920 6 cfgreg_do[19]
port 69 nsew signal output
rlabel metal3 s 92303 34008 93103 34128 6 cfgreg_do[1]
port 70 nsew signal output
rlabel metal3 s 92303 44344 93103 44464 6 cfgreg_do[20]
port 71 nsew signal output
rlabel metal3 s 92303 44888 93103 45008 6 cfgreg_do[21]
port 72 nsew signal output
rlabel metal3 s 92303 45432 93103 45552 6 cfgreg_do[22]
port 73 nsew signal output
rlabel metal3 s 92303 45976 93103 46096 6 cfgreg_do[23]
port 74 nsew signal output
rlabel metal3 s 92303 46520 93103 46640 6 cfgreg_do[24]
port 75 nsew signal output
rlabel metal3 s 92303 47064 93103 47184 6 cfgreg_do[25]
port 76 nsew signal output
rlabel metal3 s 92303 47608 93103 47728 6 cfgreg_do[26]
port 77 nsew signal output
rlabel metal3 s 92303 48152 93103 48272 6 cfgreg_do[27]
port 78 nsew signal output
rlabel metal3 s 92303 48696 93103 48816 6 cfgreg_do[28]
port 79 nsew signal output
rlabel metal3 s 92303 49240 93103 49360 6 cfgreg_do[29]
port 80 nsew signal output
rlabel metal3 s 92303 34552 93103 34672 6 cfgreg_do[2]
port 81 nsew signal output
rlabel metal3 s 92303 49784 93103 49904 6 cfgreg_do[30]
port 82 nsew signal output
rlabel metal3 s 92303 50328 93103 50448 6 cfgreg_do[31]
port 83 nsew signal output
rlabel metal3 s 92303 35096 93103 35216 6 cfgreg_do[3]
port 84 nsew signal output
rlabel metal3 s 92303 35640 93103 35760 6 cfgreg_do[4]
port 85 nsew signal output
rlabel metal3 s 92303 36184 93103 36304 6 cfgreg_do[5]
port 86 nsew signal output
rlabel metal3 s 92303 36728 93103 36848 6 cfgreg_do[6]
port 87 nsew signal output
rlabel metal3 s 92303 37272 93103 37392 6 cfgreg_do[7]
port 88 nsew signal output
rlabel metal3 s 92303 37816 93103 37936 6 cfgreg_do[8]
port 89 nsew signal output
rlabel metal3 s 92303 38360 93103 38480 6 cfgreg_do[9]
port 90 nsew signal output
rlabel metal3 s 92303 13880 93103 14000 6 cfgreg_we[0]
port 91 nsew signal input
rlabel metal3 s 92303 14424 93103 14544 6 cfgreg_we[1]
port 92 nsew signal input
rlabel metal3 s 92303 14968 93103 15088 6 cfgreg_we[2]
port 93 nsew signal input
rlabel metal3 s 92303 15512 93103 15632 6 cfgreg_we[3]
port 94 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 clk
port 95 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 flash_clk
port 96 nsew signal output
rlabel metal3 s 0 84872 800 84992 6 flash_csb
port 97 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 flash_io0_di
port 98 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 flash_io0_do
port 99 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 flash_io0_oe
port 100 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 flash_io1_di
port 101 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 flash_io1_do
port 102 nsew signal output
rlabel metal3 s 0 37272 800 37392 6 flash_io1_oe
port 103 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 flash_io2_di
port 104 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 flash_io2_do
port 105 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 flash_io2_oe
port 106 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 flash_io3_di
port 107 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 flash_io3_do
port 108 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 flash_io3_oe
port 109 nsew signal output
rlabel metal3 s 92303 64472 93103 64592 6 rdata[0]
port 110 nsew signal output
rlabel metal3 s 92303 69912 93103 70032 6 rdata[10]
port 111 nsew signal output
rlabel metal3 s 92303 70456 93103 70576 6 rdata[11]
port 112 nsew signal output
rlabel metal3 s 92303 71000 93103 71120 6 rdata[12]
port 113 nsew signal output
rlabel metal3 s 92303 71544 93103 71664 6 rdata[13]
port 114 nsew signal output
rlabel metal3 s 92303 72088 93103 72208 6 rdata[14]
port 115 nsew signal output
rlabel metal3 s 92303 72632 93103 72752 6 rdata[15]
port 116 nsew signal output
rlabel metal3 s 92303 73176 93103 73296 6 rdata[16]
port 117 nsew signal output
rlabel metal3 s 92303 73720 93103 73840 6 rdata[17]
port 118 nsew signal output
rlabel metal3 s 92303 74264 93103 74384 6 rdata[18]
port 119 nsew signal output
rlabel metal3 s 92303 74808 93103 74928 6 rdata[19]
port 120 nsew signal output
rlabel metal3 s 92303 65016 93103 65136 6 rdata[1]
port 121 nsew signal output
rlabel metal3 s 92303 75352 93103 75472 6 rdata[20]
port 122 nsew signal output
rlabel metal3 s 92303 75896 93103 76016 6 rdata[21]
port 123 nsew signal output
rlabel metal3 s 92303 76440 93103 76560 6 rdata[22]
port 124 nsew signal output
rlabel metal3 s 92303 76984 93103 77104 6 rdata[23]
port 125 nsew signal output
rlabel metal3 s 92303 77528 93103 77648 6 rdata[24]
port 126 nsew signal output
rlabel metal3 s 92303 78072 93103 78192 6 rdata[25]
port 127 nsew signal output
rlabel metal3 s 92303 78616 93103 78736 6 rdata[26]
port 128 nsew signal output
rlabel metal3 s 92303 79160 93103 79280 6 rdata[27]
port 129 nsew signal output
rlabel metal3 s 92303 79704 93103 79824 6 rdata[28]
port 130 nsew signal output
rlabel metal3 s 92303 80248 93103 80368 6 rdata[29]
port 131 nsew signal output
rlabel metal3 s 92303 65560 93103 65680 6 rdata[2]
port 132 nsew signal output
rlabel metal3 s 92303 80792 93103 80912 6 rdata[30]
port 133 nsew signal output
rlabel metal3 s 92303 81336 93103 81456 6 rdata[31]
port 134 nsew signal output
rlabel metal3 s 92303 66104 93103 66224 6 rdata[3]
port 135 nsew signal output
rlabel metal3 s 92303 66648 93103 66768 6 rdata[4]
port 136 nsew signal output
rlabel metal3 s 92303 67192 93103 67312 6 rdata[5]
port 137 nsew signal output
rlabel metal3 s 92303 67736 93103 67856 6 rdata[6]
port 138 nsew signal output
rlabel metal3 s 92303 68280 93103 68400 6 rdata[7]
port 139 nsew signal output
rlabel metal3 s 92303 68824 93103 68944 6 rdata[8]
port 140 nsew signal output
rlabel metal3 s 92303 69368 93103 69488 6 rdata[9]
port 141 nsew signal output
rlabel metal3 s 92303 50872 93103 50992 6 ready
port 142 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 resetn
port 143 nsew signal input
rlabel metal3 s 92303 13336 93103 13456 6 valid
port 144 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 93103 95247
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5713252
string GDS_FILE /openlane/designs/spimemio/runs/RUN_2023.12.03_10.14.21/results/signoff/spimemio.magic.gds
string GDS_START 688246
<< end >>

