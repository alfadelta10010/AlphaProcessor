module alphacore (clk,
    cpi_valid,
    cpi_wait,
    mem_instr,
    mem_la_read,
    mem_la_write,
    mem_ready,
    mem_valid,
    resetn,
    trace_valid,
    trap,
    cpi_insn,
    cpi_rs1,
    cpi_rs2,
    eoi,
    irq,
    mem_addr,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    mem_rdata,
    mem_wdata,
    mem_wstrb,
    trace_data);
 input clk;
 output cpi_valid;
 input cpi_wait;
 output mem_instr;
 output mem_la_read;
 output mem_la_write;
 input mem_ready;
 output mem_valid;
 input resetn;
 output trace_valid;
 output trap;
 output [31:0] cpi_insn;
 output [31:0] cpi_rs1;
 output [31:0] cpi_rs2;
 output [31:0] eoi;
 input [31:0] irq;
 output [31:0] mem_addr;
 output [31:0] mem_la_addr;
 output [31:0] mem_la_wdata;
 output [3:0] mem_la_wstrb;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;
 output [35:0] trace_data;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire \alu_out[0] ;
 wire \alu_out[10] ;
 wire \alu_out[11] ;
 wire \alu_out[12] ;
 wire \alu_out[13] ;
 wire \alu_out[14] ;
 wire \alu_out[15] ;
 wire \alu_out[16] ;
 wire \alu_out[17] ;
 wire \alu_out[18] ;
 wire \alu_out[19] ;
 wire \alu_out[1] ;
 wire \alu_out[20] ;
 wire \alu_out[21] ;
 wire \alu_out[22] ;
 wire \alu_out[23] ;
 wire \alu_out[24] ;
 wire \alu_out[25] ;
 wire \alu_out[26] ;
 wire \alu_out[27] ;
 wire \alu_out[28] ;
 wire \alu_out[29] ;
 wire \alu_out[2] ;
 wire \alu_out[30] ;
 wire \alu_out[31] ;
 wire \alu_out[3] ;
 wire \alu_out[4] ;
 wire \alu_out[5] ;
 wire \alu_out[6] ;
 wire \alu_out[7] ;
 wire \alu_out[8] ;
 wire \alu_out[9] ;
 wire \alu_out_q[0] ;
 wire \alu_out_q[10] ;
 wire \alu_out_q[11] ;
 wire \alu_out_q[12] ;
 wire \alu_out_q[13] ;
 wire \alu_out_q[14] ;
 wire \alu_out_q[15] ;
 wire \alu_out_q[16] ;
 wire \alu_out_q[17] ;
 wire \alu_out_q[18] ;
 wire \alu_out_q[19] ;
 wire \alu_out_q[1] ;
 wire \alu_out_q[20] ;
 wire \alu_out_q[21] ;
 wire \alu_out_q[22] ;
 wire \alu_out_q[23] ;
 wire \alu_out_q[24] ;
 wire \alu_out_q[25] ;
 wire \alu_out_q[26] ;
 wire \alu_out_q[27] ;
 wire \alu_out_q[28] ;
 wire \alu_out_q[29] ;
 wire \alu_out_q[2] ;
 wire \alu_out_q[30] ;
 wire \alu_out_q[31] ;
 wire \alu_out_q[3] ;
 wire \alu_out_q[4] ;
 wire \alu_out_q[5] ;
 wire \alu_out_q[6] ;
 wire \alu_out_q[7] ;
 wire \alu_out_q[8] ;
 wire \alu_out_q[9] ;
 wire clear_prefetched_high_word;
 wire clear_prefetched_high_word_q;
 wire compressed_instr;
 wire \count_cycle[0] ;
 wire \count_cycle[10] ;
 wire \count_cycle[11] ;
 wire \count_cycle[12] ;
 wire \count_cycle[13] ;
 wire \count_cycle[14] ;
 wire \count_cycle[15] ;
 wire \count_cycle[16] ;
 wire \count_cycle[17] ;
 wire \count_cycle[18] ;
 wire \count_cycle[19] ;
 wire \count_cycle[1] ;
 wire \count_cycle[20] ;
 wire \count_cycle[21] ;
 wire \count_cycle[22] ;
 wire \count_cycle[23] ;
 wire \count_cycle[24] ;
 wire \count_cycle[25] ;
 wire \count_cycle[26] ;
 wire \count_cycle[27] ;
 wire \count_cycle[28] ;
 wire \count_cycle[29] ;
 wire \count_cycle[2] ;
 wire \count_cycle[30] ;
 wire \count_cycle[31] ;
 wire \count_cycle[32] ;
 wire \count_cycle[33] ;
 wire \count_cycle[34] ;
 wire \count_cycle[35] ;
 wire \count_cycle[36] ;
 wire \count_cycle[37] ;
 wire \count_cycle[38] ;
 wire \count_cycle[39] ;
 wire \count_cycle[3] ;
 wire \count_cycle[40] ;
 wire \count_cycle[41] ;
 wire \count_cycle[42] ;
 wire \count_cycle[43] ;
 wire \count_cycle[44] ;
 wire \count_cycle[45] ;
 wire \count_cycle[46] ;
 wire \count_cycle[47] ;
 wire \count_cycle[48] ;
 wire \count_cycle[49] ;
 wire \count_cycle[4] ;
 wire \count_cycle[50] ;
 wire \count_cycle[51] ;
 wire \count_cycle[52] ;
 wire \count_cycle[53] ;
 wire \count_cycle[54] ;
 wire \count_cycle[55] ;
 wire \count_cycle[56] ;
 wire \count_cycle[57] ;
 wire \count_cycle[58] ;
 wire \count_cycle[59] ;
 wire \count_cycle[5] ;
 wire \count_cycle[60] ;
 wire \count_cycle[61] ;
 wire \count_cycle[62] ;
 wire \count_cycle[63] ;
 wire \count_cycle[6] ;
 wire \count_cycle[7] ;
 wire \count_cycle[8] ;
 wire \count_cycle[9] ;
 wire \count_instr[0] ;
 wire \count_instr[10] ;
 wire \count_instr[11] ;
 wire \count_instr[12] ;
 wire \count_instr[13] ;
 wire \count_instr[14] ;
 wire \count_instr[15] ;
 wire \count_instr[16] ;
 wire \count_instr[17] ;
 wire \count_instr[18] ;
 wire \count_instr[19] ;
 wire \count_instr[1] ;
 wire \count_instr[20] ;
 wire \count_instr[21] ;
 wire \count_instr[22] ;
 wire \count_instr[23] ;
 wire \count_instr[24] ;
 wire \count_instr[25] ;
 wire \count_instr[26] ;
 wire \count_instr[27] ;
 wire \count_instr[28] ;
 wire \count_instr[29] ;
 wire \count_instr[2] ;
 wire \count_instr[30] ;
 wire \count_instr[31] ;
 wire \count_instr[32] ;
 wire \count_instr[33] ;
 wire \count_instr[34] ;
 wire \count_instr[35] ;
 wire \count_instr[36] ;
 wire \count_instr[37] ;
 wire \count_instr[38] ;
 wire \count_instr[39] ;
 wire \count_instr[3] ;
 wire \count_instr[40] ;
 wire \count_instr[41] ;
 wire \count_instr[42] ;
 wire \count_instr[43] ;
 wire \count_instr[44] ;
 wire \count_instr[45] ;
 wire \count_instr[46] ;
 wire \count_instr[47] ;
 wire \count_instr[48] ;
 wire \count_instr[49] ;
 wire \count_instr[4] ;
 wire \count_instr[50] ;
 wire \count_instr[51] ;
 wire \count_instr[52] ;
 wire \count_instr[53] ;
 wire \count_instr[54] ;
 wire \count_instr[55] ;
 wire \count_instr[56] ;
 wire \count_instr[57] ;
 wire \count_instr[58] ;
 wire \count_instr[59] ;
 wire \count_instr[5] ;
 wire \count_instr[60] ;
 wire \count_instr[61] ;
 wire \count_instr[62] ;
 wire \count_instr[63] ;
 wire \count_instr[6] ;
 wire \count_instr[7] ;
 wire \count_instr[8] ;
 wire \count_instr[9] ;
 wire net303;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net304;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net305;
 wire net333;
 wire net334;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net335;
 wire \cpu_state[0] ;
 wire \cpu_state[1] ;
 wire \cpu_state[2] ;
 wire \cpu_state[3] ;
 wire \cpu_state[4] ;
 wire \cpu_state[5] ;
 wire \cpu_state[6] ;
 wire \cpuregs.raddr1[0] ;
 wire \cpuregs.raddr1[1] ;
 wire \cpuregs.raddr1[2] ;
 wire \cpuregs.raddr1[3] ;
 wire \cpuregs.raddr1[4] ;
 wire \cpuregs.raddr2[0] ;
 wire \cpuregs.raddr2[1] ;
 wire \cpuregs.raddr2[2] ;
 wire \cpuregs.raddr2[3] ;
 wire \cpuregs.raddr2[4] ;
 wire \cpuregs.regs[0][0] ;
 wire \cpuregs.regs[0][10] ;
 wire \cpuregs.regs[0][11] ;
 wire \cpuregs.regs[0][12] ;
 wire \cpuregs.regs[0][13] ;
 wire \cpuregs.regs[0][14] ;
 wire \cpuregs.regs[0][15] ;
 wire \cpuregs.regs[0][16] ;
 wire \cpuregs.regs[0][17] ;
 wire \cpuregs.regs[0][18] ;
 wire \cpuregs.regs[0][19] ;
 wire \cpuregs.regs[0][1] ;
 wire \cpuregs.regs[0][20] ;
 wire \cpuregs.regs[0][21] ;
 wire \cpuregs.regs[0][22] ;
 wire \cpuregs.regs[0][23] ;
 wire \cpuregs.regs[0][24] ;
 wire \cpuregs.regs[0][25] ;
 wire \cpuregs.regs[0][26] ;
 wire \cpuregs.regs[0][27] ;
 wire \cpuregs.regs[0][28] ;
 wire \cpuregs.regs[0][29] ;
 wire \cpuregs.regs[0][2] ;
 wire \cpuregs.regs[0][30] ;
 wire \cpuregs.regs[0][31] ;
 wire \cpuregs.regs[0][3] ;
 wire \cpuregs.regs[0][4] ;
 wire \cpuregs.regs[0][5] ;
 wire \cpuregs.regs[0][6] ;
 wire \cpuregs.regs[0][7] ;
 wire \cpuregs.regs[0][8] ;
 wire \cpuregs.regs[0][9] ;
 wire \cpuregs.regs[10][0] ;
 wire \cpuregs.regs[10][10] ;
 wire \cpuregs.regs[10][11] ;
 wire \cpuregs.regs[10][12] ;
 wire \cpuregs.regs[10][13] ;
 wire \cpuregs.regs[10][14] ;
 wire \cpuregs.regs[10][15] ;
 wire \cpuregs.regs[10][16] ;
 wire \cpuregs.regs[10][17] ;
 wire \cpuregs.regs[10][18] ;
 wire \cpuregs.regs[10][19] ;
 wire \cpuregs.regs[10][1] ;
 wire \cpuregs.regs[10][20] ;
 wire \cpuregs.regs[10][21] ;
 wire \cpuregs.regs[10][22] ;
 wire \cpuregs.regs[10][23] ;
 wire \cpuregs.regs[10][24] ;
 wire \cpuregs.regs[10][25] ;
 wire \cpuregs.regs[10][26] ;
 wire \cpuregs.regs[10][27] ;
 wire \cpuregs.regs[10][28] ;
 wire \cpuregs.regs[10][29] ;
 wire \cpuregs.regs[10][2] ;
 wire \cpuregs.regs[10][30] ;
 wire \cpuregs.regs[10][31] ;
 wire \cpuregs.regs[10][3] ;
 wire \cpuregs.regs[10][4] ;
 wire \cpuregs.regs[10][5] ;
 wire \cpuregs.regs[10][6] ;
 wire \cpuregs.regs[10][7] ;
 wire \cpuregs.regs[10][8] ;
 wire \cpuregs.regs[10][9] ;
 wire \cpuregs.regs[11][0] ;
 wire \cpuregs.regs[11][10] ;
 wire \cpuregs.regs[11][11] ;
 wire \cpuregs.regs[11][12] ;
 wire \cpuregs.regs[11][13] ;
 wire \cpuregs.regs[11][14] ;
 wire \cpuregs.regs[11][15] ;
 wire \cpuregs.regs[11][16] ;
 wire \cpuregs.regs[11][17] ;
 wire \cpuregs.regs[11][18] ;
 wire \cpuregs.regs[11][19] ;
 wire \cpuregs.regs[11][1] ;
 wire \cpuregs.regs[11][20] ;
 wire \cpuregs.regs[11][21] ;
 wire \cpuregs.regs[11][22] ;
 wire \cpuregs.regs[11][23] ;
 wire \cpuregs.regs[11][24] ;
 wire \cpuregs.regs[11][25] ;
 wire \cpuregs.regs[11][26] ;
 wire \cpuregs.regs[11][27] ;
 wire \cpuregs.regs[11][28] ;
 wire \cpuregs.regs[11][29] ;
 wire \cpuregs.regs[11][2] ;
 wire \cpuregs.regs[11][30] ;
 wire \cpuregs.regs[11][31] ;
 wire \cpuregs.regs[11][3] ;
 wire \cpuregs.regs[11][4] ;
 wire \cpuregs.regs[11][5] ;
 wire \cpuregs.regs[11][6] ;
 wire \cpuregs.regs[11][7] ;
 wire \cpuregs.regs[11][8] ;
 wire \cpuregs.regs[11][9] ;
 wire \cpuregs.regs[12][0] ;
 wire \cpuregs.regs[12][10] ;
 wire \cpuregs.regs[12][11] ;
 wire \cpuregs.regs[12][12] ;
 wire \cpuregs.regs[12][13] ;
 wire \cpuregs.regs[12][14] ;
 wire \cpuregs.regs[12][15] ;
 wire \cpuregs.regs[12][16] ;
 wire \cpuregs.regs[12][17] ;
 wire \cpuregs.regs[12][18] ;
 wire \cpuregs.regs[12][19] ;
 wire \cpuregs.regs[12][1] ;
 wire \cpuregs.regs[12][20] ;
 wire \cpuregs.regs[12][21] ;
 wire \cpuregs.regs[12][22] ;
 wire \cpuregs.regs[12][23] ;
 wire \cpuregs.regs[12][24] ;
 wire \cpuregs.regs[12][25] ;
 wire \cpuregs.regs[12][26] ;
 wire \cpuregs.regs[12][27] ;
 wire \cpuregs.regs[12][28] ;
 wire \cpuregs.regs[12][29] ;
 wire \cpuregs.regs[12][2] ;
 wire \cpuregs.regs[12][30] ;
 wire \cpuregs.regs[12][31] ;
 wire \cpuregs.regs[12][3] ;
 wire \cpuregs.regs[12][4] ;
 wire \cpuregs.regs[12][5] ;
 wire \cpuregs.regs[12][6] ;
 wire \cpuregs.regs[12][7] ;
 wire \cpuregs.regs[12][8] ;
 wire \cpuregs.regs[12][9] ;
 wire \cpuregs.regs[13][0] ;
 wire \cpuregs.regs[13][10] ;
 wire \cpuregs.regs[13][11] ;
 wire \cpuregs.regs[13][12] ;
 wire \cpuregs.regs[13][13] ;
 wire \cpuregs.regs[13][14] ;
 wire \cpuregs.regs[13][15] ;
 wire \cpuregs.regs[13][16] ;
 wire \cpuregs.regs[13][17] ;
 wire \cpuregs.regs[13][18] ;
 wire \cpuregs.regs[13][19] ;
 wire \cpuregs.regs[13][1] ;
 wire \cpuregs.regs[13][20] ;
 wire \cpuregs.regs[13][21] ;
 wire \cpuregs.regs[13][22] ;
 wire \cpuregs.regs[13][23] ;
 wire \cpuregs.regs[13][24] ;
 wire \cpuregs.regs[13][25] ;
 wire \cpuregs.regs[13][26] ;
 wire \cpuregs.regs[13][27] ;
 wire \cpuregs.regs[13][28] ;
 wire \cpuregs.regs[13][29] ;
 wire \cpuregs.regs[13][2] ;
 wire \cpuregs.regs[13][30] ;
 wire \cpuregs.regs[13][31] ;
 wire \cpuregs.regs[13][3] ;
 wire \cpuregs.regs[13][4] ;
 wire \cpuregs.regs[13][5] ;
 wire \cpuregs.regs[13][6] ;
 wire \cpuregs.regs[13][7] ;
 wire \cpuregs.regs[13][8] ;
 wire \cpuregs.regs[13][9] ;
 wire \cpuregs.regs[14][0] ;
 wire \cpuregs.regs[14][10] ;
 wire \cpuregs.regs[14][11] ;
 wire \cpuregs.regs[14][12] ;
 wire \cpuregs.regs[14][13] ;
 wire \cpuregs.regs[14][14] ;
 wire \cpuregs.regs[14][15] ;
 wire \cpuregs.regs[14][16] ;
 wire \cpuregs.regs[14][17] ;
 wire \cpuregs.regs[14][18] ;
 wire \cpuregs.regs[14][19] ;
 wire \cpuregs.regs[14][1] ;
 wire \cpuregs.regs[14][20] ;
 wire \cpuregs.regs[14][21] ;
 wire \cpuregs.regs[14][22] ;
 wire \cpuregs.regs[14][23] ;
 wire \cpuregs.regs[14][24] ;
 wire \cpuregs.regs[14][25] ;
 wire \cpuregs.regs[14][26] ;
 wire \cpuregs.regs[14][27] ;
 wire \cpuregs.regs[14][28] ;
 wire \cpuregs.regs[14][29] ;
 wire \cpuregs.regs[14][2] ;
 wire \cpuregs.regs[14][30] ;
 wire \cpuregs.regs[14][31] ;
 wire \cpuregs.regs[14][3] ;
 wire \cpuregs.regs[14][4] ;
 wire \cpuregs.regs[14][5] ;
 wire \cpuregs.regs[14][6] ;
 wire \cpuregs.regs[14][7] ;
 wire \cpuregs.regs[14][8] ;
 wire \cpuregs.regs[14][9] ;
 wire \cpuregs.regs[15][0] ;
 wire \cpuregs.regs[15][10] ;
 wire \cpuregs.regs[15][11] ;
 wire \cpuregs.regs[15][12] ;
 wire \cpuregs.regs[15][13] ;
 wire \cpuregs.regs[15][14] ;
 wire \cpuregs.regs[15][15] ;
 wire \cpuregs.regs[15][16] ;
 wire \cpuregs.regs[15][17] ;
 wire \cpuregs.regs[15][18] ;
 wire \cpuregs.regs[15][19] ;
 wire \cpuregs.regs[15][1] ;
 wire \cpuregs.regs[15][20] ;
 wire \cpuregs.regs[15][21] ;
 wire \cpuregs.regs[15][22] ;
 wire \cpuregs.regs[15][23] ;
 wire \cpuregs.regs[15][24] ;
 wire \cpuregs.regs[15][25] ;
 wire \cpuregs.regs[15][26] ;
 wire \cpuregs.regs[15][27] ;
 wire \cpuregs.regs[15][28] ;
 wire \cpuregs.regs[15][29] ;
 wire \cpuregs.regs[15][2] ;
 wire \cpuregs.regs[15][30] ;
 wire \cpuregs.regs[15][31] ;
 wire \cpuregs.regs[15][3] ;
 wire \cpuregs.regs[15][4] ;
 wire \cpuregs.regs[15][5] ;
 wire \cpuregs.regs[15][6] ;
 wire \cpuregs.regs[15][7] ;
 wire \cpuregs.regs[15][8] ;
 wire \cpuregs.regs[15][9] ;
 wire \cpuregs.regs[16][0] ;
 wire \cpuregs.regs[16][10] ;
 wire \cpuregs.regs[16][11] ;
 wire \cpuregs.regs[16][12] ;
 wire \cpuregs.regs[16][13] ;
 wire \cpuregs.regs[16][14] ;
 wire \cpuregs.regs[16][15] ;
 wire \cpuregs.regs[16][16] ;
 wire \cpuregs.regs[16][17] ;
 wire \cpuregs.regs[16][18] ;
 wire \cpuregs.regs[16][19] ;
 wire \cpuregs.regs[16][1] ;
 wire \cpuregs.regs[16][20] ;
 wire \cpuregs.regs[16][21] ;
 wire \cpuregs.regs[16][22] ;
 wire \cpuregs.regs[16][23] ;
 wire \cpuregs.regs[16][24] ;
 wire \cpuregs.regs[16][25] ;
 wire \cpuregs.regs[16][26] ;
 wire \cpuregs.regs[16][27] ;
 wire \cpuregs.regs[16][28] ;
 wire \cpuregs.regs[16][29] ;
 wire \cpuregs.regs[16][2] ;
 wire \cpuregs.regs[16][30] ;
 wire \cpuregs.regs[16][31] ;
 wire \cpuregs.regs[16][3] ;
 wire \cpuregs.regs[16][4] ;
 wire \cpuregs.regs[16][5] ;
 wire \cpuregs.regs[16][6] ;
 wire \cpuregs.regs[16][7] ;
 wire \cpuregs.regs[16][8] ;
 wire \cpuregs.regs[16][9] ;
 wire \cpuregs.regs[17][0] ;
 wire \cpuregs.regs[17][10] ;
 wire \cpuregs.regs[17][11] ;
 wire \cpuregs.regs[17][12] ;
 wire \cpuregs.regs[17][13] ;
 wire \cpuregs.regs[17][14] ;
 wire \cpuregs.regs[17][15] ;
 wire \cpuregs.regs[17][16] ;
 wire \cpuregs.regs[17][17] ;
 wire \cpuregs.regs[17][18] ;
 wire \cpuregs.regs[17][19] ;
 wire \cpuregs.regs[17][1] ;
 wire \cpuregs.regs[17][20] ;
 wire \cpuregs.regs[17][21] ;
 wire \cpuregs.regs[17][22] ;
 wire \cpuregs.regs[17][23] ;
 wire \cpuregs.regs[17][24] ;
 wire \cpuregs.regs[17][25] ;
 wire \cpuregs.regs[17][26] ;
 wire \cpuregs.regs[17][27] ;
 wire \cpuregs.regs[17][28] ;
 wire \cpuregs.regs[17][29] ;
 wire \cpuregs.regs[17][2] ;
 wire \cpuregs.regs[17][30] ;
 wire \cpuregs.regs[17][31] ;
 wire \cpuregs.regs[17][3] ;
 wire \cpuregs.regs[17][4] ;
 wire \cpuregs.regs[17][5] ;
 wire \cpuregs.regs[17][6] ;
 wire \cpuregs.regs[17][7] ;
 wire \cpuregs.regs[17][8] ;
 wire \cpuregs.regs[17][9] ;
 wire \cpuregs.regs[18][0] ;
 wire \cpuregs.regs[18][10] ;
 wire \cpuregs.regs[18][11] ;
 wire \cpuregs.regs[18][12] ;
 wire \cpuregs.regs[18][13] ;
 wire \cpuregs.regs[18][14] ;
 wire \cpuregs.regs[18][15] ;
 wire \cpuregs.regs[18][16] ;
 wire \cpuregs.regs[18][17] ;
 wire \cpuregs.regs[18][18] ;
 wire \cpuregs.regs[18][19] ;
 wire \cpuregs.regs[18][1] ;
 wire \cpuregs.regs[18][20] ;
 wire \cpuregs.regs[18][21] ;
 wire \cpuregs.regs[18][22] ;
 wire \cpuregs.regs[18][23] ;
 wire \cpuregs.regs[18][24] ;
 wire \cpuregs.regs[18][25] ;
 wire \cpuregs.regs[18][26] ;
 wire \cpuregs.regs[18][27] ;
 wire \cpuregs.regs[18][28] ;
 wire \cpuregs.regs[18][29] ;
 wire \cpuregs.regs[18][2] ;
 wire \cpuregs.regs[18][30] ;
 wire \cpuregs.regs[18][31] ;
 wire \cpuregs.regs[18][3] ;
 wire \cpuregs.regs[18][4] ;
 wire \cpuregs.regs[18][5] ;
 wire \cpuregs.regs[18][6] ;
 wire \cpuregs.regs[18][7] ;
 wire \cpuregs.regs[18][8] ;
 wire \cpuregs.regs[18][9] ;
 wire \cpuregs.regs[19][0] ;
 wire \cpuregs.regs[19][10] ;
 wire \cpuregs.regs[19][11] ;
 wire \cpuregs.regs[19][12] ;
 wire \cpuregs.regs[19][13] ;
 wire \cpuregs.regs[19][14] ;
 wire \cpuregs.regs[19][15] ;
 wire \cpuregs.regs[19][16] ;
 wire \cpuregs.regs[19][17] ;
 wire \cpuregs.regs[19][18] ;
 wire \cpuregs.regs[19][19] ;
 wire \cpuregs.regs[19][1] ;
 wire \cpuregs.regs[19][20] ;
 wire \cpuregs.regs[19][21] ;
 wire \cpuregs.regs[19][22] ;
 wire \cpuregs.regs[19][23] ;
 wire \cpuregs.regs[19][24] ;
 wire \cpuregs.regs[19][25] ;
 wire \cpuregs.regs[19][26] ;
 wire \cpuregs.regs[19][27] ;
 wire \cpuregs.regs[19][28] ;
 wire \cpuregs.regs[19][29] ;
 wire \cpuregs.regs[19][2] ;
 wire \cpuregs.regs[19][30] ;
 wire \cpuregs.regs[19][31] ;
 wire \cpuregs.regs[19][3] ;
 wire \cpuregs.regs[19][4] ;
 wire \cpuregs.regs[19][5] ;
 wire \cpuregs.regs[19][6] ;
 wire \cpuregs.regs[19][7] ;
 wire \cpuregs.regs[19][8] ;
 wire \cpuregs.regs[19][9] ;
 wire \cpuregs.regs[1][0] ;
 wire \cpuregs.regs[1][10] ;
 wire \cpuregs.regs[1][11] ;
 wire \cpuregs.regs[1][12] ;
 wire \cpuregs.regs[1][13] ;
 wire \cpuregs.regs[1][14] ;
 wire \cpuregs.regs[1][15] ;
 wire \cpuregs.regs[1][16] ;
 wire \cpuregs.regs[1][17] ;
 wire \cpuregs.regs[1][18] ;
 wire \cpuregs.regs[1][19] ;
 wire \cpuregs.regs[1][1] ;
 wire \cpuregs.regs[1][20] ;
 wire \cpuregs.regs[1][21] ;
 wire \cpuregs.regs[1][22] ;
 wire \cpuregs.regs[1][23] ;
 wire \cpuregs.regs[1][24] ;
 wire \cpuregs.regs[1][25] ;
 wire \cpuregs.regs[1][26] ;
 wire \cpuregs.regs[1][27] ;
 wire \cpuregs.regs[1][28] ;
 wire \cpuregs.regs[1][29] ;
 wire \cpuregs.regs[1][2] ;
 wire \cpuregs.regs[1][30] ;
 wire \cpuregs.regs[1][31] ;
 wire \cpuregs.regs[1][3] ;
 wire \cpuregs.regs[1][4] ;
 wire \cpuregs.regs[1][5] ;
 wire \cpuregs.regs[1][6] ;
 wire \cpuregs.regs[1][7] ;
 wire \cpuregs.regs[1][8] ;
 wire \cpuregs.regs[1][9] ;
 wire \cpuregs.regs[20][0] ;
 wire \cpuregs.regs[20][10] ;
 wire \cpuregs.regs[20][11] ;
 wire \cpuregs.regs[20][12] ;
 wire \cpuregs.regs[20][13] ;
 wire \cpuregs.regs[20][14] ;
 wire \cpuregs.regs[20][15] ;
 wire \cpuregs.regs[20][16] ;
 wire \cpuregs.regs[20][17] ;
 wire \cpuregs.regs[20][18] ;
 wire \cpuregs.regs[20][19] ;
 wire \cpuregs.regs[20][1] ;
 wire \cpuregs.regs[20][20] ;
 wire \cpuregs.regs[20][21] ;
 wire \cpuregs.regs[20][22] ;
 wire \cpuregs.regs[20][23] ;
 wire \cpuregs.regs[20][24] ;
 wire \cpuregs.regs[20][25] ;
 wire \cpuregs.regs[20][26] ;
 wire \cpuregs.regs[20][27] ;
 wire \cpuregs.regs[20][28] ;
 wire \cpuregs.regs[20][29] ;
 wire \cpuregs.regs[20][2] ;
 wire \cpuregs.regs[20][30] ;
 wire \cpuregs.regs[20][31] ;
 wire \cpuregs.regs[20][3] ;
 wire \cpuregs.regs[20][4] ;
 wire \cpuregs.regs[20][5] ;
 wire \cpuregs.regs[20][6] ;
 wire \cpuregs.regs[20][7] ;
 wire \cpuregs.regs[20][8] ;
 wire \cpuregs.regs[20][9] ;
 wire \cpuregs.regs[21][0] ;
 wire \cpuregs.regs[21][10] ;
 wire \cpuregs.regs[21][11] ;
 wire \cpuregs.regs[21][12] ;
 wire \cpuregs.regs[21][13] ;
 wire \cpuregs.regs[21][14] ;
 wire \cpuregs.regs[21][15] ;
 wire \cpuregs.regs[21][16] ;
 wire \cpuregs.regs[21][17] ;
 wire \cpuregs.regs[21][18] ;
 wire \cpuregs.regs[21][19] ;
 wire \cpuregs.regs[21][1] ;
 wire \cpuregs.regs[21][20] ;
 wire \cpuregs.regs[21][21] ;
 wire \cpuregs.regs[21][22] ;
 wire \cpuregs.regs[21][23] ;
 wire \cpuregs.regs[21][24] ;
 wire \cpuregs.regs[21][25] ;
 wire \cpuregs.regs[21][26] ;
 wire \cpuregs.regs[21][27] ;
 wire \cpuregs.regs[21][28] ;
 wire \cpuregs.regs[21][29] ;
 wire \cpuregs.regs[21][2] ;
 wire \cpuregs.regs[21][30] ;
 wire \cpuregs.regs[21][31] ;
 wire \cpuregs.regs[21][3] ;
 wire \cpuregs.regs[21][4] ;
 wire \cpuregs.regs[21][5] ;
 wire \cpuregs.regs[21][6] ;
 wire \cpuregs.regs[21][7] ;
 wire \cpuregs.regs[21][8] ;
 wire \cpuregs.regs[21][9] ;
 wire \cpuregs.regs[22][0] ;
 wire \cpuregs.regs[22][10] ;
 wire \cpuregs.regs[22][11] ;
 wire \cpuregs.regs[22][12] ;
 wire \cpuregs.regs[22][13] ;
 wire \cpuregs.regs[22][14] ;
 wire \cpuregs.regs[22][15] ;
 wire \cpuregs.regs[22][16] ;
 wire \cpuregs.regs[22][17] ;
 wire \cpuregs.regs[22][18] ;
 wire \cpuregs.regs[22][19] ;
 wire \cpuregs.regs[22][1] ;
 wire \cpuregs.regs[22][20] ;
 wire \cpuregs.regs[22][21] ;
 wire \cpuregs.regs[22][22] ;
 wire \cpuregs.regs[22][23] ;
 wire \cpuregs.regs[22][24] ;
 wire \cpuregs.regs[22][25] ;
 wire \cpuregs.regs[22][26] ;
 wire \cpuregs.regs[22][27] ;
 wire \cpuregs.regs[22][28] ;
 wire \cpuregs.regs[22][29] ;
 wire \cpuregs.regs[22][2] ;
 wire \cpuregs.regs[22][30] ;
 wire \cpuregs.regs[22][31] ;
 wire \cpuregs.regs[22][3] ;
 wire \cpuregs.regs[22][4] ;
 wire \cpuregs.regs[22][5] ;
 wire \cpuregs.regs[22][6] ;
 wire \cpuregs.regs[22][7] ;
 wire \cpuregs.regs[22][8] ;
 wire \cpuregs.regs[22][9] ;
 wire \cpuregs.regs[23][0] ;
 wire \cpuregs.regs[23][10] ;
 wire \cpuregs.regs[23][11] ;
 wire \cpuregs.regs[23][12] ;
 wire \cpuregs.regs[23][13] ;
 wire \cpuregs.regs[23][14] ;
 wire \cpuregs.regs[23][15] ;
 wire \cpuregs.regs[23][16] ;
 wire \cpuregs.regs[23][17] ;
 wire \cpuregs.regs[23][18] ;
 wire \cpuregs.regs[23][19] ;
 wire \cpuregs.regs[23][1] ;
 wire \cpuregs.regs[23][20] ;
 wire \cpuregs.regs[23][21] ;
 wire \cpuregs.regs[23][22] ;
 wire \cpuregs.regs[23][23] ;
 wire \cpuregs.regs[23][24] ;
 wire \cpuregs.regs[23][25] ;
 wire \cpuregs.regs[23][26] ;
 wire \cpuregs.regs[23][27] ;
 wire \cpuregs.regs[23][28] ;
 wire \cpuregs.regs[23][29] ;
 wire \cpuregs.regs[23][2] ;
 wire \cpuregs.regs[23][30] ;
 wire \cpuregs.regs[23][31] ;
 wire \cpuregs.regs[23][3] ;
 wire \cpuregs.regs[23][4] ;
 wire \cpuregs.regs[23][5] ;
 wire \cpuregs.regs[23][6] ;
 wire \cpuregs.regs[23][7] ;
 wire \cpuregs.regs[23][8] ;
 wire \cpuregs.regs[23][9] ;
 wire \cpuregs.regs[24][0] ;
 wire \cpuregs.regs[24][10] ;
 wire \cpuregs.regs[24][11] ;
 wire \cpuregs.regs[24][12] ;
 wire \cpuregs.regs[24][13] ;
 wire \cpuregs.regs[24][14] ;
 wire \cpuregs.regs[24][15] ;
 wire \cpuregs.regs[24][16] ;
 wire \cpuregs.regs[24][17] ;
 wire \cpuregs.regs[24][18] ;
 wire \cpuregs.regs[24][19] ;
 wire \cpuregs.regs[24][1] ;
 wire \cpuregs.regs[24][20] ;
 wire \cpuregs.regs[24][21] ;
 wire \cpuregs.regs[24][22] ;
 wire \cpuregs.regs[24][23] ;
 wire \cpuregs.regs[24][24] ;
 wire \cpuregs.regs[24][25] ;
 wire \cpuregs.regs[24][26] ;
 wire \cpuregs.regs[24][27] ;
 wire \cpuregs.regs[24][28] ;
 wire \cpuregs.regs[24][29] ;
 wire \cpuregs.regs[24][2] ;
 wire \cpuregs.regs[24][30] ;
 wire \cpuregs.regs[24][31] ;
 wire \cpuregs.regs[24][3] ;
 wire \cpuregs.regs[24][4] ;
 wire \cpuregs.regs[24][5] ;
 wire \cpuregs.regs[24][6] ;
 wire \cpuregs.regs[24][7] ;
 wire \cpuregs.regs[24][8] ;
 wire \cpuregs.regs[24][9] ;
 wire \cpuregs.regs[25][0] ;
 wire \cpuregs.regs[25][10] ;
 wire \cpuregs.regs[25][11] ;
 wire \cpuregs.regs[25][12] ;
 wire \cpuregs.regs[25][13] ;
 wire \cpuregs.regs[25][14] ;
 wire \cpuregs.regs[25][15] ;
 wire \cpuregs.regs[25][16] ;
 wire \cpuregs.regs[25][17] ;
 wire \cpuregs.regs[25][18] ;
 wire \cpuregs.regs[25][19] ;
 wire \cpuregs.regs[25][1] ;
 wire \cpuregs.regs[25][20] ;
 wire \cpuregs.regs[25][21] ;
 wire \cpuregs.regs[25][22] ;
 wire \cpuregs.regs[25][23] ;
 wire \cpuregs.regs[25][24] ;
 wire \cpuregs.regs[25][25] ;
 wire \cpuregs.regs[25][26] ;
 wire \cpuregs.regs[25][27] ;
 wire \cpuregs.regs[25][28] ;
 wire \cpuregs.regs[25][29] ;
 wire \cpuregs.regs[25][2] ;
 wire \cpuregs.regs[25][30] ;
 wire \cpuregs.regs[25][31] ;
 wire \cpuregs.regs[25][3] ;
 wire \cpuregs.regs[25][4] ;
 wire \cpuregs.regs[25][5] ;
 wire \cpuregs.regs[25][6] ;
 wire \cpuregs.regs[25][7] ;
 wire \cpuregs.regs[25][8] ;
 wire \cpuregs.regs[25][9] ;
 wire \cpuregs.regs[26][0] ;
 wire \cpuregs.regs[26][10] ;
 wire \cpuregs.regs[26][11] ;
 wire \cpuregs.regs[26][12] ;
 wire \cpuregs.regs[26][13] ;
 wire \cpuregs.regs[26][14] ;
 wire \cpuregs.regs[26][15] ;
 wire \cpuregs.regs[26][16] ;
 wire \cpuregs.regs[26][17] ;
 wire \cpuregs.regs[26][18] ;
 wire \cpuregs.regs[26][19] ;
 wire \cpuregs.regs[26][1] ;
 wire \cpuregs.regs[26][20] ;
 wire \cpuregs.regs[26][21] ;
 wire \cpuregs.regs[26][22] ;
 wire \cpuregs.regs[26][23] ;
 wire \cpuregs.regs[26][24] ;
 wire \cpuregs.regs[26][25] ;
 wire \cpuregs.regs[26][26] ;
 wire \cpuregs.regs[26][27] ;
 wire \cpuregs.regs[26][28] ;
 wire \cpuregs.regs[26][29] ;
 wire \cpuregs.regs[26][2] ;
 wire \cpuregs.regs[26][30] ;
 wire \cpuregs.regs[26][31] ;
 wire \cpuregs.regs[26][3] ;
 wire \cpuregs.regs[26][4] ;
 wire \cpuregs.regs[26][5] ;
 wire \cpuregs.regs[26][6] ;
 wire \cpuregs.regs[26][7] ;
 wire \cpuregs.regs[26][8] ;
 wire \cpuregs.regs[26][9] ;
 wire \cpuregs.regs[27][0] ;
 wire \cpuregs.regs[27][10] ;
 wire \cpuregs.regs[27][11] ;
 wire \cpuregs.regs[27][12] ;
 wire \cpuregs.regs[27][13] ;
 wire \cpuregs.regs[27][14] ;
 wire \cpuregs.regs[27][15] ;
 wire \cpuregs.regs[27][16] ;
 wire \cpuregs.regs[27][17] ;
 wire \cpuregs.regs[27][18] ;
 wire \cpuregs.regs[27][19] ;
 wire \cpuregs.regs[27][1] ;
 wire \cpuregs.regs[27][20] ;
 wire \cpuregs.regs[27][21] ;
 wire \cpuregs.regs[27][22] ;
 wire \cpuregs.regs[27][23] ;
 wire \cpuregs.regs[27][24] ;
 wire \cpuregs.regs[27][25] ;
 wire \cpuregs.regs[27][26] ;
 wire \cpuregs.regs[27][27] ;
 wire \cpuregs.regs[27][28] ;
 wire \cpuregs.regs[27][29] ;
 wire \cpuregs.regs[27][2] ;
 wire \cpuregs.regs[27][30] ;
 wire \cpuregs.regs[27][31] ;
 wire \cpuregs.regs[27][3] ;
 wire \cpuregs.regs[27][4] ;
 wire \cpuregs.regs[27][5] ;
 wire \cpuregs.regs[27][6] ;
 wire \cpuregs.regs[27][7] ;
 wire \cpuregs.regs[27][8] ;
 wire \cpuregs.regs[27][9] ;
 wire \cpuregs.regs[28][0] ;
 wire \cpuregs.regs[28][10] ;
 wire \cpuregs.regs[28][11] ;
 wire \cpuregs.regs[28][12] ;
 wire \cpuregs.regs[28][13] ;
 wire \cpuregs.regs[28][14] ;
 wire \cpuregs.regs[28][15] ;
 wire \cpuregs.regs[28][16] ;
 wire \cpuregs.regs[28][17] ;
 wire \cpuregs.regs[28][18] ;
 wire \cpuregs.regs[28][19] ;
 wire \cpuregs.regs[28][1] ;
 wire \cpuregs.regs[28][20] ;
 wire \cpuregs.regs[28][21] ;
 wire \cpuregs.regs[28][22] ;
 wire \cpuregs.regs[28][23] ;
 wire \cpuregs.regs[28][24] ;
 wire \cpuregs.regs[28][25] ;
 wire \cpuregs.regs[28][26] ;
 wire \cpuregs.regs[28][27] ;
 wire \cpuregs.regs[28][28] ;
 wire \cpuregs.regs[28][29] ;
 wire \cpuregs.regs[28][2] ;
 wire \cpuregs.regs[28][30] ;
 wire \cpuregs.regs[28][31] ;
 wire \cpuregs.regs[28][3] ;
 wire \cpuregs.regs[28][4] ;
 wire \cpuregs.regs[28][5] ;
 wire \cpuregs.regs[28][6] ;
 wire \cpuregs.regs[28][7] ;
 wire \cpuregs.regs[28][8] ;
 wire \cpuregs.regs[28][9] ;
 wire \cpuregs.regs[29][0] ;
 wire \cpuregs.regs[29][10] ;
 wire \cpuregs.regs[29][11] ;
 wire \cpuregs.regs[29][12] ;
 wire \cpuregs.regs[29][13] ;
 wire \cpuregs.regs[29][14] ;
 wire \cpuregs.regs[29][15] ;
 wire \cpuregs.regs[29][16] ;
 wire \cpuregs.regs[29][17] ;
 wire \cpuregs.regs[29][18] ;
 wire \cpuregs.regs[29][19] ;
 wire \cpuregs.regs[29][1] ;
 wire \cpuregs.regs[29][20] ;
 wire \cpuregs.regs[29][21] ;
 wire \cpuregs.regs[29][22] ;
 wire \cpuregs.regs[29][23] ;
 wire \cpuregs.regs[29][24] ;
 wire \cpuregs.regs[29][25] ;
 wire \cpuregs.regs[29][26] ;
 wire \cpuregs.regs[29][27] ;
 wire \cpuregs.regs[29][28] ;
 wire \cpuregs.regs[29][29] ;
 wire \cpuregs.regs[29][2] ;
 wire \cpuregs.regs[29][30] ;
 wire \cpuregs.regs[29][31] ;
 wire \cpuregs.regs[29][3] ;
 wire \cpuregs.regs[29][4] ;
 wire \cpuregs.regs[29][5] ;
 wire \cpuregs.regs[29][6] ;
 wire \cpuregs.regs[29][7] ;
 wire \cpuregs.regs[29][8] ;
 wire \cpuregs.regs[29][9] ;
 wire \cpuregs.regs[2][0] ;
 wire \cpuregs.regs[2][10] ;
 wire \cpuregs.regs[2][11] ;
 wire \cpuregs.regs[2][12] ;
 wire \cpuregs.regs[2][13] ;
 wire \cpuregs.regs[2][14] ;
 wire \cpuregs.regs[2][15] ;
 wire \cpuregs.regs[2][16] ;
 wire \cpuregs.regs[2][17] ;
 wire \cpuregs.regs[2][18] ;
 wire \cpuregs.regs[2][19] ;
 wire \cpuregs.regs[2][1] ;
 wire \cpuregs.regs[2][20] ;
 wire \cpuregs.regs[2][21] ;
 wire \cpuregs.regs[2][22] ;
 wire \cpuregs.regs[2][23] ;
 wire \cpuregs.regs[2][24] ;
 wire \cpuregs.regs[2][25] ;
 wire \cpuregs.regs[2][26] ;
 wire \cpuregs.regs[2][27] ;
 wire \cpuregs.regs[2][28] ;
 wire \cpuregs.regs[2][29] ;
 wire \cpuregs.regs[2][2] ;
 wire \cpuregs.regs[2][30] ;
 wire \cpuregs.regs[2][31] ;
 wire \cpuregs.regs[2][3] ;
 wire \cpuregs.regs[2][4] ;
 wire \cpuregs.regs[2][5] ;
 wire \cpuregs.regs[2][6] ;
 wire \cpuregs.regs[2][7] ;
 wire \cpuregs.regs[2][8] ;
 wire \cpuregs.regs[2][9] ;
 wire \cpuregs.regs[30][0] ;
 wire \cpuregs.regs[30][10] ;
 wire \cpuregs.regs[30][11] ;
 wire \cpuregs.regs[30][12] ;
 wire \cpuregs.regs[30][13] ;
 wire \cpuregs.regs[30][14] ;
 wire \cpuregs.regs[30][15] ;
 wire \cpuregs.regs[30][16] ;
 wire \cpuregs.regs[30][17] ;
 wire \cpuregs.regs[30][18] ;
 wire \cpuregs.regs[30][19] ;
 wire \cpuregs.regs[30][1] ;
 wire \cpuregs.regs[30][20] ;
 wire \cpuregs.regs[30][21] ;
 wire \cpuregs.regs[30][22] ;
 wire \cpuregs.regs[30][23] ;
 wire \cpuregs.regs[30][24] ;
 wire \cpuregs.regs[30][25] ;
 wire \cpuregs.regs[30][26] ;
 wire \cpuregs.regs[30][27] ;
 wire \cpuregs.regs[30][28] ;
 wire \cpuregs.regs[30][29] ;
 wire \cpuregs.regs[30][2] ;
 wire \cpuregs.regs[30][30] ;
 wire \cpuregs.regs[30][31] ;
 wire \cpuregs.regs[30][3] ;
 wire \cpuregs.regs[30][4] ;
 wire \cpuregs.regs[30][5] ;
 wire \cpuregs.regs[30][6] ;
 wire \cpuregs.regs[30][7] ;
 wire \cpuregs.regs[30][8] ;
 wire \cpuregs.regs[30][9] ;
 wire \cpuregs.regs[31][0] ;
 wire \cpuregs.regs[31][10] ;
 wire \cpuregs.regs[31][11] ;
 wire \cpuregs.regs[31][12] ;
 wire \cpuregs.regs[31][13] ;
 wire \cpuregs.regs[31][14] ;
 wire \cpuregs.regs[31][15] ;
 wire \cpuregs.regs[31][16] ;
 wire \cpuregs.regs[31][17] ;
 wire \cpuregs.regs[31][18] ;
 wire \cpuregs.regs[31][19] ;
 wire \cpuregs.regs[31][1] ;
 wire \cpuregs.regs[31][20] ;
 wire \cpuregs.regs[31][21] ;
 wire \cpuregs.regs[31][22] ;
 wire \cpuregs.regs[31][23] ;
 wire \cpuregs.regs[31][24] ;
 wire \cpuregs.regs[31][25] ;
 wire \cpuregs.regs[31][26] ;
 wire \cpuregs.regs[31][27] ;
 wire \cpuregs.regs[31][28] ;
 wire \cpuregs.regs[31][29] ;
 wire \cpuregs.regs[31][2] ;
 wire \cpuregs.regs[31][30] ;
 wire \cpuregs.regs[31][31] ;
 wire \cpuregs.regs[31][3] ;
 wire \cpuregs.regs[31][4] ;
 wire \cpuregs.regs[31][5] ;
 wire \cpuregs.regs[31][6] ;
 wire \cpuregs.regs[31][7] ;
 wire \cpuregs.regs[31][8] ;
 wire \cpuregs.regs[31][9] ;
 wire \cpuregs.regs[3][0] ;
 wire \cpuregs.regs[3][10] ;
 wire \cpuregs.regs[3][11] ;
 wire \cpuregs.regs[3][12] ;
 wire \cpuregs.regs[3][13] ;
 wire \cpuregs.regs[3][14] ;
 wire \cpuregs.regs[3][15] ;
 wire \cpuregs.regs[3][16] ;
 wire \cpuregs.regs[3][17] ;
 wire \cpuregs.regs[3][18] ;
 wire \cpuregs.regs[3][19] ;
 wire \cpuregs.regs[3][1] ;
 wire \cpuregs.regs[3][20] ;
 wire \cpuregs.regs[3][21] ;
 wire \cpuregs.regs[3][22] ;
 wire \cpuregs.regs[3][23] ;
 wire \cpuregs.regs[3][24] ;
 wire \cpuregs.regs[3][25] ;
 wire \cpuregs.regs[3][26] ;
 wire \cpuregs.regs[3][27] ;
 wire \cpuregs.regs[3][28] ;
 wire \cpuregs.regs[3][29] ;
 wire \cpuregs.regs[3][2] ;
 wire \cpuregs.regs[3][30] ;
 wire \cpuregs.regs[3][31] ;
 wire \cpuregs.regs[3][3] ;
 wire \cpuregs.regs[3][4] ;
 wire \cpuregs.regs[3][5] ;
 wire \cpuregs.regs[3][6] ;
 wire \cpuregs.regs[3][7] ;
 wire \cpuregs.regs[3][8] ;
 wire \cpuregs.regs[3][9] ;
 wire \cpuregs.regs[4][0] ;
 wire \cpuregs.regs[4][10] ;
 wire \cpuregs.regs[4][11] ;
 wire \cpuregs.regs[4][12] ;
 wire \cpuregs.regs[4][13] ;
 wire \cpuregs.regs[4][14] ;
 wire \cpuregs.regs[4][15] ;
 wire \cpuregs.regs[4][16] ;
 wire \cpuregs.regs[4][17] ;
 wire \cpuregs.regs[4][18] ;
 wire \cpuregs.regs[4][19] ;
 wire \cpuregs.regs[4][1] ;
 wire \cpuregs.regs[4][20] ;
 wire \cpuregs.regs[4][21] ;
 wire \cpuregs.regs[4][22] ;
 wire \cpuregs.regs[4][23] ;
 wire \cpuregs.regs[4][24] ;
 wire \cpuregs.regs[4][25] ;
 wire \cpuregs.regs[4][26] ;
 wire \cpuregs.regs[4][27] ;
 wire \cpuregs.regs[4][28] ;
 wire \cpuregs.regs[4][29] ;
 wire \cpuregs.regs[4][2] ;
 wire \cpuregs.regs[4][30] ;
 wire \cpuregs.regs[4][31] ;
 wire \cpuregs.regs[4][3] ;
 wire \cpuregs.regs[4][4] ;
 wire \cpuregs.regs[4][5] ;
 wire \cpuregs.regs[4][6] ;
 wire \cpuregs.regs[4][7] ;
 wire \cpuregs.regs[4][8] ;
 wire \cpuregs.regs[4][9] ;
 wire \cpuregs.regs[5][0] ;
 wire \cpuregs.regs[5][10] ;
 wire \cpuregs.regs[5][11] ;
 wire \cpuregs.regs[5][12] ;
 wire \cpuregs.regs[5][13] ;
 wire \cpuregs.regs[5][14] ;
 wire \cpuregs.regs[5][15] ;
 wire \cpuregs.regs[5][16] ;
 wire \cpuregs.regs[5][17] ;
 wire \cpuregs.regs[5][18] ;
 wire \cpuregs.regs[5][19] ;
 wire \cpuregs.regs[5][1] ;
 wire \cpuregs.regs[5][20] ;
 wire \cpuregs.regs[5][21] ;
 wire \cpuregs.regs[5][22] ;
 wire \cpuregs.regs[5][23] ;
 wire \cpuregs.regs[5][24] ;
 wire \cpuregs.regs[5][25] ;
 wire \cpuregs.regs[5][26] ;
 wire \cpuregs.regs[5][27] ;
 wire \cpuregs.regs[5][28] ;
 wire \cpuregs.regs[5][29] ;
 wire \cpuregs.regs[5][2] ;
 wire \cpuregs.regs[5][30] ;
 wire \cpuregs.regs[5][31] ;
 wire \cpuregs.regs[5][3] ;
 wire \cpuregs.regs[5][4] ;
 wire \cpuregs.regs[5][5] ;
 wire \cpuregs.regs[5][6] ;
 wire \cpuregs.regs[5][7] ;
 wire \cpuregs.regs[5][8] ;
 wire \cpuregs.regs[5][9] ;
 wire \cpuregs.regs[6][0] ;
 wire \cpuregs.regs[6][10] ;
 wire \cpuregs.regs[6][11] ;
 wire \cpuregs.regs[6][12] ;
 wire \cpuregs.regs[6][13] ;
 wire \cpuregs.regs[6][14] ;
 wire \cpuregs.regs[6][15] ;
 wire \cpuregs.regs[6][16] ;
 wire \cpuregs.regs[6][17] ;
 wire \cpuregs.regs[6][18] ;
 wire \cpuregs.regs[6][19] ;
 wire \cpuregs.regs[6][1] ;
 wire \cpuregs.regs[6][20] ;
 wire \cpuregs.regs[6][21] ;
 wire \cpuregs.regs[6][22] ;
 wire \cpuregs.regs[6][23] ;
 wire \cpuregs.regs[6][24] ;
 wire \cpuregs.regs[6][25] ;
 wire \cpuregs.regs[6][26] ;
 wire \cpuregs.regs[6][27] ;
 wire \cpuregs.regs[6][28] ;
 wire \cpuregs.regs[6][29] ;
 wire \cpuregs.regs[6][2] ;
 wire \cpuregs.regs[6][30] ;
 wire \cpuregs.regs[6][31] ;
 wire \cpuregs.regs[6][3] ;
 wire \cpuregs.regs[6][4] ;
 wire \cpuregs.regs[6][5] ;
 wire \cpuregs.regs[6][6] ;
 wire \cpuregs.regs[6][7] ;
 wire \cpuregs.regs[6][8] ;
 wire \cpuregs.regs[6][9] ;
 wire \cpuregs.regs[7][0] ;
 wire \cpuregs.regs[7][10] ;
 wire \cpuregs.regs[7][11] ;
 wire \cpuregs.regs[7][12] ;
 wire \cpuregs.regs[7][13] ;
 wire \cpuregs.regs[7][14] ;
 wire \cpuregs.regs[7][15] ;
 wire \cpuregs.regs[7][16] ;
 wire \cpuregs.regs[7][17] ;
 wire \cpuregs.regs[7][18] ;
 wire \cpuregs.regs[7][19] ;
 wire \cpuregs.regs[7][1] ;
 wire \cpuregs.regs[7][20] ;
 wire \cpuregs.regs[7][21] ;
 wire \cpuregs.regs[7][22] ;
 wire \cpuregs.regs[7][23] ;
 wire \cpuregs.regs[7][24] ;
 wire \cpuregs.regs[7][25] ;
 wire \cpuregs.regs[7][26] ;
 wire \cpuregs.regs[7][27] ;
 wire \cpuregs.regs[7][28] ;
 wire \cpuregs.regs[7][29] ;
 wire \cpuregs.regs[7][2] ;
 wire \cpuregs.regs[7][30] ;
 wire \cpuregs.regs[7][31] ;
 wire \cpuregs.regs[7][3] ;
 wire \cpuregs.regs[7][4] ;
 wire \cpuregs.regs[7][5] ;
 wire \cpuregs.regs[7][6] ;
 wire \cpuregs.regs[7][7] ;
 wire \cpuregs.regs[7][8] ;
 wire \cpuregs.regs[7][9] ;
 wire \cpuregs.regs[8][0] ;
 wire \cpuregs.regs[8][10] ;
 wire \cpuregs.regs[8][11] ;
 wire \cpuregs.regs[8][12] ;
 wire \cpuregs.regs[8][13] ;
 wire \cpuregs.regs[8][14] ;
 wire \cpuregs.regs[8][15] ;
 wire \cpuregs.regs[8][16] ;
 wire \cpuregs.regs[8][17] ;
 wire \cpuregs.regs[8][18] ;
 wire \cpuregs.regs[8][19] ;
 wire \cpuregs.regs[8][1] ;
 wire \cpuregs.regs[8][20] ;
 wire \cpuregs.regs[8][21] ;
 wire \cpuregs.regs[8][22] ;
 wire \cpuregs.regs[8][23] ;
 wire \cpuregs.regs[8][24] ;
 wire \cpuregs.regs[8][25] ;
 wire \cpuregs.regs[8][26] ;
 wire \cpuregs.regs[8][27] ;
 wire \cpuregs.regs[8][28] ;
 wire \cpuregs.regs[8][29] ;
 wire \cpuregs.regs[8][2] ;
 wire \cpuregs.regs[8][30] ;
 wire \cpuregs.regs[8][31] ;
 wire \cpuregs.regs[8][3] ;
 wire \cpuregs.regs[8][4] ;
 wire \cpuregs.regs[8][5] ;
 wire \cpuregs.regs[8][6] ;
 wire \cpuregs.regs[8][7] ;
 wire \cpuregs.regs[8][8] ;
 wire \cpuregs.regs[8][9] ;
 wire \cpuregs.regs[9][0] ;
 wire \cpuregs.regs[9][10] ;
 wire \cpuregs.regs[9][11] ;
 wire \cpuregs.regs[9][12] ;
 wire \cpuregs.regs[9][13] ;
 wire \cpuregs.regs[9][14] ;
 wire \cpuregs.regs[9][15] ;
 wire \cpuregs.regs[9][16] ;
 wire \cpuregs.regs[9][17] ;
 wire \cpuregs.regs[9][18] ;
 wire \cpuregs.regs[9][19] ;
 wire \cpuregs.regs[9][1] ;
 wire \cpuregs.regs[9][20] ;
 wire \cpuregs.regs[9][21] ;
 wire \cpuregs.regs[9][22] ;
 wire \cpuregs.regs[9][23] ;
 wire \cpuregs.regs[9][24] ;
 wire \cpuregs.regs[9][25] ;
 wire \cpuregs.regs[9][26] ;
 wire \cpuregs.regs[9][27] ;
 wire \cpuregs.regs[9][28] ;
 wire \cpuregs.regs[9][29] ;
 wire \cpuregs.regs[9][2] ;
 wire \cpuregs.regs[9][30] ;
 wire \cpuregs.regs[9][31] ;
 wire \cpuregs.regs[9][3] ;
 wire \cpuregs.regs[9][4] ;
 wire \cpuregs.regs[9][5] ;
 wire \cpuregs.regs[9][6] ;
 wire \cpuregs.regs[9][7] ;
 wire \cpuregs.regs[9][8] ;
 wire \cpuregs.regs[9][9] ;
 wire \cpuregs.waddr[0] ;
 wire \cpuregs.waddr[1] ;
 wire \cpuregs.waddr[2] ;
 wire \cpuregs.waddr[3] ;
 wire \cpuregs.waddr[4] ;
 wire \decoded_imm[0] ;
 wire \decoded_imm[10] ;
 wire \decoded_imm[11] ;
 wire \decoded_imm[12] ;
 wire \decoded_imm[13] ;
 wire \decoded_imm[14] ;
 wire \decoded_imm[15] ;
 wire \decoded_imm[16] ;
 wire \decoded_imm[17] ;
 wire \decoded_imm[18] ;
 wire \decoded_imm[19] ;
 wire \decoded_imm[1] ;
 wire \decoded_imm[20] ;
 wire \decoded_imm[21] ;
 wire \decoded_imm[22] ;
 wire \decoded_imm[23] ;
 wire \decoded_imm[24] ;
 wire \decoded_imm[25] ;
 wire \decoded_imm[26] ;
 wire \decoded_imm[27] ;
 wire \decoded_imm[28] ;
 wire \decoded_imm[29] ;
 wire \decoded_imm[2] ;
 wire \decoded_imm[30] ;
 wire \decoded_imm[31] ;
 wire \decoded_imm[3] ;
 wire \decoded_imm[4] ;
 wire \decoded_imm[5] ;
 wire \decoded_imm[6] ;
 wire \decoded_imm[7] ;
 wire \decoded_imm[8] ;
 wire \decoded_imm[9] ;
 wire \decoded_imm_j[10] ;
 wire \decoded_imm_j[11] ;
 wire \decoded_imm_j[12] ;
 wire \decoded_imm_j[13] ;
 wire \decoded_imm_j[14] ;
 wire \decoded_imm_j[15] ;
 wire \decoded_imm_j[16] ;
 wire \decoded_imm_j[17] ;
 wire \decoded_imm_j[18] ;
 wire \decoded_imm_j[19] ;
 wire \decoded_imm_j[1] ;
 wire \decoded_imm_j[20] ;
 wire \decoded_imm_j[2] ;
 wire \decoded_imm_j[3] ;
 wire \decoded_imm_j[4] ;
 wire \decoded_imm_j[5] ;
 wire \decoded_imm_j[6] ;
 wire \decoded_imm_j[7] ;
 wire \decoded_imm_j[8] ;
 wire \decoded_imm_j[9] ;
 wire \decoded_rd[0] ;
 wire \decoded_rd[1] ;
 wire \decoded_rd[2] ;
 wire \decoded_rd[3] ;
 wire \decoded_rd[4] ;
 wire decoder_pseudo_trigger;
 wire decoder_trigger;
 wire do_waitirq;
 wire instr_add;
 wire instr_addi;
 wire instr_and;
 wire instr_andi;
 wire instr_auipc;
 wire instr_beq;
 wire instr_bge;
 wire instr_bgeu;
 wire instr_blt;
 wire instr_bltu;
 wire instr_bne;
 wire instr_fence;
 wire instr_jal;
 wire instr_jalr;
 wire instr_lb;
 wire instr_lbu;
 wire instr_lh;
 wire instr_lhu;
 wire instr_lui;
 wire instr_lw;
 wire instr_maskirq;
 wire instr_or;
 wire instr_ori;
 wire instr_rdcycle;
 wire instr_rdcycleh;
 wire instr_rdinstr;
 wire instr_rdinstrh;
 wire instr_retirq;
 wire instr_sb;
 wire instr_sh;
 wire instr_sll;
 wire instr_slli;
 wire instr_slt;
 wire instr_slti;
 wire instr_sltiu;
 wire instr_sltu;
 wire instr_sra;
 wire instr_srai;
 wire instr_srl;
 wire instr_srli;
 wire instr_sub;
 wire instr_sw;
 wire instr_timer;
 wire instr_waitirq;
 wire instr_xor;
 wire instr_xori;
 wire irq_active;
 wire irq_delay;
 wire \irq_mask[0] ;
 wire \irq_mask[10] ;
 wire \irq_mask[11] ;
 wire \irq_mask[12] ;
 wire \irq_mask[13] ;
 wire \irq_mask[14] ;
 wire \irq_mask[15] ;
 wire \irq_mask[16] ;
 wire \irq_mask[17] ;
 wire \irq_mask[18] ;
 wire \irq_mask[19] ;
 wire \irq_mask[1] ;
 wire \irq_mask[20] ;
 wire \irq_mask[21] ;
 wire \irq_mask[22] ;
 wire \irq_mask[23] ;
 wire \irq_mask[24] ;
 wire \irq_mask[25] ;
 wire \irq_mask[26] ;
 wire \irq_mask[27] ;
 wire \irq_mask[28] ;
 wire \irq_mask[29] ;
 wire \irq_mask[2] ;
 wire \irq_mask[30] ;
 wire \irq_mask[31] ;
 wire \irq_mask[3] ;
 wire \irq_mask[4] ;
 wire \irq_mask[5] ;
 wire \irq_mask[6] ;
 wire \irq_mask[7] ;
 wire \irq_mask[8] ;
 wire \irq_mask[9] ;
 wire \irq_pending[0] ;
 wire \irq_pending[10] ;
 wire \irq_pending[11] ;
 wire \irq_pending[12] ;
 wire \irq_pending[13] ;
 wire \irq_pending[14] ;
 wire \irq_pending[15] ;
 wire \irq_pending[16] ;
 wire \irq_pending[17] ;
 wire \irq_pending[18] ;
 wire \irq_pending[19] ;
 wire \irq_pending[1] ;
 wire \irq_pending[20] ;
 wire \irq_pending[21] ;
 wire \irq_pending[22] ;
 wire \irq_pending[23] ;
 wire \irq_pending[24] ;
 wire \irq_pending[25] ;
 wire \irq_pending[26] ;
 wire \irq_pending[27] ;
 wire \irq_pending[28] ;
 wire \irq_pending[29] ;
 wire \irq_pending[2] ;
 wire \irq_pending[30] ;
 wire \irq_pending[31] ;
 wire \irq_pending[3] ;
 wire \irq_pending[4] ;
 wire \irq_pending[5] ;
 wire \irq_pending[6] ;
 wire \irq_pending[7] ;
 wire \irq_pending[8] ;
 wire \irq_pending[9] ;
 wire \irq_state[0] ;
 wire \irq_state[1] ;
 wire is_alu_reg_imm;
 wire is_alu_reg_reg;
 wire is_beq_bne_blt_bge_bltu_bgeu;
 wire is_compare;
 wire is_jalr_addi_slti_sltiu_xori_ori_andi;
 wire is_lb_lh_lw_lbu_lhu;
 wire is_lui_auipc_jal;
 wire is_sb_sh_sw;
 wire is_slli_srli_srai;
 wire is_slti_blt_slt;
 wire is_sltiu_bltu_sltu;
 wire last_mem_valid;
 wire latched_branch;
 wire latched_compr;
 wire latched_is_lb;
 wire latched_is_lh;
 wire latched_stalu;
 wire latched_store;
 wire \mem_16bit_buffer[0] ;
 wire \mem_16bit_buffer[10] ;
 wire \mem_16bit_buffer[11] ;
 wire \mem_16bit_buffer[12] ;
 wire \mem_16bit_buffer[13] ;
 wire \mem_16bit_buffer[14] ;
 wire \mem_16bit_buffer[15] ;
 wire \mem_16bit_buffer[1] ;
 wire \mem_16bit_buffer[2] ;
 wire \mem_16bit_buffer[3] ;
 wire \mem_16bit_buffer[4] ;
 wire \mem_16bit_buffer[5] ;
 wire \mem_16bit_buffer[6] ;
 wire \mem_16bit_buffer[7] ;
 wire \mem_16bit_buffer[8] ;
 wire \mem_16bit_buffer[9] ;
 wire net336;
 wire net337;
 wire mem_do_prefetch;
 wire mem_do_rdata;
 wire mem_do_rinst;
 wire mem_do_wdata;
 wire net338;
 wire net339;
 wire mem_la_firstword_reg;
 wire mem_la_secondword;
 wire \mem_rdata_q[0] ;
 wire \mem_rdata_q[10] ;
 wire \mem_rdata_q[11] ;
 wire \mem_rdata_q[12] ;
 wire \mem_rdata_q[13] ;
 wire \mem_rdata_q[14] ;
 wire \mem_rdata_q[15] ;
 wire \mem_rdata_q[16] ;
 wire \mem_rdata_q[17] ;
 wire \mem_rdata_q[18] ;
 wire \mem_rdata_q[19] ;
 wire \mem_rdata_q[1] ;
 wire \mem_rdata_q[20] ;
 wire \mem_rdata_q[21] ;
 wire \mem_rdata_q[22] ;
 wire \mem_rdata_q[23] ;
 wire \mem_rdata_q[24] ;
 wire \mem_rdata_q[25] ;
 wire \mem_rdata_q[26] ;
 wire \mem_rdata_q[27] ;
 wire \mem_rdata_q[28] ;
 wire \mem_rdata_q[29] ;
 wire \mem_rdata_q[2] ;
 wire \mem_rdata_q[30] ;
 wire \mem_rdata_q[31] ;
 wire \mem_rdata_q[3] ;
 wire \mem_rdata_q[4] ;
 wire \mem_rdata_q[5] ;
 wire \mem_rdata_q[6] ;
 wire \mem_rdata_q[7] ;
 wire \mem_rdata_q[8] ;
 wire \mem_rdata_q[9] ;
 wire \mem_state[0] ;
 wire \mem_state[1] ;
 wire \mem_wordsize[0] ;
 wire \mem_wordsize[1] ;
 wire \mem_wordsize[2] ;
 wire prefetched_high_word;
 wire \reg_next_pc[0] ;
 wire \reg_next_pc[10] ;
 wire \reg_next_pc[11] ;
 wire \reg_next_pc[12] ;
 wire \reg_next_pc[13] ;
 wire \reg_next_pc[14] ;
 wire \reg_next_pc[15] ;
 wire \reg_next_pc[16] ;
 wire \reg_next_pc[17] ;
 wire \reg_next_pc[18] ;
 wire \reg_next_pc[19] ;
 wire \reg_next_pc[1] ;
 wire \reg_next_pc[20] ;
 wire \reg_next_pc[21] ;
 wire \reg_next_pc[22] ;
 wire \reg_next_pc[23] ;
 wire \reg_next_pc[24] ;
 wire \reg_next_pc[25] ;
 wire \reg_next_pc[26] ;
 wire \reg_next_pc[27] ;
 wire \reg_next_pc[28] ;
 wire \reg_next_pc[29] ;
 wire \reg_next_pc[2] ;
 wire \reg_next_pc[30] ;
 wire \reg_next_pc[31] ;
 wire \reg_next_pc[3] ;
 wire \reg_next_pc[4] ;
 wire \reg_next_pc[5] ;
 wire \reg_next_pc[6] ;
 wire \reg_next_pc[7] ;
 wire \reg_next_pc[8] ;
 wire \reg_next_pc[9] ;
 wire \reg_out[0] ;
 wire \reg_out[10] ;
 wire \reg_out[11] ;
 wire \reg_out[12] ;
 wire \reg_out[13] ;
 wire \reg_out[14] ;
 wire \reg_out[15] ;
 wire \reg_out[16] ;
 wire \reg_out[17] ;
 wire \reg_out[18] ;
 wire \reg_out[19] ;
 wire \reg_out[1] ;
 wire \reg_out[20] ;
 wire \reg_out[21] ;
 wire \reg_out[22] ;
 wire \reg_out[23] ;
 wire \reg_out[24] ;
 wire \reg_out[25] ;
 wire \reg_out[26] ;
 wire \reg_out[27] ;
 wire \reg_out[28] ;
 wire \reg_out[29] ;
 wire \reg_out[2] ;
 wire \reg_out[30] ;
 wire \reg_out[31] ;
 wire \reg_out[3] ;
 wire \reg_out[4] ;
 wire \reg_out[5] ;
 wire \reg_out[6] ;
 wire \reg_out[7] ;
 wire \reg_out[8] ;
 wire \reg_out[9] ;
 wire \reg_pc[10] ;
 wire \reg_pc[11] ;
 wire \reg_pc[12] ;
 wire \reg_pc[13] ;
 wire \reg_pc[14] ;
 wire \reg_pc[15] ;
 wire \reg_pc[16] ;
 wire \reg_pc[17] ;
 wire \reg_pc[18] ;
 wire \reg_pc[19] ;
 wire \reg_pc[1] ;
 wire \reg_pc[20] ;
 wire \reg_pc[21] ;
 wire \reg_pc[22] ;
 wire \reg_pc[23] ;
 wire \reg_pc[24] ;
 wire \reg_pc[25] ;
 wire \reg_pc[26] ;
 wire \reg_pc[27] ;
 wire \reg_pc[28] ;
 wire \reg_pc[29] ;
 wire \reg_pc[2] ;
 wire \reg_pc[30] ;
 wire \reg_pc[31] ;
 wire \reg_pc[3] ;
 wire \reg_pc[4] ;
 wire \reg_pc[5] ;
 wire \reg_pc[6] ;
 wire \reg_pc[7] ;
 wire \reg_pc[8] ;
 wire \reg_pc[9] ;
 wire \reg_sh[0] ;
 wire \reg_sh[1] ;
 wire \reg_sh[2] ;
 wire \reg_sh[3] ;
 wire \reg_sh[4] ;
 wire \timer[0] ;
 wire \timer[10] ;
 wire \timer[11] ;
 wire \timer[12] ;
 wire \timer[13] ;
 wire \timer[14] ;
 wire \timer[15] ;
 wire \timer[16] ;
 wire \timer[17] ;
 wire \timer[18] ;
 wire \timer[19] ;
 wire \timer[1] ;
 wire \timer[20] ;
 wire \timer[21] ;
 wire \timer[22] ;
 wire \timer[23] ;
 wire \timer[24] ;
 wire \timer[25] ;
 wire \timer[26] ;
 wire \timer[27] ;
 wire \timer[28] ;
 wire \timer[29] ;
 wire \timer[2] ;
 wire \timer[30] ;
 wire \timer[31] ;
 wire \timer[3] ;
 wire \timer[4] ;
 wire \timer[5] ;
 wire \timer[6] ;
 wire \timer[7] ;
 wire \timer[8] ;
 wire \timer[9] ;
 wire net340;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net341;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net342;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire clknet_leaf_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sky130_fd_sc_hd__inv_2 _08401_ (.A(mem_la_secondword),
    .Y(_03187_));
 sky130_fd_sc_hd__nand2_1 _08402_ (.A(latched_branch),
    .B(latched_store),
    .Y(_03188_));
 sky130_fd_sc_hd__and2_2 _08403_ (.A(latched_branch),
    .B(latched_store),
    .X(_03189_));
 sky130_fd_sc_hd__or2_1 _08404_ (.A(\reg_next_pc[1] ),
    .B(_03189_),
    .X(_03190_));
 sky130_fd_sc_hd__o21ai_2 _08405_ (.A1(\reg_out[1] ),
    .A2(_03188_),
    .B1(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__or2_1 _08406_ (.A(mem_do_rinst),
    .B(mem_do_prefetch),
    .X(_03192_));
 sky130_fd_sc_hd__and3b_1 _08407_ (.A_N(_03191_),
    .B(_03192_),
    .C(_03187_),
    .X(_03193_));
 sky130_fd_sc_hd__or2_1 _08408_ (.A(\irq_state[1] ),
    .B(\irq_state[0] ),
    .X(_03194_));
 sky130_fd_sc_hd__buf_4 _08409_ (.A(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__clkinv_4 _08410_ (.A(net66),
    .Y(_03196_));
 sky130_fd_sc_hd__a2111oi_1 _08411_ (.A1(prefetched_high_word),
    .A2(clear_prefetched_high_word_q),
    .B1(_03195_),
    .C1(latched_branch),
    .D1(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__and3_2 _08412_ (.A(prefetched_high_word),
    .B(_03193_),
    .C(_03197_),
    .X(_03198_));
 sky130_fd_sc_hd__buf_4 _08413_ (.A(mem_do_rinst),
    .X(_03199_));
 sky130_fd_sc_hd__a22oi_4 _08414_ (.A1(net262),
    .A2(net65),
    .B1(_03198_),
    .B2(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__mux2_1 _08415_ (.A0(net33),
    .A1(\mem_rdata_q[0] ),
    .S(_03200_),
    .X(_03201_));
 sky130_fd_sc_hd__mux2_1 _08416_ (.A0(net40),
    .A1(\mem_rdata_q[16] ),
    .S(_03200_),
    .X(_03202_));
 sky130_fd_sc_hd__clkbuf_4 _08417_ (.A(_03193_),
    .X(_03203_));
 sky130_fd_sc_hd__mux2_1 _08418_ (.A0(_03201_),
    .A1(_03202_),
    .S(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__nor2_2 _08419_ (.A(mem_la_secondword),
    .B(_03198_),
    .Y(_03205_));
 sky130_fd_sc_hd__mux2_2 _08420_ (.A0(\mem_16bit_buffer[0] ),
    .A1(_03204_),
    .S(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__a22o_1 _08421_ (.A1(net262),
    .A2(net65),
    .B1(_03198_),
    .B2(mem_do_rinst),
    .X(_03207_));
 sky130_fd_sc_hd__clkbuf_4 _08422_ (.A(_03207_),
    .X(_03208_));
 sky130_fd_sc_hd__mux2_1 _08423_ (.A0(\mem_rdata_q[1] ),
    .A1(net44),
    .S(_03208_),
    .X(_03209_));
 sky130_fd_sc_hd__mux2_1 _08424_ (.A0(\mem_rdata_q[17] ),
    .A1(net41),
    .S(_03207_),
    .X(_03210_));
 sky130_fd_sc_hd__mux2_1 _08425_ (.A0(_03209_),
    .A1(_03210_),
    .S(_03203_),
    .X(_03211_));
 sky130_fd_sc_hd__mux2_1 _08426_ (.A0(\mem_16bit_buffer[1] ),
    .A1(_03211_),
    .S(_03205_),
    .X(_03212_));
 sky130_fd_sc_hd__clkbuf_4 _08427_ (.A(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__and2_1 _08428_ (.A(_03206_),
    .B(_03213_),
    .X(_03214_));
 sky130_fd_sc_hd__clkbuf_4 _08429_ (.A(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__mux2_1 _08430_ (.A0(_03203_),
    .A1(mem_la_firstword_reg),
    .S(last_mem_valid),
    .X(_03216_));
 sky130_fd_sc_hd__and2_2 _08431_ (.A(_03207_),
    .B(_03216_),
    .X(_03217_));
 sky130_fd_sc_hd__clkbuf_4 _08432_ (.A(mem_do_rdata),
    .X(_03218_));
 sky130_fd_sc_hd__buf_4 _08433_ (.A(_03192_),
    .X(_03219_));
 sky130_fd_sc_hd__nor2_1 _08434_ (.A(\mem_state[0] ),
    .B(\mem_state[1] ),
    .Y(_03220_));
 sky130_fd_sc_hd__o21ai_2 _08435_ (.A1(_03218_),
    .A2(_03219_),
    .B1(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__nor2_1 _08436_ (.A(_03198_),
    .B(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hd__a31o_1 _08437_ (.A1(_03187_),
    .A2(_03215_),
    .A3(_03217_),
    .B1(_03222_),
    .X(_03223_));
 sky130_fd_sc_hd__and2_1 _08438_ (.A(net66),
    .B(_03223_),
    .X(_03224_));
 sky130_fd_sc_hd__clkbuf_2 _08439_ (.A(_03224_),
    .X(net224));
 sky130_fd_sc_hd__inv_2 _08440_ (.A(_03197_),
    .Y(clear_prefetched_high_word));
 sky130_fd_sc_hd__clkbuf_4 _08441_ (.A(\cpu_state[6] ),
    .X(_03225_));
 sky130_fd_sc_hd__clkbuf_4 _08442_ (.A(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__clkbuf_4 _08443_ (.A(_03208_),
    .X(_03227_));
 sky130_fd_sc_hd__nand2_2 _08444_ (.A(_03206_),
    .B(_03212_),
    .Y(_03228_));
 sky130_fd_sc_hd__nor2_2 _08445_ (.A(_03199_),
    .B(mem_do_prefetch),
    .Y(_03229_));
 sky130_fd_sc_hd__or3_2 _08446_ (.A(mem_la_secondword),
    .B(_03229_),
    .C(_03191_),
    .X(_03230_));
 sky130_fd_sc_hd__clkbuf_4 _08447_ (.A(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__a21oi_1 _08448_ (.A1(_03227_),
    .A2(_03228_),
    .B1(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__or2_1 _08449_ (.A(\mem_state[0] ),
    .B(\mem_state[1] ),
    .X(_03233_));
 sky130_fd_sc_hd__o311a_1 _08450_ (.A1(mem_do_wdata),
    .A2(mem_do_rdata),
    .A3(_03199_),
    .B1(_03227_),
    .C1(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__a31o_1 _08451_ (.A1(_03199_),
    .A2(\mem_state[0] ),
    .A3(\mem_state[1] ),
    .B1(_03234_),
    .X(_03235_));
 sky130_fd_sc_hd__or3b_1 _08452_ (.A(_03196_),
    .B(_03232_),
    .C_N(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__buf_2 _08453_ (.A(_03236_),
    .X(_03237_));
 sky130_fd_sc_hd__or2_1 _08454_ (.A(mem_do_prefetch),
    .B(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__clkbuf_8 _08455_ (.A(_03196_),
    .X(_03239_));
 sky130_fd_sc_hd__clkbuf_8 _08456_ (.A(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__and3_1 _08457_ (.A(\reg_next_pc[0] ),
    .B(_03199_),
    .C(net66),
    .X(_03241_));
 sky130_fd_sc_hd__clkbuf_4 _08458_ (.A(net78),
    .X(_03242_));
 sky130_fd_sc_hd__or2_1 _08459_ (.A(_03242_),
    .B(net67),
    .X(_03243_));
 sky130_fd_sc_hd__a22o_1 _08460_ (.A1(net67),
    .A2(\mem_wordsize[2] ),
    .B1(_03243_),
    .B2(\mem_wordsize[0] ),
    .X(_03244_));
 sky130_fd_sc_hd__or2_1 _08461_ (.A(_03241_),
    .B(_03244_),
    .X(_03245_));
 sky130_fd_sc_hd__o21ai_1 _08462_ (.A1(\irq_mask[2] ),
    .A2(irq_active),
    .B1(_03245_),
    .Y(_03246_));
 sky130_fd_sc_hd__or3_1 _08463_ (.A(mem_do_wdata),
    .B(_03218_),
    .C(_03241_),
    .X(_03247_));
 sky130_fd_sc_hd__nand2_2 _08464_ (.A(net66),
    .B(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__or2_2 _08465_ (.A(_03246_),
    .B(_03248_),
    .X(_03249_));
 sky130_fd_sc_hd__inv_2 _08466_ (.A(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__nor2_1 _08467_ (.A(_03240_),
    .B(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__or3_4 _08468_ (.A(instr_timer),
    .B(instr_maskirq),
    .C(instr_retirq),
    .X(_03252_));
 sky130_fd_sc_hd__nor3_4 _08469_ (.A(instr_rdinstrh),
    .B(instr_rdinstr),
    .C(instr_rdcycleh),
    .Y(_03253_));
 sky130_fd_sc_hd__or3b_4 _08470_ (.A(_03252_),
    .B(instr_rdcycle),
    .C_N(_03253_),
    .X(_03254_));
 sky130_fd_sc_hd__or4_2 _08471_ (.A(instr_sltu),
    .B(instr_slt),
    .C(instr_sltiu),
    .D(instr_slti),
    .X(_03255_));
 sky130_fd_sc_hd__or4_1 _08472_ (.A(instr_lh),
    .B(instr_jalr),
    .C(instr_jal),
    .D(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__or2_1 _08473_ (.A(instr_auipc),
    .B(instr_lui),
    .X(_03257_));
 sky130_fd_sc_hd__or2_1 _08474_ (.A(instr_lbu),
    .B(instr_lb),
    .X(_03258_));
 sky130_fd_sc_hd__or3_1 _08475_ (.A(instr_sw),
    .B(instr_sh),
    .C(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__or4_1 _08476_ (.A(instr_fence),
    .B(instr_and),
    .C(_03257_),
    .D(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__or4_1 _08477_ (.A(instr_sll),
    .B(instr_sub),
    .C(instr_add),
    .D(instr_andi),
    .X(_03261_));
 sky130_fd_sc_hd__or4_1 _08478_ (.A(instr_or),
    .B(instr_sra),
    .C(instr_srl),
    .D(instr_xor),
    .X(_03262_));
 sky130_fd_sc_hd__or4_1 _08479_ (.A(instr_bltu),
    .B(instr_bge),
    .C(instr_blt),
    .D(instr_bne),
    .X(_03263_));
 sky130_fd_sc_hd__or4_1 _08480_ (.A(instr_ori),
    .B(instr_xori),
    .C(instr_addi),
    .D(instr_bgeu),
    .X(_03264_));
 sky130_fd_sc_hd__or4_1 _08481_ (.A(_03261_),
    .B(_03262_),
    .C(_03263_),
    .D(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__or4_1 _08482_ (.A(instr_beq),
    .B(instr_waitirq),
    .C(instr_srai),
    .D(instr_slli),
    .X(_03266_));
 sky130_fd_sc_hd__or4_1 _08483_ (.A(instr_srli),
    .B(instr_lhu),
    .C(instr_sb),
    .D(instr_lw),
    .X(_03267_));
 sky130_fd_sc_hd__or4_1 _08484_ (.A(_03260_),
    .B(_03265_),
    .C(_03266_),
    .D(_03267_),
    .X(_03268_));
 sky130_fd_sc_hd__nor3_2 _08485_ (.A(_03254_),
    .B(_03256_),
    .C(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__inv_2 _08486_ (.A(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hd__inv_2 _08487_ (.A(\cpu_state[2] ),
    .Y(_03271_));
 sky130_fd_sc_hd__nor2_4 _08488_ (.A(_03239_),
    .B(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__and4_1 _08489_ (.A(is_lb_lh_lw_lbu_lhu),
    .B(_03270_),
    .C(_03272_),
    .D(_03249_),
    .X(_03273_));
 sky130_fd_sc_hd__a31o_1 _08490_ (.A1(_03226_),
    .A2(_03238_),
    .A3(_03251_),
    .B1(_03273_),
    .X(_00080_));
 sky130_fd_sc_hd__or2_2 _08491_ (.A(\cpu_state[6] ),
    .B(\cpu_state[5] ),
    .X(_03274_));
 sky130_fd_sc_hd__clkbuf_4 _08492_ (.A(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__buf_4 _08493_ (.A(_03275_),
    .X(_03276_));
 sky130_fd_sc_hd__buf_4 _08494_ (.A(net66),
    .X(_03277_));
 sky130_fd_sc_hd__and2_1 _08495_ (.A(mem_do_prefetch),
    .B(_03237_),
    .X(_03278_));
 sky130_fd_sc_hd__o21ai_1 _08496_ (.A1(_03218_),
    .A2(_03278_),
    .B1(\cpu_state[6] ),
    .Y(_03279_));
 sky130_fd_sc_hd__o21ai_1 _08497_ (.A1(mem_do_wdata),
    .A2(_03278_),
    .B1(\cpu_state[5] ),
    .Y(_03280_));
 sky130_fd_sc_hd__and3_1 _08498_ (.A(_03277_),
    .B(_03279_),
    .C(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__or3b_2 _08499_ (.A(_03218_),
    .B(_03278_),
    .C_N(\cpu_state[6] ),
    .X(_03282_));
 sky130_fd_sc_hd__or2_1 _08500_ (.A(instr_lhu),
    .B(instr_lh),
    .X(_03283_));
 sky130_fd_sc_hd__or2_1 _08501_ (.A(instr_lw),
    .B(_03283_),
    .X(_03284_));
 sky130_fd_sc_hd__or4_1 _08502_ (.A(_03239_),
    .B(_03258_),
    .C(_03282_),
    .D(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__inv_2 _08503_ (.A(mem_do_wdata),
    .Y(_03286_));
 sky130_fd_sc_hd__and4bb_1 _08504_ (.A_N(_03196_),
    .B_N(_03278_),
    .C(\cpu_state[5] ),
    .D(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__or4b_1 _08505_ (.A(instr_sw),
    .B(instr_sh),
    .C(instr_sb),
    .D_N(_03287_),
    .X(_03288_));
 sky130_fd_sc_hd__and3_1 _08506_ (.A(_03281_),
    .B(_03285_),
    .C(_03288_),
    .X(_03289_));
 sky130_fd_sc_hd__nand2_1 _08507_ (.A(_03276_),
    .B(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__nor2_2 _08508_ (.A(_03239_),
    .B(_03282_),
    .Y(_03291_));
 sky130_fd_sc_hd__inv_2 _08509_ (.A(\cpu_state[1] ),
    .Y(_03292_));
 sky130_fd_sc_hd__nor2_4 _08510_ (.A(_03292_),
    .B(_03196_),
    .Y(_03293_));
 sky130_fd_sc_hd__buf_4 _08511_ (.A(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__a221o_1 _08512_ (.A1(instr_lw),
    .A2(_03291_),
    .B1(_03287_),
    .B2(instr_sw),
    .C1(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__a21o_1 _08513_ (.A1(\mem_wordsize[0] ),
    .A2(_03290_),
    .B1(_03295_),
    .X(_00081_));
 sky130_fd_sc_hd__and3_1 _08514_ (.A(mem_do_wdata),
    .B(net66),
    .C(_03220_),
    .X(_03296_));
 sky130_fd_sc_hd__buf_2 _08515_ (.A(_03296_),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_4 _08516_ (.A(\mem_wordsize[2] ),
    .X(_03297_));
 sky130_fd_sc_hd__buf_4 _08517_ (.A(\cpu_state[1] ),
    .X(_03298_));
 sky130_fd_sc_hd__o21ai_2 _08518_ (.A1(_03298_),
    .A2(_03276_),
    .B1(_03289_),
    .Y(_03299_));
 sky130_fd_sc_hd__a22o_1 _08519_ (.A1(_03291_),
    .A2(_03283_),
    .B1(_03287_),
    .B2(instr_sh),
    .X(_03300_));
 sky130_fd_sc_hd__a21o_1 _08520_ (.A1(_03297_),
    .A2(_03299_),
    .B1(_03300_),
    .X(_00083_));
 sky130_fd_sc_hd__buf_4 _08521_ (.A(\cpu_state[2] ),
    .X(_03301_));
 sky130_fd_sc_hd__buf_4 _08522_ (.A(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__buf_4 _08523_ (.A(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__buf_4 _08524_ (.A(_03277_),
    .X(_03304_));
 sky130_fd_sc_hd__buf_4 _08525_ (.A(_03304_),
    .X(_03305_));
 sky130_fd_sc_hd__a21bo_1 _08526_ (.A1(_03305_),
    .A2(_03246_),
    .B1_N(_03247_),
    .X(_03306_));
 sky130_fd_sc_hd__nand2_1 _08527_ (.A(\cpu_state[2] ),
    .B(_03269_),
    .Y(_03307_));
 sky130_fd_sc_hd__nor3_4 _08528_ (.A(\irq_mask[1] ),
    .B(irq_active),
    .C(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__buf_4 _08529_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_03309_));
 sky130_fd_sc_hd__inv_2 _08530_ (.A(_03237_),
    .Y(_03310_));
 sky130_fd_sc_hd__nor2_4 _08531_ (.A(\cpu_state[6] ),
    .B(\cpu_state[5] ),
    .Y(_03311_));
 sky130_fd_sc_hd__nor2_1 _08532_ (.A(_03238_),
    .B(_03311_),
    .Y(_01226_));
 sky130_fd_sc_hd__clkbuf_4 _08533_ (.A(\cpu_state[4] ),
    .X(_03312_));
 sky130_fd_sc_hd__nor3_2 _08534_ (.A(\reg_sh[4] ),
    .B(\reg_sh[3] ),
    .C(\reg_sh[2] ),
    .Y(_03313_));
 sky130_fd_sc_hd__nand2_1 _08535_ (.A(_03312_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__or2_2 _08536_ (.A(\reg_sh[1] ),
    .B(\reg_sh[0] ),
    .X(_03315_));
 sky130_fd_sc_hd__nor2_1 _08537_ (.A(_03314_),
    .B(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__inv_2 _08538_ (.A(\cpu_state[3] ),
    .Y(_03317_));
 sky130_fd_sc_hd__nor2_1 _08539_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(_03317_),
    .Y(_03318_));
 sky130_fd_sc_hd__o21a_2 _08540_ (.A1(decoder_trigger),
    .A2(do_waitirq),
    .B1(instr_waitirq),
    .X(_03319_));
 sky130_fd_sc_hd__and2b_2 _08541_ (.A_N(\irq_mask[22] ),
    .B(\irq_pending[22] ),
    .X(_03320_));
 sky130_fd_sc_hd__and2b_2 _08542_ (.A_N(\irq_mask[6] ),
    .B(\irq_pending[6] ),
    .X(_03321_));
 sky130_fd_sc_hd__and2b_2 _08543_ (.A_N(\irq_mask[5] ),
    .B(\irq_pending[5] ),
    .X(_03322_));
 sky130_fd_sc_hd__and2b_2 _08544_ (.A_N(\irq_mask[9] ),
    .B(\irq_pending[9] ),
    .X(_03323_));
 sky130_fd_sc_hd__or4_1 _08545_ (.A(_03320_),
    .B(_03321_),
    .C(_03322_),
    .D(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__and2b_1 _08546_ (.A_N(\irq_mask[26] ),
    .B(\irq_pending[26] ),
    .X(_03325_));
 sky130_fd_sc_hd__and2b_2 _08547_ (.A_N(\irq_mask[2] ),
    .B(\irq_pending[2] ),
    .X(_03326_));
 sky130_fd_sc_hd__and2b_4 _08548_ (.A_N(\irq_mask[4] ),
    .B(\irq_pending[4] ),
    .X(_03327_));
 sky130_fd_sc_hd__and2b_1 _08549_ (.A_N(\irq_mask[30] ),
    .B(\irq_pending[30] ),
    .X(_03328_));
 sky130_fd_sc_hd__or4_1 _08550_ (.A(_03325_),
    .B(_03326_),
    .C(_03327_),
    .D(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__and2b_2 _08551_ (.A_N(\irq_mask[16] ),
    .B(\irq_pending[16] ),
    .X(_03330_));
 sky130_fd_sc_hd__and2b_1 _08552_ (.A_N(\irq_mask[31] ),
    .B(\irq_pending[31] ),
    .X(_03331_));
 sky130_fd_sc_hd__and2b_1 _08553_ (.A_N(\irq_mask[20] ),
    .B(\irq_pending[20] ),
    .X(_03332_));
 sky130_fd_sc_hd__and2b_2 _08554_ (.A_N(\irq_mask[10] ),
    .B(\irq_pending[10] ),
    .X(_03333_));
 sky130_fd_sc_hd__or4_1 _08555_ (.A(_03330_),
    .B(_03331_),
    .C(_03332_),
    .D(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__and2b_2 _08556_ (.A_N(\irq_mask[11] ),
    .B(\irq_pending[11] ),
    .X(_03335_));
 sky130_fd_sc_hd__and2b_2 _08557_ (.A_N(\irq_mask[18] ),
    .B(\irq_pending[18] ),
    .X(_03336_));
 sky130_fd_sc_hd__and2b_1 _08558_ (.A_N(\irq_mask[29] ),
    .B(\irq_pending[29] ),
    .X(_03337_));
 sky130_fd_sc_hd__and2b_2 _08559_ (.A_N(\irq_mask[0] ),
    .B(\irq_pending[0] ),
    .X(_03338_));
 sky130_fd_sc_hd__or4_1 _08560_ (.A(_03335_),
    .B(_03336_),
    .C(_03337_),
    .D(_03338_),
    .X(_03339_));
 sky130_fd_sc_hd__or4_4 _08561_ (.A(_03324_),
    .B(_03329_),
    .C(_03334_),
    .D(_03339_),
    .X(_03340_));
 sky130_fd_sc_hd__and2b_1 _08562_ (.A_N(\irq_mask[27] ),
    .B(\irq_pending[27] ),
    .X(_03341_));
 sky130_fd_sc_hd__and2b_1 _08563_ (.A_N(\irq_mask[24] ),
    .B(\irq_pending[24] ),
    .X(_03342_));
 sky130_fd_sc_hd__and2b_1 _08564_ (.A_N(\irq_mask[23] ),
    .B(\irq_pending[23] ),
    .X(_03343_));
 sky130_fd_sc_hd__and2b_2 _08565_ (.A_N(\irq_mask[3] ),
    .B(\irq_pending[3] ),
    .X(_03344_));
 sky130_fd_sc_hd__or4_1 _08566_ (.A(_03341_),
    .B(_03342_),
    .C(_03343_),
    .D(_03344_),
    .X(_03345_));
 sky130_fd_sc_hd__and2b_1 _08567_ (.A_N(\irq_mask[21] ),
    .B(\irq_pending[21] ),
    .X(_03346_));
 sky130_fd_sc_hd__and2b_1 _08568_ (.A_N(\irq_mask[25] ),
    .B(\irq_pending[25] ),
    .X(_03347_));
 sky130_fd_sc_hd__and2b_2 _08569_ (.A_N(\irq_mask[17] ),
    .B(\irq_pending[17] ),
    .X(_03348_));
 sky130_fd_sc_hd__and2b_2 _08570_ (.A_N(\irq_mask[7] ),
    .B(\irq_pending[7] ),
    .X(_03349_));
 sky130_fd_sc_hd__or4_1 _08571_ (.A(_03346_),
    .B(_03347_),
    .C(_03348_),
    .D(_03349_),
    .X(_03350_));
 sky130_fd_sc_hd__and2b_2 _08572_ (.A_N(\irq_mask[1] ),
    .B(\irq_pending[1] ),
    .X(_03351_));
 sky130_fd_sc_hd__and2b_2 _08573_ (.A_N(\irq_mask[13] ),
    .B(\irq_pending[13] ),
    .X(_03352_));
 sky130_fd_sc_hd__and2b_2 _08574_ (.A_N(\irq_mask[14] ),
    .B(\irq_pending[14] ),
    .X(_03353_));
 sky130_fd_sc_hd__and2b_1 _08575_ (.A_N(\irq_mask[28] ),
    .B(\irq_pending[28] ),
    .X(_03354_));
 sky130_fd_sc_hd__or4_1 _08576_ (.A(_03351_),
    .B(_03352_),
    .C(_03353_),
    .D(_03354_),
    .X(_03355_));
 sky130_fd_sc_hd__and2b_2 _08577_ (.A_N(\irq_mask[15] ),
    .B(\irq_pending[15] ),
    .X(_03356_));
 sky130_fd_sc_hd__and2b_2 _08578_ (.A_N(\irq_mask[12] ),
    .B(\irq_pending[12] ),
    .X(_03357_));
 sky130_fd_sc_hd__and2b_2 _08579_ (.A_N(\irq_mask[19] ),
    .B(\irq_pending[19] ),
    .X(_03358_));
 sky130_fd_sc_hd__and2b_2 _08580_ (.A_N(\irq_mask[8] ),
    .B(\irq_pending[8] ),
    .X(_03359_));
 sky130_fd_sc_hd__or4_1 _08581_ (.A(_03356_),
    .B(_03357_),
    .C(_03358_),
    .D(_03359_),
    .X(_03360_));
 sky130_fd_sc_hd__or4_2 _08582_ (.A(_03345_),
    .B(_03350_),
    .C(_03355_),
    .D(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__nor2_1 _08583_ (.A(irq_active),
    .B(irq_delay),
    .Y(_03362_));
 sky130_fd_sc_hd__o211a_2 _08584_ (.A1(_03340_),
    .A2(_03361_),
    .B1(_03362_),
    .C1(decoder_trigger),
    .X(_03363_));
 sky130_fd_sc_hd__nor2_4 _08585_ (.A(_03195_),
    .B(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__a31o_1 _08586_ (.A1(_03298_),
    .A2(_03319_),
    .A3(_03364_),
    .B1(_03308_),
    .X(_03365_));
 sky130_fd_sc_hd__inv_2 _08587_ (.A(instr_jal),
    .Y(_03366_));
 sky130_fd_sc_hd__or2b_2 _08588_ (.A(instr_waitirq),
    .B_N(decoder_trigger),
    .X(_03367_));
 sky130_fd_sc_hd__nor2_4 _08589_ (.A(_03366_),
    .B(_03367_),
    .Y(_03368_));
 sky130_fd_sc_hd__o21ai_1 _08590_ (.A1(decoder_trigger),
    .A2(do_waitirq),
    .B1(instr_waitirq),
    .Y(_03369_));
 sky130_fd_sc_hd__o211a_1 _08591_ (.A1(_03248_),
    .A2(_03369_),
    .B1(_03367_),
    .C1(_03249_),
    .X(_03370_));
 sky130_fd_sc_hd__or3b_1 _08592_ (.A(_03368_),
    .B(_03370_),
    .C_N(_03364_),
    .X(_03371_));
 sky130_fd_sc_hd__a32o_1 _08593_ (.A1(_03277_),
    .A2(_03247_),
    .A3(_03365_),
    .B1(_03371_),
    .B2(_03298_),
    .X(_03372_));
 sky130_fd_sc_hd__or4_1 _08594_ (.A(_03196_),
    .B(_03316_),
    .C(_03318_),
    .D(_03372_),
    .X(_03373_));
 sky130_fd_sc_hd__a311o_1 _08595_ (.A1(_03309_),
    .A2(\cpu_state[3] ),
    .A3(_03310_),
    .B1(_01226_),
    .C1(_03373_),
    .X(_03374_));
 sky130_fd_sc_hd__a22o_1 _08596_ (.A1(_03248_),
    .A2(_03308_),
    .B1(_03374_),
    .B2(_03249_),
    .X(_03375_));
 sky130_fd_sc_hd__a31o_1 _08597_ (.A1(_03303_),
    .A2(_03254_),
    .A3(_03306_),
    .B1(_03375_),
    .X(_00075_));
 sky130_fd_sc_hd__nor2_1 _08598_ (.A(\irq_state[1] ),
    .B(\irq_state[0] ),
    .Y(_03376_));
 sky130_fd_sc_hd__and3b_1 _08599_ (.A_N(_03363_),
    .B(_03293_),
    .C(_03376_),
    .X(_03377_));
 sky130_fd_sc_hd__buf_2 _08600_ (.A(_03377_),
    .X(_03378_));
 sky130_fd_sc_hd__nor2_2 _08601_ (.A(instr_jal),
    .B(_03367_),
    .Y(_03379_));
 sky130_fd_sc_hd__nand2_1 _08602_ (.A(_03378_),
    .B(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__nor2_1 _08603_ (.A(_03250_),
    .B(_03380_),
    .Y(_00076_));
 sky130_fd_sc_hd__o211a_1 _08604_ (.A1(\irq_mask[1] ),
    .A2(irq_active),
    .B1(_03269_),
    .C1(_03272_),
    .X(_03381_));
 sky130_fd_sc_hd__and2_1 _08605_ (.A(_03277_),
    .B(\cpu_state[0] ),
    .X(_03382_));
 sky130_fd_sc_hd__buf_1 _08606_ (.A(_03382_),
    .X(_00865_));
 sky130_fd_sc_hd__or3_1 _08607_ (.A(_03250_),
    .B(_03381_),
    .C(_00865_),
    .X(_03383_));
 sky130_fd_sc_hd__clkbuf_1 _08608_ (.A(_03383_),
    .X(_00074_));
 sky130_fd_sc_hd__buf_4 _08609_ (.A(\cpu_state[3] ),
    .X(_03384_));
 sky130_fd_sc_hd__buf_4 _08610_ (.A(_03384_),
    .X(_03385_));
 sky130_fd_sc_hd__nand2_1 _08611_ (.A(_03277_),
    .B(_03249_),
    .Y(_03386_));
 sky130_fd_sc_hd__clkbuf_4 _08612_ (.A(is_lui_auipc_jal),
    .X(_03387_));
 sky130_fd_sc_hd__or3_1 _08613_ (.A(is_slli_srli_srai),
    .B(_03387_),
    .C(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .X(_03388_));
 sky130_fd_sc_hd__or2_1 _08614_ (.A(_03271_),
    .B(_03254_),
    .X(_03389_));
 sky130_fd_sc_hd__or4_1 _08615_ (.A(is_lb_lh_lw_lbu_lhu),
    .B(_03269_),
    .C(_03388_),
    .D(_03389_),
    .X(_03390_));
 sky130_fd_sc_hd__or2_1 _08616_ (.A(_03386_),
    .B(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__o21a_1 _08617_ (.A1(\irq_mask[2] ),
    .A2(irq_active),
    .B1(_03241_),
    .X(_03392_));
 sky130_fd_sc_hd__o21ai_1 _08618_ (.A1(mem_do_wdata),
    .A2(_03218_),
    .B1(_03244_),
    .Y(_03393_));
 sky130_fd_sc_hd__nor4b_4 _08619_ (.A(\irq_mask[2] ),
    .B(irq_active),
    .C(_03248_),
    .D_N(_03245_),
    .Y(_03394_));
 sky130_fd_sc_hd__a21oi_1 _08620_ (.A1(_03304_),
    .A2(_03393_),
    .B1(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__nor3_2 _08621_ (.A(is_slli_srli_srai),
    .B(_03387_),
    .C(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .Y(_03396_));
 sky130_fd_sc_hd__or4_1 _08622_ (.A(_03271_),
    .B(_03392_),
    .C(_03395_),
    .D(_03396_),
    .X(_03397_));
 sky130_fd_sc_hd__o21ai_1 _08623_ (.A1(is_sb_sh_sw),
    .A2(_03391_),
    .B1(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__a41o_1 _08624_ (.A1(_03309_),
    .A2(_03385_),
    .A3(_03237_),
    .A4(_03251_),
    .B1(_03398_),
    .X(_00077_));
 sky130_fd_sc_hd__or3_4 _08625_ (.A(\reg_sh[4] ),
    .B(\reg_sh[3] ),
    .C(\reg_sh[2] ),
    .X(_03399_));
 sky130_fd_sc_hd__o21ai_4 _08626_ (.A1(_03399_),
    .A2(_03315_),
    .B1(_03312_),
    .Y(_03400_));
 sky130_fd_sc_hd__nor2_1 _08627_ (.A(_03386_),
    .B(_03400_),
    .Y(_00078_));
 sky130_fd_sc_hd__inv_2 _08628_ (.A(_03391_),
    .Y(_03401_));
 sky130_fd_sc_hd__a32o_1 _08629_ (.A1(\cpu_state[5] ),
    .A2(_03238_),
    .A3(_03251_),
    .B1(_03401_),
    .B2(is_sb_sh_sw),
    .X(_00079_));
 sky130_fd_sc_hd__buf_2 _08630_ (.A(instr_jal),
    .X(_03402_));
 sky130_fd_sc_hd__buf_2 _08631_ (.A(_03257_),
    .X(_03403_));
 sky130_fd_sc_hd__or2_1 _08632_ (.A(_03402_),
    .B(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__clkbuf_1 _08633_ (.A(_03404_),
    .X(_00033_));
 sky130_fd_sc_hd__or3_1 _08634_ (.A(instr_slt),
    .B(instr_slti),
    .C(instr_blt),
    .X(_03405_));
 sky130_fd_sc_hd__clkbuf_1 _08635_ (.A(_03405_),
    .X(_00034_));
 sky130_fd_sc_hd__or3_1 _08636_ (.A(instr_sltu),
    .B(instr_sltiu),
    .C(instr_bltu),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_1 _08637_ (.A(_03406_),
    .X(_00035_));
 sky130_fd_sc_hd__clkbuf_4 _08638_ (.A(\mem_wordsize[1] ),
    .X(_03407_));
 sky130_fd_sc_hd__a22o_1 _08639_ (.A1(_03258_),
    .A2(_03291_),
    .B1(_03287_),
    .B2(instr_sb),
    .X(_03408_));
 sky130_fd_sc_hd__a21o_1 _08640_ (.A1(_03407_),
    .A2(_03299_),
    .B1(_03408_),
    .X(_00082_));
 sky130_fd_sc_hd__clkbuf_4 _08641_ (.A(\irq_state[1] ),
    .X(_03409_));
 sky130_fd_sc_hd__or2_4 _08642_ (.A(\cpu_state[2] ),
    .B(\cpu_state[4] ),
    .X(_03410_));
 sky130_fd_sc_hd__nor3_2 _08643_ (.A(\cpu_state[0] ),
    .B(_03274_),
    .C(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__nand3_2 _08644_ (.A(_03317_),
    .B(_03409_),
    .C(_03411_),
    .Y(_03412_));
 sky130_fd_sc_hd__o211a_1 _08645_ (.A1(\irq_mask[2] ),
    .A2(_03412_),
    .B1(\irq_pending[2] ),
    .C1(_03304_),
    .X(_03413_));
 sky130_fd_sc_hd__or3_1 _08646_ (.A(net23),
    .B(_03394_),
    .C(_03413_),
    .X(_03414_));
 sky130_fd_sc_hd__clkbuf_1 _08647_ (.A(_03414_),
    .X(_00023_));
 sky130_fd_sc_hd__or4_1 _08648_ (.A(\timer[5] ),
    .B(\timer[6] ),
    .C(\timer[1] ),
    .D(\timer[2] ),
    .X(_03415_));
 sky130_fd_sc_hd__or4_1 _08649_ (.A(\timer[4] ),
    .B(\timer[7] ),
    .C(\timer[3] ),
    .D(_03415_),
    .X(_03416_));
 sky130_fd_sc_hd__or4_1 _08650_ (.A(\timer[25] ),
    .B(\timer[24] ),
    .C(\timer[27] ),
    .D(\timer[26] ),
    .X(_03417_));
 sky130_fd_sc_hd__or4_1 _08651_ (.A(\timer[21] ),
    .B(\timer[20] ),
    .C(\timer[23] ),
    .D(\timer[22] ),
    .X(_03418_));
 sky130_fd_sc_hd__or4_1 _08652_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .C(\timer[15] ),
    .D(\timer[14] ),
    .X(_03419_));
 sky130_fd_sc_hd__or4_1 _08653_ (.A(\timer[17] ),
    .B(\timer[16] ),
    .C(\timer[19] ),
    .D(\timer[18] ),
    .X(_03420_));
 sky130_fd_sc_hd__or3_1 _08654_ (.A(_03418_),
    .B(_03419_),
    .C(_03420_),
    .X(_03421_));
 sky130_fd_sc_hd__or3_1 _08655_ (.A(\timer[9] ),
    .B(\timer[11] ),
    .C(\timer[10] ),
    .X(_03422_));
 sky130_fd_sc_hd__or4_1 _08656_ (.A(\timer[8] ),
    .B(_03417_),
    .C(_03421_),
    .D(_03422_),
    .X(_03423_));
 sky130_fd_sc_hd__or3_1 _08657_ (.A(\timer[29] ),
    .B(\timer[28] ),
    .C(\timer[30] ),
    .X(_03424_));
 sky130_fd_sc_hd__nor2_1 _08658_ (.A(\timer[31] ),
    .B(_03424_),
    .Y(_03425_));
 sky130_fd_sc_hd__or3b_1 _08659_ (.A(_03416_),
    .B(_03423_),
    .C_N(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__inv_2 _08660_ (.A(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__buf_2 _08661_ (.A(_03412_),
    .X(_03428_));
 sky130_fd_sc_hd__o211a_1 _08662_ (.A1(\irq_mask[0] ),
    .A2(_03428_),
    .B1(\irq_pending[0] ),
    .C1(_03305_),
    .X(_03429_));
 sky130_fd_sc_hd__a211o_1 _08663_ (.A1(\timer[0] ),
    .A2(_03427_),
    .B1(_03429_),
    .C1(net1),
    .X(_00001_));
 sky130_fd_sc_hd__or3_1 _08664_ (.A(instr_bgeu),
    .B(instr_bge),
    .C(instr_bne),
    .X(_03430_));
 sky130_fd_sc_hd__nor2_1 _08665_ (.A(instr_beq),
    .B(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__or2_1 _08666_ (.A(net91),
    .B(net123),
    .X(_03432_));
 sky130_fd_sc_hd__nand2_1 _08667_ (.A(net91),
    .B(net123),
    .Y(_03433_));
 sky130_fd_sc_hd__nand2_2 _08668_ (.A(_03432_),
    .B(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__nor2_1 _08669_ (.A(net122),
    .B(net90),
    .Y(_03435_));
 sky130_fd_sc_hd__and2_1 _08670_ (.A(net122),
    .B(net90),
    .X(_03436_));
 sky130_fd_sc_hd__or2_1 _08671_ (.A(_03435_),
    .B(_03436_),
    .X(_03437_));
 sky130_fd_sc_hd__clkbuf_2 _08672_ (.A(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__nand2_1 _08673_ (.A(_03434_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__nor2_1 _08674_ (.A(net119),
    .B(net87),
    .Y(_03440_));
 sky130_fd_sc_hd__nand2_1 _08675_ (.A(net119),
    .B(net87),
    .Y(_03441_));
 sky130_fd_sc_hd__and2b_1 _08676_ (.A_N(_03440_),
    .B(_03441_),
    .X(_03442_));
 sky130_fd_sc_hd__or2_1 _08677_ (.A(net120),
    .B(net88),
    .X(_03443_));
 sky130_fd_sc_hd__nand2_2 _08678_ (.A(net120),
    .B(net88),
    .Y(_03444_));
 sky130_fd_sc_hd__nand2_1 _08679_ (.A(_03443_),
    .B(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__or3b_1 _08680_ (.A(_03439_),
    .B(_03442_),
    .C_N(_03445_),
    .X(_03446_));
 sky130_fd_sc_hd__nor2_1 _08681_ (.A(net118),
    .B(net86),
    .Y(_03447_));
 sky130_fd_sc_hd__nand2_1 _08682_ (.A(net118),
    .B(net86),
    .Y(_03448_));
 sky130_fd_sc_hd__nand2b_2 _08683_ (.A_N(_03447_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__nor2_1 _08684_ (.A(net117),
    .B(net85),
    .Y(_03450_));
 sky130_fd_sc_hd__nand2_1 _08685_ (.A(net117),
    .B(net85),
    .Y(_03451_));
 sky130_fd_sc_hd__nand2b_2 _08686_ (.A_N(_03450_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__nand2_1 _08687_ (.A(_03449_),
    .B(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__and2_1 _08688_ (.A(net116),
    .B(net84),
    .X(_03454_));
 sky130_fd_sc_hd__nor2_1 _08689_ (.A(net116),
    .B(net84),
    .Y(_03455_));
 sky130_fd_sc_hd__nor2_2 _08690_ (.A(_03454_),
    .B(_03455_),
    .Y(_03456_));
 sky130_fd_sc_hd__nor2_1 _08691_ (.A(net115),
    .B(net83),
    .Y(_03457_));
 sky130_fd_sc_hd__and2_1 _08692_ (.A(net115),
    .B(net83),
    .X(_03458_));
 sky130_fd_sc_hd__nor2_1 _08693_ (.A(_03457_),
    .B(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__inv_2 _08694_ (.A(net82),
    .Y(_03460_));
 sky130_fd_sc_hd__or2_1 _08695_ (.A(net112),
    .B(net80),
    .X(_03461_));
 sky130_fd_sc_hd__nand2_1 _08696_ (.A(net112),
    .B(net80),
    .Y(_03462_));
 sky130_fd_sc_hd__and2_1 _08697_ (.A(_03461_),
    .B(_03462_),
    .X(_03463_));
 sky130_fd_sc_hd__nor2_1 _08698_ (.A(net111),
    .B(net79),
    .Y(_03464_));
 sky130_fd_sc_hd__nand2_1 _08699_ (.A(net111),
    .B(net79),
    .Y(_03465_));
 sky130_fd_sc_hd__and2b_1 _08700_ (.A_N(_03464_),
    .B(_03465_),
    .X(_03466_));
 sky130_fd_sc_hd__or2_1 _08701_ (.A(net114),
    .B(net82),
    .X(_03467_));
 sky130_fd_sc_hd__nand2_1 _08702_ (.A(net114),
    .B(net82),
    .Y(_03468_));
 sky130_fd_sc_hd__and2_1 _08703_ (.A(_03467_),
    .B(_03468_),
    .X(_03469_));
 sky130_fd_sc_hd__or2_1 _08704_ (.A(net113),
    .B(net81),
    .X(_03470_));
 sky130_fd_sc_hd__nand2_1 _08705_ (.A(net113),
    .B(net81),
    .Y(_03471_));
 sky130_fd_sc_hd__nand2_1 _08706_ (.A(_03470_),
    .B(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__inv_2 _08707_ (.A(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__or4_1 _08708_ (.A(_03463_),
    .B(_03466_),
    .C(_03469_),
    .D(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__inv_2 _08709_ (.A(net77),
    .Y(_03475_));
 sky130_fd_sc_hd__nor2_1 _08710_ (.A(net109),
    .B(net77),
    .Y(_03476_));
 sky130_fd_sc_hd__nand2_1 _08711_ (.A(net109),
    .B(net77),
    .Y(_03477_));
 sky130_fd_sc_hd__or2b_1 _08712_ (.A(_03476_),
    .B_N(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__inv_2 _08713_ (.A(_03478_),
    .Y(_03479_));
 sky130_fd_sc_hd__or2_1 _08714_ (.A(net108),
    .B(net76),
    .X(_03480_));
 sky130_fd_sc_hd__nand2_1 _08715_ (.A(net108),
    .B(net76),
    .Y(_03481_));
 sky130_fd_sc_hd__and2_1 _08716_ (.A(_03480_),
    .B(_03481_),
    .X(_03482_));
 sky130_fd_sc_hd__or2_1 _08717_ (.A(net106),
    .B(net74),
    .X(_03483_));
 sky130_fd_sc_hd__nand2_1 _08718_ (.A(net106),
    .B(net74),
    .Y(_03484_));
 sky130_fd_sc_hd__and2_1 _08719_ (.A(_03483_),
    .B(_03484_),
    .X(_03485_));
 sky130_fd_sc_hd__nor2_1 _08720_ (.A(net107),
    .B(net75),
    .Y(_03486_));
 sky130_fd_sc_hd__and2_1 _08721_ (.A(net107),
    .B(net75),
    .X(_03487_));
 sky130_fd_sc_hd__nor2_2 _08722_ (.A(_03486_),
    .B(_03487_),
    .Y(_03488_));
 sky130_fd_sc_hd__or4_1 _08723_ (.A(_03479_),
    .B(_03482_),
    .C(_03485_),
    .D(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__or2b_1 _08724_ (.A(net73),
    .B_N(net105),
    .X(_03490_));
 sky130_fd_sc_hd__nor2_1 _08725_ (.A(net104),
    .B(net72),
    .Y(_03491_));
 sky130_fd_sc_hd__nand2_1 _08726_ (.A(net104),
    .B(net72),
    .Y(_03492_));
 sky130_fd_sc_hd__or2b_2 _08727_ (.A(_03491_),
    .B_N(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__nor2_1 _08728_ (.A(net103),
    .B(net71),
    .Y(_03494_));
 sky130_fd_sc_hd__nand2_1 _08729_ (.A(net103),
    .B(net71),
    .Y(_03495_));
 sky130_fd_sc_hd__or2b_2 _08730_ (.A(_03494_),
    .B_N(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__nor2_1 _08731_ (.A(net102),
    .B(net70),
    .Y(_03497_));
 sky130_fd_sc_hd__nand2_1 _08732_ (.A(net102),
    .B(net70),
    .Y(_03498_));
 sky130_fd_sc_hd__nand2b_2 _08733_ (.A_N(_03497_),
    .B(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hd__inv_2 _08734_ (.A(net101),
    .Y(_03500_));
 sky130_fd_sc_hd__nand2_2 _08735_ (.A(net101),
    .B(net69),
    .Y(_03501_));
 sky130_fd_sc_hd__inv_2 _08736_ (.A(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__nor2_1 _08737_ (.A(net101),
    .B(net69),
    .Y(_03503_));
 sky130_fd_sc_hd__nor2_2 _08738_ (.A(_03502_),
    .B(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__nor2_1 _08739_ (.A(net100),
    .B(net68),
    .Y(_03505_));
 sky130_fd_sc_hd__nand2_1 _08740_ (.A(net100),
    .B(net68),
    .Y(_03506_));
 sky130_fd_sc_hd__nor2b_2 _08741_ (.A(_03505_),
    .B_N(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__inv_2 _08742_ (.A(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__or2_2 _08743_ (.A(net129),
    .B(net97),
    .X(_03509_));
 sky130_fd_sc_hd__clkbuf_4 _08744_ (.A(net97),
    .X(_03510_));
 sky130_fd_sc_hd__nand2_1 _08745_ (.A(net129),
    .B(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__nand2_2 _08746_ (.A(_03509_),
    .B(_03511_),
    .Y(_03512_));
 sky130_fd_sc_hd__nor2_1 _08747_ (.A(net130),
    .B(net98),
    .Y(_03513_));
 sky130_fd_sc_hd__nand2_1 _08748_ (.A(net130),
    .B(net98),
    .Y(_03514_));
 sky130_fd_sc_hd__nand2b_2 _08749_ (.A_N(_03513_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__and4b_1 _08750_ (.A_N(_03504_),
    .B(_03508_),
    .C(_03512_),
    .D(_03515_),
    .X(_03516_));
 sky130_fd_sc_hd__inv_2 _08751_ (.A(net128),
    .Y(_03517_));
 sky130_fd_sc_hd__clkbuf_4 _08752_ (.A(net96),
    .X(_03518_));
 sky130_fd_sc_hd__nor2_1 _08753_ (.A(net127),
    .B(net95),
    .Y(_03519_));
 sky130_fd_sc_hd__nand2_1 _08754_ (.A(net127),
    .B(net95),
    .Y(_03520_));
 sky130_fd_sc_hd__and2b_1 _08755_ (.A_N(_03519_),
    .B(_03520_),
    .X(_03521_));
 sky130_fd_sc_hd__inv_2 _08756_ (.A(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__or2_1 _08757_ (.A(net126),
    .B(net94),
    .X(_03523_));
 sky130_fd_sc_hd__clkbuf_4 _08758_ (.A(net94),
    .X(_03524_));
 sky130_fd_sc_hd__nand2_1 _08759_ (.A(net126),
    .B(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__and2_1 _08760_ (.A(_03523_),
    .B(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__nor2_1 _08761_ (.A(net125),
    .B(net93),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_1 _08762_ (.A(net125),
    .B(net93),
    .Y(_03528_));
 sky130_fd_sc_hd__nand2b_2 _08763_ (.A_N(_03527_),
    .B(_03528_),
    .Y(_03529_));
 sky130_fd_sc_hd__clkbuf_4 _08764_ (.A(net124),
    .X(_03530_));
 sky130_fd_sc_hd__inv_2 _08765_ (.A(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__or2_2 _08766_ (.A(net121),
    .B(net89),
    .X(_03532_));
 sky130_fd_sc_hd__nand2_1 _08767_ (.A(net121),
    .B(net89),
    .Y(_03533_));
 sky130_fd_sc_hd__nand2_2 _08768_ (.A(_03532_),
    .B(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__xor2_2 _08769_ (.A(net78),
    .B(net110),
    .X(_03535_));
 sky130_fd_sc_hd__and2b_1 _08770_ (.A_N(net67),
    .B(net99),
    .X(_03536_));
 sky130_fd_sc_hd__or2b_1 _08771_ (.A(net110),
    .B_N(net78),
    .X(_03537_));
 sky130_fd_sc_hd__o21ai_1 _08772_ (.A1(_03535_),
    .A2(_03536_),
    .B1(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__and2b_1 _08773_ (.A_N(net121),
    .B(net89),
    .X(_03539_));
 sky130_fd_sc_hd__a21oi_1 _08774_ (.A1(_03534_),
    .A2(_03538_),
    .B1(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__o21ba_1 _08775_ (.A1(_03531_),
    .A2(net92),
    .B1_N(_03540_),
    .X(_03541_));
 sky130_fd_sc_hd__a21o_1 _08776_ (.A1(_03531_),
    .A2(net92),
    .B1(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__and2b_1 _08777_ (.A_N(net125),
    .B(net93),
    .X(_03543_));
 sky130_fd_sc_hd__a21oi_1 _08778_ (.A1(_03529_),
    .A2(_03542_),
    .B1(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__or2b_1 _08779_ (.A(net126),
    .B_N(_03524_),
    .X(_03545_));
 sky130_fd_sc_hd__o21ai_2 _08780_ (.A1(_03526_),
    .A2(_03544_),
    .B1(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__and2b_1 _08781_ (.A_N(net127),
    .B(net95),
    .X(_03547_));
 sky130_fd_sc_hd__a221o_1 _08782_ (.A1(_03517_),
    .A2(_03518_),
    .B1(_03522_),
    .B2(_03546_),
    .C1(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__o21a_1 _08783_ (.A1(_03517_),
    .A2(_03518_),
    .B1(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__inv_2 _08784_ (.A(net129),
    .Y(_03550_));
 sky130_fd_sc_hd__and2b_1 _08785_ (.A_N(net130),
    .B(net98),
    .X(_03551_));
 sky130_fd_sc_hd__a31o_1 _08786_ (.A1(_03550_),
    .A2(_03510_),
    .A3(_03515_),
    .B1(_03551_),
    .X(_03552_));
 sky130_fd_sc_hd__and2b_1 _08787_ (.A_N(net100),
    .B(net68),
    .X(_03553_));
 sky130_fd_sc_hd__a21oi_1 _08788_ (.A1(_03508_),
    .A2(_03552_),
    .B1(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__nor2_1 _08789_ (.A(_03504_),
    .B(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__a221o_1 _08790_ (.A1(_03500_),
    .A2(net69),
    .B1(_03516_),
    .B2(_03549_),
    .C1(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__and2b_1 _08791_ (.A_N(net102),
    .B(net70),
    .X(_03557_));
 sky130_fd_sc_hd__and2b_1 _08792_ (.A_N(net103),
    .B(net71),
    .X(_03558_));
 sky130_fd_sc_hd__a21o_1 _08793_ (.A1(_03496_),
    .A2(_03557_),
    .B1(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__a31o_1 _08794_ (.A1(_03496_),
    .A2(_03499_),
    .A3(_03556_),
    .B1(_03559_),
    .X(_03560_));
 sky130_fd_sc_hd__and2b_1 _08795_ (.A_N(net104),
    .B(net72),
    .X(_03561_));
 sky130_fd_sc_hd__a21o_1 _08796_ (.A1(_03493_),
    .A2(_03560_),
    .B1(_03561_),
    .X(_03562_));
 sky130_fd_sc_hd__and2b_1 _08797_ (.A_N(net105),
    .B(net73),
    .X(_03563_));
 sky130_fd_sc_hd__a21oi_2 _08798_ (.A1(_03490_),
    .A2(_03562_),
    .B1(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__or2b_1 _08799_ (.A(net106),
    .B_N(net74),
    .X(_03565_));
 sky130_fd_sc_hd__inv_2 _08800_ (.A(net75),
    .Y(_03566_));
 sky130_fd_sc_hd__or2_1 _08801_ (.A(net107),
    .B(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__o21a_1 _08802_ (.A1(_03488_),
    .A2(_03565_),
    .B1(_03567_),
    .X(_03568_));
 sky130_fd_sc_hd__or2b_1 _08803_ (.A(net108),
    .B_N(net76),
    .X(_03569_));
 sky130_fd_sc_hd__o21ai_1 _08804_ (.A1(_03482_),
    .A2(_03568_),
    .B1(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__nand2_1 _08805_ (.A(_03478_),
    .B(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__o221a_1 _08806_ (.A1(net109),
    .A2(_03475_),
    .B1(_03489_),
    .B2(_03564_),
    .C1(_03571_),
    .X(_03572_));
 sky130_fd_sc_hd__inv_2 _08807_ (.A(net111),
    .Y(_03573_));
 sky130_fd_sc_hd__nand2_1 _08808_ (.A(_03461_),
    .B(_03462_),
    .Y(_03574_));
 sky130_fd_sc_hd__inv_2 _08809_ (.A(net80),
    .Y(_03575_));
 sky130_fd_sc_hd__nor2_1 _08810_ (.A(net112),
    .B(_03575_),
    .Y(_03576_));
 sky130_fd_sc_hd__a31o_1 _08811_ (.A1(_03573_),
    .A2(net79),
    .A3(_03574_),
    .B1(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__and2b_1 _08812_ (.A_N(net113),
    .B(net81),
    .X(_03578_));
 sky130_fd_sc_hd__a21oi_1 _08813_ (.A1(_03472_),
    .A2(_03577_),
    .B1(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__or2_1 _08814_ (.A(_03469_),
    .B(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__o221a_1 _08815_ (.A1(net114),
    .A2(_03460_),
    .B1(_03474_),
    .B2(_03572_),
    .C1(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__or2_1 _08816_ (.A(_03459_),
    .B(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__inv_2 _08817_ (.A(net86),
    .Y(_03583_));
 sky130_fd_sc_hd__inv_2 _08818_ (.A(net84),
    .Y(_03584_));
 sky130_fd_sc_hd__and2b_1 _08819_ (.A_N(net115),
    .B(net83),
    .X(_03585_));
 sky130_fd_sc_hd__o21ai_1 _08820_ (.A1(_03454_),
    .A2(_03455_),
    .B1(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__o21a_1 _08821_ (.A1(net116),
    .A2(_03584_),
    .B1(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__and2b_1 _08822_ (.A_N(net117),
    .B(net85),
    .X(_03588_));
 sky130_fd_sc_hd__nand2_1 _08823_ (.A(_03449_),
    .B(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__o221a_1 _08824_ (.A1(net118),
    .A2(_03583_),
    .B1(_03453_),
    .B2(_03587_),
    .C1(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__o31a_1 _08825_ (.A1(_03453_),
    .A2(_03456_),
    .A3(_03582_),
    .B1(_03590_),
    .X(_03591_));
 sky130_fd_sc_hd__inv_2 _08826_ (.A(net119),
    .Y(_03592_));
 sky130_fd_sc_hd__and2b_1 _08827_ (.A_N(net120),
    .B(net88),
    .X(_03593_));
 sky130_fd_sc_hd__a31o_1 _08828_ (.A1(_03592_),
    .A2(net87),
    .A3(_03445_),
    .B1(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__and2b_1 _08829_ (.A_N(net122),
    .B(net90),
    .X(_03595_));
 sky130_fd_sc_hd__and2b_1 _08830_ (.A_N(net123),
    .B(net91),
    .X(_03596_));
 sky130_fd_sc_hd__a21o_1 _08831_ (.A1(_03434_),
    .A2(_03595_),
    .B1(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__a31o_1 _08832_ (.A1(_03434_),
    .A2(_03438_),
    .A3(_03594_),
    .B1(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__o21ba_2 _08833_ (.A1(_03446_),
    .A2(_03591_),
    .B1_N(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__a21o_1 _08834_ (.A1(_03434_),
    .A2(_03599_),
    .B1(_03596_),
    .X(_03600_));
 sky130_fd_sc_hd__and3_1 _08835_ (.A(is_slti_blt_slt),
    .B(_03431_),
    .C(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__inv_2 _08836_ (.A(instr_bge),
    .Y(_03602_));
 sky130_fd_sc_hd__nor2_1 _08837_ (.A(_03602_),
    .B(_03600_),
    .Y(_03603_));
 sky130_fd_sc_hd__or4_2 _08838_ (.A(_03446_),
    .B(_03453_),
    .C(_03456_),
    .D(_03459_),
    .X(_03604_));
 sky130_fd_sc_hd__nor2_1 _08839_ (.A(_03474_),
    .B(_03489_),
    .Y(_03605_));
 sky130_fd_sc_hd__nor2_1 _08840_ (.A(_03530_),
    .B(net92),
    .Y(_03606_));
 sky130_fd_sc_hd__and2_1 _08841_ (.A(net124),
    .B(net92),
    .X(_03607_));
 sky130_fd_sc_hd__nor2_1 _08842_ (.A(_03606_),
    .B(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__clkbuf_4 _08843_ (.A(net99),
    .X(_03609_));
 sky130_fd_sc_hd__nor2_1 _08844_ (.A(net67),
    .B(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__and2_1 _08845_ (.A(net67),
    .B(_03609_),
    .X(_03611_));
 sky130_fd_sc_hd__nor2_1 _08846_ (.A(_03610_),
    .B(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__nor2_1 _08847_ (.A(net128),
    .B(net96),
    .Y(_03613_));
 sky130_fd_sc_hd__and2_1 _08848_ (.A(net128),
    .B(_03518_),
    .X(_03614_));
 sky130_fd_sc_hd__nor2_1 _08849_ (.A(_03613_),
    .B(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__or4_1 _08850_ (.A(_03608_),
    .B(_03521_),
    .C(_03612_),
    .D(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__or2_1 _08851_ (.A(net105),
    .B(net73),
    .X(_03617_));
 sky130_fd_sc_hd__nand2_1 _08852_ (.A(net105),
    .B(net73),
    .Y(_03618_));
 sky130_fd_sc_hd__nand2_1 _08853_ (.A(_03617_),
    .B(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__and3_1 _08854_ (.A(_03534_),
    .B(_03493_),
    .C(_03619_),
    .X(_03620_));
 sky130_fd_sc_hd__and4b_1 _08855_ (.A_N(_03535_),
    .B(_03496_),
    .C(_03499_),
    .D(_03529_),
    .X(_03621_));
 sky130_fd_sc_hd__and4bb_1 _08856_ (.A_N(_03616_),
    .B_N(_03526_),
    .C(_03620_),
    .D(_03621_),
    .X(_03622_));
 sky130_fd_sc_hd__and4b_1 _08857_ (.A_N(_03604_),
    .B(_03516_),
    .C(_03605_),
    .D(_03622_),
    .X(_03623_));
 sky130_fd_sc_hd__inv_2 _08858_ (.A(_03623_),
    .Y(_03624_));
 sky130_fd_sc_hd__and2_1 _08859_ (.A(is_sltiu_bltu_sltu),
    .B(_03431_),
    .X(_03625_));
 sky130_fd_sc_hd__a211o_1 _08860_ (.A1(is_slti_blt_slt),
    .A2(_03431_),
    .B1(_03625_),
    .C1(_03430_),
    .X(_03626_));
 sky130_fd_sc_hd__inv_2 _08861_ (.A(_03626_),
    .Y(_03627_));
 sky130_fd_sc_hd__mux2_1 _08862_ (.A0(instr_bgeu),
    .A1(_03625_),
    .S(_03599_),
    .X(_03628_));
 sky130_fd_sc_hd__a211o_1 _08863_ (.A1(instr_bne),
    .A2(_03624_),
    .B1(_03627_),
    .C1(_03628_),
    .X(_03629_));
 sky130_fd_sc_hd__o32a_2 _08864_ (.A1(_03601_),
    .A2(_03603_),
    .A3(_03629_),
    .B1(_03626_),
    .B2(_03623_),
    .X(_03630_));
 sky130_fd_sc_hd__clkbuf_4 _08865_ (.A(_03311_),
    .X(_03631_));
 sky130_fd_sc_hd__and4_1 _08866_ (.A(_03309_),
    .B(_03384_),
    .C(_03305_),
    .D(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__and2_2 _08867_ (.A(_03199_),
    .B(_03310_),
    .X(_03633_));
 sky130_fd_sc_hd__clkbuf_2 _08868_ (.A(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__clkbuf_4 _08869_ (.A(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__buf_4 _08870_ (.A(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__o2bb2a_1 _08871_ (.A1_N(_03630_),
    .A2_N(_03632_),
    .B1(_01226_),
    .B2(_03636_),
    .X(_00000_));
 sky130_fd_sc_hd__buf_2 _08872_ (.A(_03312_),
    .X(_03637_));
 sky130_fd_sc_hd__clkbuf_4 _08873_ (.A(_03637_),
    .X(_03638_));
 sky130_fd_sc_hd__buf_8 _08874_ (.A(_00068_),
    .X(_03639_));
 sky130_fd_sc_hd__buf_8 _08875_ (.A(_00064_),
    .X(_03640_));
 sky130_fd_sc_hd__buf_8 _08876_ (.A(_03640_),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_8 _08877_ (.A(_00065_),
    .X(_03642_));
 sky130_fd_sc_hd__clkbuf_8 _08878_ (.A(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__mux4_1 _08879_ (.A0(\cpuregs.regs[4][2] ),
    .A1(\cpuregs.regs[5][2] ),
    .A2(\cpuregs.regs[6][2] ),
    .A3(\cpuregs.regs[7][2] ),
    .S0(_03641_),
    .S1(_03643_),
    .X(_03644_));
 sky130_fd_sc_hd__buf_8 _08880_ (.A(_03640_),
    .X(_03645_));
 sky130_fd_sc_hd__buf_4 _08881_ (.A(_00065_),
    .X(_03646_));
 sky130_fd_sc_hd__buf_8 _08882_ (.A(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__mux4_1 _08883_ (.A0(\cpuregs.regs[0][2] ),
    .A1(\cpuregs.regs[1][2] ),
    .A2(\cpuregs.regs[2][2] ),
    .A3(\cpuregs.regs[3][2] ),
    .S0(_03645_),
    .S1(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__clkbuf_8 _08884_ (.A(_03640_),
    .X(_03649_));
 sky130_fd_sc_hd__mux4_1 _08885_ (.A0(\cpuregs.regs[12][2] ),
    .A1(\cpuregs.regs[13][2] ),
    .A2(\cpuregs.regs[14][2] ),
    .A3(\cpuregs.regs[15][2] ),
    .S0(_03649_),
    .S1(_03643_),
    .X(_03650_));
 sky130_fd_sc_hd__mux4_1 _08886_ (.A0(\cpuregs.regs[8][2] ),
    .A1(\cpuregs.regs[9][2] ),
    .A2(\cpuregs.regs[10][2] ),
    .A3(\cpuregs.regs[11][2] ),
    .S0(_03649_),
    .S1(_03643_),
    .X(_03651_));
 sky130_fd_sc_hd__inv_2 _08887_ (.A(_00066_),
    .Y(_03652_));
 sky130_fd_sc_hd__clkbuf_8 _08888_ (.A(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__clkbuf_8 _08889_ (.A(_00067_),
    .X(_03654_));
 sky130_fd_sc_hd__mux4_1 _08890_ (.A0(_03644_),
    .A1(_03648_),
    .A2(_03650_),
    .A3(_03651_),
    .S0(_03653_),
    .S1(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__inv_2 _08891_ (.A(_00067_),
    .Y(_03656_));
 sky130_fd_sc_hd__buf_4 _08892_ (.A(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__clkbuf_8 _08893_ (.A(_00064_),
    .X(_03658_));
 sky130_fd_sc_hd__buf_4 _08894_ (.A(_00065_),
    .X(_03659_));
 sky130_fd_sc_hd__mux4_1 _08895_ (.A0(\cpuregs.regs[20][2] ),
    .A1(\cpuregs.regs[21][2] ),
    .A2(\cpuregs.regs[22][2] ),
    .A3(\cpuregs.regs[23][2] ),
    .S0(_03658_),
    .S1(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__buf_6 _08896_ (.A(_00064_),
    .X(_03661_));
 sky130_fd_sc_hd__clkbuf_8 _08897_ (.A(_00065_),
    .X(_03662_));
 sky130_fd_sc_hd__mux4_1 _08898_ (.A0(\cpuregs.regs[16][2] ),
    .A1(\cpuregs.regs[17][2] ),
    .A2(\cpuregs.regs[18][2] ),
    .A3(\cpuregs.regs[19][2] ),
    .S0(_03661_),
    .S1(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__buf_6 _08899_ (.A(_03652_),
    .X(_03664_));
 sky130_fd_sc_hd__mux2_1 _08900_ (.A0(_03660_),
    .A1(_03663_),
    .S(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__buf_4 _08901_ (.A(_00066_),
    .X(_03666_));
 sky130_fd_sc_hd__mux4_1 _08902_ (.A0(\cpuregs.regs[24][2] ),
    .A1(\cpuregs.regs[25][2] ),
    .A2(\cpuregs.regs[26][2] ),
    .A3(\cpuregs.regs[27][2] ),
    .S0(_03658_),
    .S1(_03659_),
    .X(_03667_));
 sky130_fd_sc_hd__or2_1 _08903_ (.A(_03666_),
    .B(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__clkbuf_8 _08904_ (.A(_00064_),
    .X(_03669_));
 sky130_fd_sc_hd__buf_6 _08905_ (.A(_03669_),
    .X(_03670_));
 sky130_fd_sc_hd__buf_4 _08906_ (.A(_03646_),
    .X(_03671_));
 sky130_fd_sc_hd__mux4_1 _08907_ (.A0(\cpuregs.regs[28][2] ),
    .A1(\cpuregs.regs[29][2] ),
    .A2(\cpuregs.regs[30][2] ),
    .A3(\cpuregs.regs[31][2] ),
    .S0(_03670_),
    .S1(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__o21a_1 _08908_ (.A1(_03664_),
    .A2(_03672_),
    .B1(_00067_),
    .X(_03673_));
 sky130_fd_sc_hd__clkinv_4 _08909_ (.A(_00068_),
    .Y(_03674_));
 sky130_fd_sc_hd__buf_4 _08910_ (.A(_03674_),
    .X(_03675_));
 sky130_fd_sc_hd__a221o_1 _08911_ (.A1(_03657_),
    .A2(_03665_),
    .B1(_03668_),
    .B2(_03673_),
    .C1(_03675_),
    .X(_03676_));
 sky130_fd_sc_hd__o21a_1 _08912_ (.A1(_03639_),
    .A2(_03655_),
    .B1(_03676_),
    .X(_03677_));
 sky130_fd_sc_hd__or3_1 _08913_ (.A(\cpuregs.raddr2[1] ),
    .B(\cpuregs.raddr2[0] ),
    .C(\cpuregs.raddr2[2] ),
    .X(_03678_));
 sky130_fd_sc_hd__or3_4 _08914_ (.A(\cpuregs.raddr2[3] ),
    .B(\cpuregs.raddr2[4] ),
    .C(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__clkbuf_4 _08915_ (.A(_03312_),
    .X(_03680_));
 sky130_fd_sc_hd__a21oi_1 _08916_ (.A1(_03677_),
    .A2(_03679_),
    .B1(_03680_),
    .Y(_03681_));
 sky130_fd_sc_hd__a31o_1 _08917_ (.A1(_03638_),
    .A2(_03313_),
    .A3(_03315_),
    .B1(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__a21oi_1 _08918_ (.A1(\reg_sh[2] ),
    .A2(_03638_),
    .B1(_03682_),
    .Y(_00061_));
 sky130_fd_sc_hd__buf_6 _08919_ (.A(_03654_),
    .X(_03683_));
 sky130_fd_sc_hd__buf_6 _08920_ (.A(_03662_),
    .X(_03684_));
 sky130_fd_sc_hd__mux4_1 _08921_ (.A0(\cpuregs.regs[8][3] ),
    .A1(\cpuregs.regs[9][3] ),
    .A2(\cpuregs.regs[10][3] ),
    .A3(\cpuregs.regs[11][3] ),
    .S0(_03641_),
    .S1(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__mux4_1 _08922_ (.A0(\cpuregs.regs[12][3] ),
    .A1(\cpuregs.regs[13][3] ),
    .A2(\cpuregs.regs[14][3] ),
    .A3(\cpuregs.regs[15][3] ),
    .S0(_03641_),
    .S1(_03684_),
    .X(_03686_));
 sky130_fd_sc_hd__buf_6 _08923_ (.A(_03666_),
    .X(_03687_));
 sky130_fd_sc_hd__mux2_1 _08924_ (.A0(_03685_),
    .A1(_03686_),
    .S(_03687_),
    .X(_03688_));
 sky130_fd_sc_hd__mux4_1 _08925_ (.A0(\cpuregs.regs[4][3] ),
    .A1(\cpuregs.regs[5][3] ),
    .A2(\cpuregs.regs[6][3] ),
    .A3(\cpuregs.regs[7][3] ),
    .S0(_03658_),
    .S1(_03659_),
    .X(_03689_));
 sky130_fd_sc_hd__mux4_1 _08926_ (.A0(\cpuregs.regs[0][3] ),
    .A1(\cpuregs.regs[1][3] ),
    .A2(\cpuregs.regs[2][3] ),
    .A3(\cpuregs.regs[3][3] ),
    .S0(_03658_),
    .S1(_03659_),
    .X(_03690_));
 sky130_fd_sc_hd__mux2_1 _08927_ (.A0(_03689_),
    .A1(_03690_),
    .S(_03664_),
    .X(_03691_));
 sky130_fd_sc_hd__clkbuf_8 _08928_ (.A(_00068_),
    .X(_03692_));
 sky130_fd_sc_hd__a21o_1 _08929_ (.A1(_03657_),
    .A2(_03691_),
    .B1(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__a21o_1 _08930_ (.A1(_03683_),
    .A2(_03688_),
    .B1(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__mux4_1 _08931_ (.A0(\cpuregs.regs[24][3] ),
    .A1(\cpuregs.regs[25][3] ),
    .A2(\cpuregs.regs[26][3] ),
    .A3(\cpuregs.regs[27][3] ),
    .S0(_03641_),
    .S1(_03684_),
    .X(_03695_));
 sky130_fd_sc_hd__mux4_1 _08932_ (.A0(\cpuregs.regs[28][3] ),
    .A1(\cpuregs.regs[29][3] ),
    .A2(\cpuregs.regs[30][3] ),
    .A3(\cpuregs.regs[31][3] ),
    .S0(_03641_),
    .S1(_03684_),
    .X(_03696_));
 sky130_fd_sc_hd__mux2_1 _08933_ (.A0(_03695_),
    .A1(_03696_),
    .S(_03687_),
    .X(_03697_));
 sky130_fd_sc_hd__mux4_1 _08934_ (.A0(\cpuregs.regs[20][3] ),
    .A1(\cpuregs.regs[21][3] ),
    .A2(\cpuregs.regs[22][3] ),
    .A3(\cpuregs.regs[23][3] ),
    .S0(_03658_),
    .S1(_03659_),
    .X(_03698_));
 sky130_fd_sc_hd__mux4_1 _08935_ (.A0(\cpuregs.regs[16][3] ),
    .A1(\cpuregs.regs[17][3] ),
    .A2(\cpuregs.regs[18][3] ),
    .A3(\cpuregs.regs[19][3] ),
    .S0(_03658_),
    .S1(_03659_),
    .X(_03699_));
 sky130_fd_sc_hd__mux2_1 _08936_ (.A0(_03698_),
    .A1(_03699_),
    .S(_03664_),
    .X(_03700_));
 sky130_fd_sc_hd__a21o_1 _08937_ (.A1(_03657_),
    .A2(_03700_),
    .B1(_03675_),
    .X(_03701_));
 sky130_fd_sc_hd__a21o_1 _08938_ (.A1(_03683_),
    .A2(_03697_),
    .B1(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__and3_2 _08939_ (.A(_03679_),
    .B(_03694_),
    .C(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__or3b_1 _08940_ (.A(\reg_sh[3] ),
    .B(\reg_sh[2] ),
    .C_N(\reg_sh[4] ),
    .X(_03704_));
 sky130_fd_sc_hd__a21bo_1 _08941_ (.A1(\reg_sh[3] ),
    .A2(\reg_sh[2] ),
    .B1_N(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__o22a_1 _08942_ (.A1(_03638_),
    .A2(_03703_),
    .B1(_03705_),
    .B2(_03400_),
    .X(_00062_));
 sky130_fd_sc_hd__o21a_1 _08943_ (.A1(\reg_sh[3] ),
    .A2(\reg_sh[2] ),
    .B1(\reg_sh[4] ),
    .X(_03706_));
 sky130_fd_sc_hd__mux4_1 _08944_ (.A0(\cpuregs.regs[8][4] ),
    .A1(\cpuregs.regs[9][4] ),
    .A2(\cpuregs.regs[10][4] ),
    .A3(\cpuregs.regs[11][4] ),
    .S0(_03649_),
    .S1(_03643_),
    .X(_03707_));
 sky130_fd_sc_hd__mux4_1 _08945_ (.A0(\cpuregs.regs[12][4] ),
    .A1(\cpuregs.regs[13][4] ),
    .A2(\cpuregs.regs[14][4] ),
    .A3(\cpuregs.regs[15][4] ),
    .S0(_03649_),
    .S1(_03643_),
    .X(_03708_));
 sky130_fd_sc_hd__clkbuf_8 _08946_ (.A(_03666_),
    .X(_03709_));
 sky130_fd_sc_hd__mux2_1 _08947_ (.A0(_03707_),
    .A1(_03708_),
    .S(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__mux4_1 _08948_ (.A0(\cpuregs.regs[4][4] ),
    .A1(\cpuregs.regs[5][4] ),
    .A2(\cpuregs.regs[6][4] ),
    .A3(\cpuregs.regs[7][4] ),
    .S0(_03661_),
    .S1(_03662_),
    .X(_03711_));
 sky130_fd_sc_hd__mux4_1 _08949_ (.A0(\cpuregs.regs[0][4] ),
    .A1(\cpuregs.regs[1][4] ),
    .A2(\cpuregs.regs[2][4] ),
    .A3(\cpuregs.regs[3][4] ),
    .S0(_03661_),
    .S1(_03662_),
    .X(_03712_));
 sky130_fd_sc_hd__clkbuf_8 _08950_ (.A(_03652_),
    .X(_03713_));
 sky130_fd_sc_hd__mux2_1 _08951_ (.A0(_03711_),
    .A1(_03712_),
    .S(_03713_),
    .X(_03714_));
 sky130_fd_sc_hd__a21o_1 _08952_ (.A1(_03657_),
    .A2(_03714_),
    .B1(_03692_),
    .X(_03715_));
 sky130_fd_sc_hd__a21o_1 _08953_ (.A1(_03683_),
    .A2(_03710_),
    .B1(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__mux4_1 _08954_ (.A0(\cpuregs.regs[28][4] ),
    .A1(\cpuregs.regs[29][4] ),
    .A2(\cpuregs.regs[30][4] ),
    .A3(\cpuregs.regs[31][4] ),
    .S0(_03649_),
    .S1(_03643_),
    .X(_03717_));
 sky130_fd_sc_hd__mux4_1 _08955_ (.A0(\cpuregs.regs[24][4] ),
    .A1(\cpuregs.regs[25][4] ),
    .A2(\cpuregs.regs[26][4] ),
    .A3(\cpuregs.regs[27][4] ),
    .S0(_03649_),
    .S1(_03643_),
    .X(_03718_));
 sky130_fd_sc_hd__clkbuf_8 _08956_ (.A(_03713_),
    .X(_03719_));
 sky130_fd_sc_hd__mux2_1 _08957_ (.A0(_03717_),
    .A1(_03718_),
    .S(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__mux4_1 _08958_ (.A0(\cpuregs.regs[20][4] ),
    .A1(\cpuregs.regs[21][4] ),
    .A2(\cpuregs.regs[22][4] ),
    .A3(\cpuregs.regs[23][4] ),
    .S0(_03661_),
    .S1(_03662_),
    .X(_03721_));
 sky130_fd_sc_hd__mux4_1 _08959_ (.A0(\cpuregs.regs[16][4] ),
    .A1(\cpuregs.regs[17][4] ),
    .A2(\cpuregs.regs[18][4] ),
    .A3(\cpuregs.regs[19][4] ),
    .S0(_03661_),
    .S1(_03662_),
    .X(_03722_));
 sky130_fd_sc_hd__mux2_1 _08960_ (.A0(_03721_),
    .A1(_03722_),
    .S(_03713_),
    .X(_03723_));
 sky130_fd_sc_hd__a21o_1 _08961_ (.A1(_03656_),
    .A2(_03723_),
    .B1(_03675_),
    .X(_03724_));
 sky130_fd_sc_hd__a21o_1 _08962_ (.A1(_03683_),
    .A2(_03720_),
    .B1(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__and3_2 _08963_ (.A(_03679_),
    .B(_03716_),
    .C(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__o22a_1 _08964_ (.A1(_03400_),
    .A2(_03706_),
    .B1(_03726_),
    .B2(_03638_),
    .X(_00063_));
 sky130_fd_sc_hd__buf_4 _08965_ (.A(_03205_),
    .X(_03727_));
 sky130_fd_sc_hd__buf_4 _08966_ (.A(_03727_),
    .X(_03728_));
 sky130_fd_sc_hd__clkbuf_4 _08967_ (.A(_03200_),
    .X(_03729_));
 sky130_fd_sc_hd__clkbuf_4 _08968_ (.A(_03729_),
    .X(_03730_));
 sky130_fd_sc_hd__mux2_1 _08969_ (.A0(net36),
    .A1(\mem_rdata_q[12] ),
    .S(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__nand2_1 _08970_ (.A(_03231_),
    .B(_03731_),
    .Y(_03732_));
 sky130_fd_sc_hd__mux2_1 _08971_ (.A0(net53),
    .A1(\mem_rdata_q[28] ),
    .S(_03730_),
    .X(_03733_));
 sky130_fd_sc_hd__nand2_1 _08972_ (.A(_03203_),
    .B(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__nor2_1 _08973_ (.A(\mem_16bit_buffer[12] ),
    .B(_03728_),
    .Y(_03735_));
 sky130_fd_sc_hd__a31oi_4 _08974_ (.A1(_03728_),
    .A2(_03732_),
    .A3(_03734_),
    .B1(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__clkbuf_4 _08975_ (.A(_03736_),
    .X(_03737_));
 sky130_fd_sc_hd__or2_2 _08976_ (.A(_03229_),
    .B(_03237_),
    .X(_03738_));
 sky130_fd_sc_hd__nor2b_4 _08977_ (.A(_03213_),
    .B_N(_03206_),
    .Y(_03739_));
 sky130_fd_sc_hd__mux2_1 _08978_ (.A0(\mem_rdata_q[14] ),
    .A1(net38),
    .S(_03208_),
    .X(_03740_));
 sky130_fd_sc_hd__mux2_1 _08979_ (.A0(\mem_rdata_q[30] ),
    .A1(net56),
    .S(_03208_),
    .X(_03741_));
 sky130_fd_sc_hd__mux2_1 _08980_ (.A0(_03740_),
    .A1(_03741_),
    .S(_03203_),
    .X(_03742_));
 sky130_fd_sc_hd__mux2_4 _08981_ (.A0(\mem_16bit_buffer[14] ),
    .A1(_03742_),
    .S(_03205_),
    .X(_03743_));
 sky130_fd_sc_hd__mux2_1 _08982_ (.A0(\mem_rdata_q[29] ),
    .A1(net54),
    .S(_03208_),
    .X(_03744_));
 sky130_fd_sc_hd__mux2_1 _08983_ (.A0(\mem_rdata_q[13] ),
    .A1(net37),
    .S(_03208_),
    .X(_03745_));
 sky130_fd_sc_hd__mux2_1 _08984_ (.A0(_03744_),
    .A1(_03745_),
    .S(_03230_),
    .X(_03746_));
 sky130_fd_sc_hd__mux2_4 _08985_ (.A0(\mem_16bit_buffer[13] ),
    .A1(_03746_),
    .S(_03727_),
    .X(_03747_));
 sky130_fd_sc_hd__inv_2 _08986_ (.A(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__or2_2 _08987_ (.A(_03743_),
    .B(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__nand2_1 _08988_ (.A(_03739_),
    .B(_03749_),
    .Y(_03750_));
 sky130_fd_sc_hd__nor2_1 _08989_ (.A(_03738_),
    .B(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__mux2_1 _08990_ (.A0(\mem_rdata_q[31] ),
    .A1(net57),
    .S(_03227_),
    .X(_03752_));
 sky130_fd_sc_hd__clkbuf_4 _08991_ (.A(mem_la_secondword),
    .X(_03753_));
 sky130_fd_sc_hd__nor2_2 _08992_ (.A(_03753_),
    .B(_03203_),
    .Y(_03754_));
 sky130_fd_sc_hd__mux2_1 _08993_ (.A0(net39),
    .A1(\mem_rdata_q[15] ),
    .S(_03729_),
    .X(_03755_));
 sky130_fd_sc_hd__a22o_1 _08994_ (.A1(_03752_),
    .A2(_03754_),
    .B1(_03755_),
    .B2(_03753_),
    .X(_03756_));
 sky130_fd_sc_hd__clkbuf_4 _08995_ (.A(_03227_),
    .X(_03757_));
 sky130_fd_sc_hd__mux2_1 _08996_ (.A0(\mem_rdata_q[31] ),
    .A1(_03756_),
    .S(_03757_),
    .X(_03758_));
 sky130_fd_sc_hd__mux2_1 _08997_ (.A0(\mem_rdata_q[27] ),
    .A1(net52),
    .S(_03208_),
    .X(_03759_));
 sky130_fd_sc_hd__mux2_1 _08998_ (.A0(\mem_rdata_q[11] ),
    .A1(net35),
    .S(_03208_),
    .X(_03760_));
 sky130_fd_sc_hd__mux2_1 _08999_ (.A0(_03759_),
    .A1(_03760_),
    .S(_03230_),
    .X(_03761_));
 sky130_fd_sc_hd__mux2_4 _09000_ (.A0(\mem_16bit_buffer[11] ),
    .A1(_03761_),
    .S(_03727_),
    .X(_03762_));
 sky130_fd_sc_hd__clkbuf_4 _09001_ (.A(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__nand2_1 _09002_ (.A(_03231_),
    .B(_03755_),
    .Y(_03764_));
 sky130_fd_sc_hd__nand2_1 _09003_ (.A(_03203_),
    .B(_03752_),
    .Y(_03765_));
 sky130_fd_sc_hd__nor2_1 _09004_ (.A(\mem_16bit_buffer[15] ),
    .B(_03727_),
    .Y(_03766_));
 sky130_fd_sc_hd__a31o_4 _09005_ (.A1(_03727_),
    .A2(_03764_),
    .A3(_03765_),
    .B1(_03766_),
    .X(_03767_));
 sky130_fd_sc_hd__or2_2 _09006_ (.A(_03743_),
    .B(_03747_),
    .X(_03768_));
 sky130_fd_sc_hd__or2_1 _09007_ (.A(_03767_),
    .B(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__clkbuf_4 _09008_ (.A(_03769_),
    .X(_03770_));
 sky130_fd_sc_hd__mux2_1 _09009_ (.A0(net51),
    .A1(\mem_rdata_q[26] ),
    .S(_03729_),
    .X(_03771_));
 sky130_fd_sc_hd__mux2_1 _09010_ (.A0(net34),
    .A1(\mem_rdata_q[10] ),
    .S(_03729_),
    .X(_03772_));
 sky130_fd_sc_hd__mux2_1 _09011_ (.A0(_03771_),
    .A1(_03772_),
    .S(_03231_),
    .X(_03773_));
 sky130_fd_sc_hd__mux2_1 _09012_ (.A0(\mem_16bit_buffer[10] ),
    .A1(_03773_),
    .S(_03727_),
    .X(_03774_));
 sky130_fd_sc_hd__inv_2 _09013_ (.A(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__nand2_2 _09014_ (.A(_03762_),
    .B(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hd__inv_2 _09015_ (.A(_03776_),
    .Y(_03777_));
 sky130_fd_sc_hd__a211o_1 _09016_ (.A1(_03758_),
    .A2(_03763_),
    .B1(_03770_),
    .C1(_03777_),
    .X(_03778_));
 sky130_fd_sc_hd__nand2_2 _09017_ (.A(_03743_),
    .B(_03748_),
    .Y(_03779_));
 sky130_fd_sc_hd__a31oi_2 _09018_ (.A1(_03728_),
    .A2(_03764_),
    .A3(_03765_),
    .B1(_03766_),
    .Y(_03780_));
 sky130_fd_sc_hd__clkbuf_4 _09019_ (.A(_03780_),
    .X(_03781_));
 sky130_fd_sc_hd__nor2_1 _09020_ (.A(_03747_),
    .B(_03781_),
    .Y(_03782_));
 sky130_fd_sc_hd__clkbuf_4 _09021_ (.A(_03206_),
    .X(_03783_));
 sky130_fd_sc_hd__or2_1 _09022_ (.A(_03783_),
    .B(_03213_),
    .X(_03784_));
 sky130_fd_sc_hd__nor2_1 _09023_ (.A(_03782_),
    .B(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__and2_1 _09024_ (.A(_03779_),
    .B(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__or2b_1 _09025_ (.A(_03213_),
    .B_N(_03206_),
    .X(_03787_));
 sky130_fd_sc_hd__nor2_1 _09026_ (.A(_03787_),
    .B(_03749_),
    .Y(_03788_));
 sky130_fd_sc_hd__nand2b_2 _09027_ (.A_N(_03206_),
    .B(_03213_),
    .Y(_03789_));
 sky130_fd_sc_hd__nor2b_2 _09028_ (.A(_03206_),
    .B_N(_03213_),
    .Y(_03790_));
 sky130_fd_sc_hd__mux2_1 _09029_ (.A0(net46),
    .A1(\mem_rdata_q[21] ),
    .S(_03729_),
    .X(_03791_));
 sky130_fd_sc_hd__mux2_1 _09030_ (.A0(net60),
    .A1(\mem_rdata_q[5] ),
    .S(_03729_),
    .X(_03792_));
 sky130_fd_sc_hd__mux2_1 _09031_ (.A0(_03791_),
    .A1(_03792_),
    .S(_03231_),
    .X(_03793_));
 sky130_fd_sc_hd__mux2_1 _09032_ (.A0(\mem_16bit_buffer[5] ),
    .A1(_03793_),
    .S(_03727_),
    .X(_03794_));
 sky130_fd_sc_hd__mux2_1 _09033_ (.A0(\mem_rdata_q[22] ),
    .A1(net47),
    .S(_03227_),
    .X(_03795_));
 sky130_fd_sc_hd__mux2_1 _09034_ (.A0(\mem_rdata_q[6] ),
    .A1(net61),
    .S(_03227_),
    .X(_03796_));
 sky130_fd_sc_hd__mux2_1 _09035_ (.A0(_03795_),
    .A1(_03796_),
    .S(_03231_),
    .X(_03797_));
 sky130_fd_sc_hd__mux2_2 _09036_ (.A0(\mem_16bit_buffer[6] ),
    .A1(_03797_),
    .S(_03727_),
    .X(_03798_));
 sky130_fd_sc_hd__nor2_2 _09037_ (.A(_03794_),
    .B(_03798_),
    .Y(_03799_));
 sky130_fd_sc_hd__inv_2 _09038_ (.A(_03799_),
    .Y(_03800_));
 sky130_fd_sc_hd__mux2_1 _09039_ (.A0(net59),
    .A1(\mem_rdata_q[4] ),
    .S(_03730_),
    .X(_03801_));
 sky130_fd_sc_hd__mux2_1 _09040_ (.A0(net45),
    .A1(\mem_rdata_q[20] ),
    .S(_03730_),
    .X(_03802_));
 sky130_fd_sc_hd__mux2_1 _09041_ (.A0(_03801_),
    .A1(_03802_),
    .S(_03203_),
    .X(_03803_));
 sky130_fd_sc_hd__mux2_2 _09042_ (.A0(\mem_16bit_buffer[4] ),
    .A1(_03803_),
    .S(_03728_),
    .X(_03804_));
 sky130_fd_sc_hd__mux2_1 _09043_ (.A0(net43),
    .A1(\mem_rdata_q[19] ),
    .S(_03730_),
    .X(_03805_));
 sky130_fd_sc_hd__nand2_1 _09044_ (.A(_03203_),
    .B(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__mux2_1 _09045_ (.A0(net58),
    .A1(\mem_rdata_q[3] ),
    .S(_03730_),
    .X(_03807_));
 sky130_fd_sc_hd__nand2_1 _09046_ (.A(_03231_),
    .B(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__nor2_1 _09047_ (.A(\mem_16bit_buffer[3] ),
    .B(_03728_),
    .Y(_03809_));
 sky130_fd_sc_hd__a31oi_4 _09048_ (.A1(_03728_),
    .A2(_03806_),
    .A3(_03808_),
    .B1(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hd__mux2_1 _09049_ (.A0(net42),
    .A1(\mem_rdata_q[18] ),
    .S(_03729_),
    .X(_03811_));
 sky130_fd_sc_hd__mux2_1 _09050_ (.A0(net55),
    .A1(\mem_rdata_q[2] ),
    .S(_03729_),
    .X(_03812_));
 sky130_fd_sc_hd__mux2_1 _09051_ (.A0(_03811_),
    .A1(_03812_),
    .S(_03231_),
    .X(_03813_));
 sky130_fd_sc_hd__mux2_1 _09052_ (.A0(\mem_16bit_buffer[2] ),
    .A1(_03813_),
    .S(_03728_),
    .X(_03814_));
 sky130_fd_sc_hd__or2_1 _09053_ (.A(_03810_),
    .B(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__nor3_4 _09054_ (.A(_03800_),
    .B(_03804_),
    .C(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hd__nand2_1 _09055_ (.A(_03790_),
    .B(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__a31o_1 _09056_ (.A1(_03728_),
    .A2(_03732_),
    .A3(_03734_),
    .B1(_03735_),
    .X(_03818_));
 sky130_fd_sc_hd__mux2_1 _09057_ (.A0(\mem_rdata_q[23] ),
    .A1(net48),
    .S(_03208_),
    .X(_03819_));
 sky130_fd_sc_hd__mux2_1 _09058_ (.A0(net62),
    .A1(\mem_rdata_q[7] ),
    .S(_03200_),
    .X(_03820_));
 sky130_fd_sc_hd__mux2_1 _09059_ (.A0(_03819_),
    .A1(_03820_),
    .S(_03231_),
    .X(_03821_));
 sky130_fd_sc_hd__mux2_2 _09060_ (.A0(\mem_16bit_buffer[7] ),
    .A1(_03821_),
    .S(_03727_),
    .X(_03822_));
 sky130_fd_sc_hd__mux2_1 _09061_ (.A0(net64),
    .A1(\mem_rdata_q[9] ),
    .S(_03729_),
    .X(_03823_));
 sky130_fd_sc_hd__mux2_1 _09062_ (.A0(net50),
    .A1(\mem_rdata_q[25] ),
    .S(_03729_),
    .X(_03824_));
 sky130_fd_sc_hd__mux2_1 _09063_ (.A0(_03823_),
    .A1(_03824_),
    .S(_03203_),
    .X(_03825_));
 sky130_fd_sc_hd__mux2_4 _09064_ (.A0(\mem_16bit_buffer[9] ),
    .A1(_03825_),
    .S(_03727_),
    .X(_03826_));
 sky130_fd_sc_hd__or4_1 _09065_ (.A(_03762_),
    .B(_03774_),
    .C(_03822_),
    .D(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__mux2_1 _09066_ (.A0(\mem_rdata_q[24] ),
    .A1(net49),
    .S(_03227_),
    .X(_03828_));
 sky130_fd_sc_hd__or2_1 _09067_ (.A(\mem_rdata_q[8] ),
    .B(_03208_),
    .X(_03829_));
 sky130_fd_sc_hd__o21a_1 _09068_ (.A1(net63),
    .A2(_03730_),
    .B1(_03829_),
    .X(_03830_));
 sky130_fd_sc_hd__mux2_1 _09069_ (.A0(_03828_),
    .A1(_03830_),
    .S(_03231_),
    .X(_03831_));
 sky130_fd_sc_hd__mux2_1 _09070_ (.A0(\mem_16bit_buffer[8] ),
    .A1(_03831_),
    .S(_03728_),
    .X(_03832_));
 sky130_fd_sc_hd__nor2_2 _09071_ (.A(_03827_),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__or3b_1 _09072_ (.A(_03818_),
    .B(_03770_),
    .C_N(_03833_),
    .X(_03834_));
 sky130_fd_sc_hd__nor2_2 _09073_ (.A(_03215_),
    .B(_03738_),
    .Y(_03835_));
 sky130_fd_sc_hd__o221a_1 _09074_ (.A1(_03748_),
    .A2(_03789_),
    .B1(_03817_),
    .B2(_03834_),
    .C1(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__inv_2 _09075_ (.A(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__or2_1 _09076_ (.A(_03788_),
    .B(_03837_),
    .X(_03838_));
 sky130_fd_sc_hd__or2_1 _09077_ (.A(_03786_),
    .B(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__clkbuf_2 _09078_ (.A(_03839_),
    .X(_03840_));
 sky130_fd_sc_hd__a32o_1 _09079_ (.A1(_03737_),
    .A2(_03751_),
    .A3(_03778_),
    .B1(_03840_),
    .B2(_03758_),
    .X(_00057_));
 sky130_fd_sc_hd__buf_2 _09080_ (.A(_03229_),
    .X(_03841_));
 sky130_fd_sc_hd__nor2_1 _09081_ (.A(_03841_),
    .B(_03237_),
    .Y(_03842_));
 sky130_fd_sc_hd__and2_1 _09082_ (.A(_03743_),
    .B(_03781_),
    .X(_03843_));
 sky130_fd_sc_hd__clkbuf_4 _09083_ (.A(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__and2_2 _09084_ (.A(_03739_),
    .B(_03844_),
    .X(_03845_));
 sky130_fd_sc_hd__clkbuf_4 _09085_ (.A(_03757_),
    .X(_03846_));
 sky130_fd_sc_hd__mux2_1 _09086_ (.A0(\mem_rdata_q[7] ),
    .A1(_03822_),
    .S(_03846_),
    .X(_03847_));
 sky130_fd_sc_hd__o211ai_4 _09087_ (.A1(_03783_),
    .A2(_03748_),
    .B1(_03835_),
    .C1(_03844_),
    .Y(_03848_));
 sky130_fd_sc_hd__a32o_1 _09088_ (.A1(_03842_),
    .A2(_03737_),
    .A3(_03845_),
    .B1(_03847_),
    .B2(_03848_),
    .X(_00058_));
 sky130_fd_sc_hd__clkbuf_4 _09089_ (.A(_03753_),
    .X(_03849_));
 sky130_fd_sc_hd__clkbuf_4 _09090_ (.A(_03754_),
    .X(_03850_));
 sky130_fd_sc_hd__a22o_1 _09091_ (.A1(_03849_),
    .A2(_03801_),
    .B1(_03802_),
    .B2(_03850_),
    .X(_03851_));
 sky130_fd_sc_hd__mux2_1 _09092_ (.A0(\mem_rdata_q[20] ),
    .A1(_03851_),
    .S(_03846_),
    .X(_03852_));
 sky130_fd_sc_hd__nor2_2 _09093_ (.A(_03767_),
    .B(_03768_),
    .Y(_03853_));
 sky130_fd_sc_hd__or2_2 _09094_ (.A(_03750_),
    .B(_03844_),
    .X(_03854_));
 sky130_fd_sc_hd__nor2_1 _09095_ (.A(_03738_),
    .B(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__or2_1 _09096_ (.A(_03816_),
    .B(_03770_),
    .X(_03856_));
 sky130_fd_sc_hd__a21o_1 _09097_ (.A1(_03743_),
    .A2(_03782_),
    .B1(_03853_),
    .X(_03857_));
 sky130_fd_sc_hd__a31o_1 _09098_ (.A1(_03834_),
    .A2(_03856_),
    .A3(_03857_),
    .B1(_03789_),
    .X(_03858_));
 sky130_fd_sc_hd__nand2_1 _09099_ (.A(_03835_),
    .B(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__or4_1 _09100_ (.A(_03785_),
    .B(_03788_),
    .C(_03845_),
    .D(_03859_),
    .X(_03860_));
 sky130_fd_sc_hd__a31o_1 _09101_ (.A1(_03853_),
    .A2(_03776_),
    .A3(_03855_),
    .B1(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__clkbuf_4 _09102_ (.A(_03782_),
    .X(_03862_));
 sky130_fd_sc_hd__nor2_1 _09103_ (.A(_03770_),
    .B(_03776_),
    .Y(_03863_));
 sky130_fd_sc_hd__clkbuf_4 _09104_ (.A(_03814_),
    .X(_03864_));
 sky130_fd_sc_hd__o21a_1 _09105_ (.A1(_03862_),
    .A2(_03863_),
    .B1(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__or3b_1 _09106_ (.A(_03780_),
    .B(_03748_),
    .C_N(_03743_),
    .X(_03866_));
 sky130_fd_sc_hd__clkbuf_4 _09107_ (.A(_03832_),
    .X(_03867_));
 sky130_fd_sc_hd__or2b_1 _09108_ (.A(_03827_),
    .B_N(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__and2b_2 _09109_ (.A_N(_03866_),
    .B(_03868_),
    .X(_03869_));
 sky130_fd_sc_hd__and2_1 _09110_ (.A(_03736_),
    .B(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__or2_1 _09111_ (.A(_03865_),
    .B(_03870_),
    .X(_03871_));
 sky130_fd_sc_hd__a22o_1 _09112_ (.A1(_03852_),
    .A2(_03861_),
    .B1(_03871_),
    .B2(_03855_),
    .X(_00046_));
 sky130_fd_sc_hd__o21a_1 _09113_ (.A1(_03862_),
    .A2(_03863_),
    .B1(_03810_),
    .X(_03872_));
 sky130_fd_sc_hd__or2_1 _09114_ (.A(_03870_),
    .B(_03872_),
    .X(_03873_));
 sky130_fd_sc_hd__a22o_1 _09115_ (.A1(_03850_),
    .A2(_03791_),
    .B1(_03792_),
    .B2(_03849_),
    .X(_03874_));
 sky130_fd_sc_hd__mux2_1 _09116_ (.A0(\mem_rdata_q[21] ),
    .A1(_03874_),
    .S(_03846_),
    .X(_03875_));
 sky130_fd_sc_hd__a22o_1 _09117_ (.A1(_03855_),
    .A2(_03873_),
    .B1(_03875_),
    .B2(_03861_),
    .X(_00047_));
 sky130_fd_sc_hd__a22o_1 _09118_ (.A1(_03850_),
    .A2(_03795_),
    .B1(_03796_),
    .B2(_03849_),
    .X(_03876_));
 sky130_fd_sc_hd__mux2_1 _09119_ (.A0(\mem_rdata_q[22] ),
    .A1(_03876_),
    .S(_03846_),
    .X(_03877_));
 sky130_fd_sc_hd__clkbuf_4 _09120_ (.A(_03798_),
    .X(_03878_));
 sky130_fd_sc_hd__nor2_2 _09121_ (.A(_03783_),
    .B(_03213_),
    .Y(_03879_));
 sky130_fd_sc_hd__and2_2 _09122_ (.A(_03862_),
    .B(_03879_),
    .X(_03880_));
 sky130_fd_sc_hd__and2b_1 _09123_ (.A_N(_03854_),
    .B(_03870_),
    .X(_03881_));
 sky130_fd_sc_hd__nor2_1 _09124_ (.A(_03779_),
    .B(_03789_),
    .Y(_03882_));
 sky130_fd_sc_hd__a22o_1 _09125_ (.A1(_03862_),
    .A2(_03739_),
    .B1(_03882_),
    .B2(_03767_),
    .X(_03883_));
 sky130_fd_sc_hd__and2b_1 _09126_ (.A_N(_03854_),
    .B(_03863_),
    .X(_03884_));
 sky130_fd_sc_hd__clkbuf_4 _09127_ (.A(_03804_),
    .X(_03885_));
 sky130_fd_sc_hd__o21a_1 _09128_ (.A1(_03883_),
    .A2(_03884_),
    .B1(_03885_),
    .X(_03886_));
 sky130_fd_sc_hd__a211o_1 _09129_ (.A1(_03878_),
    .A2(_03880_),
    .B1(_03881_),
    .C1(_03886_),
    .X(_03887_));
 sky130_fd_sc_hd__clkbuf_4 _09130_ (.A(_03835_),
    .X(_03888_));
 sky130_fd_sc_hd__a22o_1 _09131_ (.A1(_03861_),
    .A2(_03877_),
    .B1(_03887_),
    .B2(_03888_),
    .X(_00048_));
 sky130_fd_sc_hd__a22o_1 _09132_ (.A1(_03850_),
    .A2(_03819_),
    .B1(_03820_),
    .B2(_03849_),
    .X(_03889_));
 sky130_fd_sc_hd__mux2_1 _09133_ (.A0(\mem_rdata_q[23] ),
    .A1(_03889_),
    .S(_03846_),
    .X(_03890_));
 sky130_fd_sc_hd__clkbuf_4 _09134_ (.A(_03743_),
    .X(_03891_));
 sky130_fd_sc_hd__clkbuf_4 _09135_ (.A(_03774_),
    .X(_03892_));
 sky130_fd_sc_hd__nand2_1 _09136_ (.A(_03862_),
    .B(_03879_),
    .Y(_03893_));
 sky130_fd_sc_hd__nor2_2 _09137_ (.A(_03891_),
    .B(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__buf_4 _09138_ (.A(_03794_),
    .X(_03895_));
 sky130_fd_sc_hd__o21a_1 _09139_ (.A1(_03883_),
    .A2(_03894_),
    .B1(_03895_),
    .X(_03896_));
 sky130_fd_sc_hd__a31o_1 _09140_ (.A1(_03891_),
    .A2(_03892_),
    .A3(_03880_),
    .B1(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__a21o_1 _09141_ (.A1(_03895_),
    .A2(_03863_),
    .B1(_03870_),
    .X(_03898_));
 sky130_fd_sc_hd__a22o_1 _09142_ (.A1(_03835_),
    .A2(_03897_),
    .B1(_03898_),
    .B2(_03855_),
    .X(_03899_));
 sky130_fd_sc_hd__a21o_1 _09143_ (.A1(_03861_),
    .A2(_03890_),
    .B1(_03899_),
    .X(_00049_));
 sky130_fd_sc_hd__a22o_1 _09144_ (.A1(_03850_),
    .A2(_03828_),
    .B1(_03830_),
    .B2(_03849_),
    .X(_03900_));
 sky130_fd_sc_hd__mux2_1 _09145_ (.A0(\mem_rdata_q[24] ),
    .A1(_03900_),
    .S(_03846_),
    .X(_03901_));
 sky130_fd_sc_hd__or2_2 _09146_ (.A(_03868_),
    .B(_03866_),
    .X(_03902_));
 sky130_fd_sc_hd__nor2_1 _09147_ (.A(_03854_),
    .B(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hd__o31a_1 _09148_ (.A1(_03883_),
    .A2(_03884_),
    .A3(_03903_),
    .B1(_03878_),
    .X(_03904_));
 sky130_fd_sc_hd__a211o_1 _09149_ (.A1(_03763_),
    .A2(_03880_),
    .B1(_03881_),
    .C1(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__a22o_1 _09150_ (.A1(_03861_),
    .A2(_03901_),
    .B1(_03905_),
    .B2(_03888_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _09151_ (.A0(\mem_rdata_q[15] ),
    .A1(_03781_),
    .S(_03846_),
    .X(_03906_));
 sky130_fd_sc_hd__and3_1 _09152_ (.A(_03739_),
    .B(_03842_),
    .C(_03869_),
    .X(_03907_));
 sky130_fd_sc_hd__clkbuf_2 _09153_ (.A(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__mux2_1 _09154_ (.A0(_03906_),
    .A1(_03895_),
    .S(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__clkbuf_1 _09155_ (.A(_03909_),
    .X(_00041_));
 sky130_fd_sc_hd__a22o_1 _09156_ (.A1(_03849_),
    .A2(_03201_),
    .B1(_03202_),
    .B2(_03850_),
    .X(_03910_));
 sky130_fd_sc_hd__mux2_1 _09157_ (.A0(\mem_rdata_q[16] ),
    .A1(_03910_),
    .S(_03846_),
    .X(_03911_));
 sky130_fd_sc_hd__mux2_1 _09158_ (.A0(_03911_),
    .A1(_03878_),
    .S(_03908_),
    .X(_03912_));
 sky130_fd_sc_hd__clkbuf_1 _09159_ (.A(_03912_),
    .X(_00042_));
 sky130_fd_sc_hd__a22o_1 _09160_ (.A1(_03849_),
    .A2(_03209_),
    .B1(_03210_),
    .B2(_03850_),
    .X(_03913_));
 sky130_fd_sc_hd__buf_4 _09161_ (.A(_03846_),
    .X(_03914_));
 sky130_fd_sc_hd__mux2_1 _09162_ (.A0(\mem_rdata_q[17] ),
    .A1(_03913_),
    .S(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__clkbuf_4 _09163_ (.A(_03818_),
    .X(_03916_));
 sky130_fd_sc_hd__nand2_1 _09164_ (.A(_03916_),
    .B(_03908_),
    .Y(_03917_));
 sky130_fd_sc_hd__o21a_1 _09165_ (.A1(_03908_),
    .A2(_03915_),
    .B1(_03917_),
    .X(_00043_));
 sky130_fd_sc_hd__a22o_1 _09166_ (.A1(_03850_),
    .A2(_03811_),
    .B1(_03812_),
    .B2(_03849_),
    .X(_03918_));
 sky130_fd_sc_hd__mux2_1 _09167_ (.A0(\mem_rdata_q[18] ),
    .A1(_03918_),
    .S(_03914_),
    .X(_03919_));
 sky130_fd_sc_hd__o21a_1 _09168_ (.A1(_03908_),
    .A2(_03919_),
    .B1(_03917_),
    .X(_00044_));
 sky130_fd_sc_hd__a22o_1 _09169_ (.A1(_03849_),
    .A2(_03807_),
    .B1(_03805_),
    .B2(_03850_),
    .X(_03920_));
 sky130_fd_sc_hd__mux2_1 _09170_ (.A0(\mem_rdata_q[19] ),
    .A1(_03920_),
    .S(_03914_),
    .X(_03921_));
 sky130_fd_sc_hd__o21a_1 _09171_ (.A1(_03908_),
    .A2(_03921_),
    .B1(_03917_),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_1 _09172_ (.A0(\mem_rdata_q[12] ),
    .A1(_03736_),
    .S(_03757_),
    .X(_03922_));
 sky130_fd_sc_hd__nor2_2 _09173_ (.A(_03781_),
    .B(_03768_),
    .Y(_03923_));
 sky130_fd_sc_hd__a21o_1 _09174_ (.A1(_03864_),
    .A2(_03868_),
    .B1(_03781_),
    .X(_03924_));
 sky130_fd_sc_hd__nand2_1 _09175_ (.A(_03762_),
    .B(_03892_),
    .Y(_03925_));
 sky130_fd_sc_hd__nor2_1 _09176_ (.A(_03736_),
    .B(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__nor2_2 _09177_ (.A(_03770_),
    .B(_03926_),
    .Y(_03927_));
 sky130_fd_sc_hd__a21o_1 _09178_ (.A1(_03798_),
    .A2(_03853_),
    .B1(_03927_),
    .X(_03928_));
 sky130_fd_sc_hd__or3_1 _09179_ (.A(_03916_),
    .B(_03922_),
    .C(_03925_),
    .X(_03929_));
 sky130_fd_sc_hd__o211a_1 _09180_ (.A1(_03895_),
    .A2(_03927_),
    .B1(_03928_),
    .C1(_03929_),
    .X(_03930_));
 sky130_fd_sc_hd__a31o_1 _09181_ (.A1(_03891_),
    .A2(_03747_),
    .A3(_03924_),
    .B1(_03930_),
    .X(_03931_));
 sky130_fd_sc_hd__and2_2 _09182_ (.A(_03739_),
    .B(_03749_),
    .X(_03932_));
 sky130_fd_sc_hd__a22o_1 _09183_ (.A1(_03790_),
    .A2(_03923_),
    .B1(_03931_),
    .B2(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__a22o_1 _09184_ (.A1(_03840_),
    .A2(_03922_),
    .B1(_03933_),
    .B2(_03888_),
    .X(_00038_));
 sky130_fd_sc_hd__mux2_1 _09185_ (.A0(\mem_rdata_q[13] ),
    .A1(_03747_),
    .S(_03227_),
    .X(_03934_));
 sky130_fd_sc_hd__nor2_2 _09186_ (.A(_03783_),
    .B(_03779_),
    .Y(_03935_));
 sky130_fd_sc_hd__or3_1 _09187_ (.A(_03775_),
    .B(_03916_),
    .C(_03934_),
    .X(_03936_));
 sky130_fd_sc_hd__a32o_1 _09188_ (.A1(_03763_),
    .A2(_03928_),
    .A3(_03936_),
    .B1(_03869_),
    .B2(_03810_),
    .X(_03937_));
 sky130_fd_sc_hd__a22o_1 _09189_ (.A1(_03785_),
    .A2(_03934_),
    .B1(_03937_),
    .B2(_03932_),
    .X(_03938_));
 sky130_fd_sc_hd__or2_1 _09190_ (.A(_03935_),
    .B(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__a22o_1 _09191_ (.A1(_03838_),
    .A2(_03934_),
    .B1(_03939_),
    .B2(_03888_),
    .X(_00039_));
 sky130_fd_sc_hd__clkbuf_4 _09192_ (.A(\mem_rdata_q[14] ),
    .X(_03940_));
 sky130_fd_sc_hd__mux2_1 _09193_ (.A0(_03940_),
    .A1(_03891_),
    .S(_03757_),
    .X(_03941_));
 sky130_fd_sc_hd__nand2_1 _09194_ (.A(_03799_),
    .B(_03926_),
    .Y(_03942_));
 sky130_fd_sc_hd__or3_1 _09195_ (.A(_03916_),
    .B(_03925_),
    .C(_03941_),
    .X(_03943_));
 sky130_fd_sc_hd__a32o_1 _09196_ (.A1(_03853_),
    .A2(_03942_),
    .A3(_03943_),
    .B1(_03869_),
    .B2(_03885_),
    .X(_03944_));
 sky130_fd_sc_hd__a22o_1 _09197_ (.A1(_03840_),
    .A2(_03941_),
    .B1(_03944_),
    .B2(_03751_),
    .X(_00040_));
 sky130_fd_sc_hd__o211a_1 _09198_ (.A1(_03730_),
    .A2(_03867_),
    .B1(_03848_),
    .C1(_03829_),
    .X(_03945_));
 sky130_fd_sc_hd__a31o_1 _09199_ (.A1(_03842_),
    .A2(_03810_),
    .A3(_03845_),
    .B1(_03945_),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _09200_ (.A0(\mem_rdata_q[9] ),
    .A1(_03826_),
    .S(_03846_),
    .X(_03946_));
 sky130_fd_sc_hd__or2_1 _09201_ (.A(_03779_),
    .B(_03789_),
    .X(_03947_));
 sky130_fd_sc_hd__nor2_1 _09202_ (.A(_03767_),
    .B(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__and4_1 _09203_ (.A(_03748_),
    .B(_03879_),
    .C(_03878_),
    .D(_03844_),
    .X(_03949_));
 sky130_fd_sc_hd__a221o_1 _09204_ (.A1(_03885_),
    .A2(_03845_),
    .B1(_03948_),
    .B2(_03826_),
    .C1(_03949_),
    .X(_03950_));
 sky130_fd_sc_hd__a22o_1 _09205_ (.A1(_03848_),
    .A2(_03946_),
    .B1(_03950_),
    .B2(_03888_),
    .X(_00060_));
 sky130_fd_sc_hd__nand2_1 _09206_ (.A(_03730_),
    .B(_03848_),
    .Y(_03951_));
 sky130_fd_sc_hd__mux2_1 _09207_ (.A0(\mem_rdata_q[10] ),
    .A1(_03892_),
    .S(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__clkbuf_1 _09208_ (.A(_03952_),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _09209_ (.A0(\mem_rdata_q[11] ),
    .A1(_03763_),
    .S(_03951_),
    .X(_03953_));
 sky130_fd_sc_hd__clkbuf_1 _09210_ (.A(_03953_),
    .X(_00037_));
 sky130_fd_sc_hd__a22o_2 _09211_ (.A1(_03753_),
    .A2(_03823_),
    .B1(_03824_),
    .B2(_03754_),
    .X(_03954_));
 sky130_fd_sc_hd__mux2_1 _09212_ (.A0(\mem_rdata_q[25] ),
    .A1(_03954_),
    .S(_03757_),
    .X(_03955_));
 sky130_fd_sc_hd__or2_1 _09213_ (.A(_03935_),
    .B(_03880_),
    .X(_03956_));
 sky130_fd_sc_hd__o21a_1 _09214_ (.A1(_03782_),
    .A2(_03869_),
    .B1(_03736_),
    .X(_03957_));
 sky130_fd_sc_hd__or2b_1 _09215_ (.A(_03843_),
    .B_N(_03902_),
    .X(_03958_));
 sky130_fd_sc_hd__and2_1 _09216_ (.A(_03762_),
    .B(_03892_),
    .X(_03959_));
 sky130_fd_sc_hd__nor2_2 _09217_ (.A(_03818_),
    .B(_03776_),
    .Y(_03960_));
 sky130_fd_sc_hd__a21o_1 _09218_ (.A1(_03959_),
    .A2(_03955_),
    .B1(_03960_),
    .X(_03961_));
 sky130_fd_sc_hd__a22o_1 _09219_ (.A1(_03864_),
    .A2(_03958_),
    .B1(_03961_),
    .B2(_03927_),
    .X(_03962_));
 sky130_fd_sc_hd__o21a_1 _09220_ (.A1(_03957_),
    .A2(_03962_),
    .B1(_03932_),
    .X(_03963_));
 sky130_fd_sc_hd__a221o_1 _09221_ (.A1(_03786_),
    .A2(_03955_),
    .B1(_03956_),
    .B2(_03737_),
    .C1(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__a22o_1 _09222_ (.A1(_03838_),
    .A2(_03955_),
    .B1(_03964_),
    .B2(_03888_),
    .X(_00051_));
 sky130_fd_sc_hd__a22o_2 _09223_ (.A1(_03754_),
    .A2(_03771_),
    .B1(_03772_),
    .B2(_03753_),
    .X(_03965_));
 sky130_fd_sc_hd__mux2_2 _09224_ (.A0(\mem_rdata_q[26] ),
    .A1(_03965_),
    .S(_03757_),
    .X(_03966_));
 sky130_fd_sc_hd__a21o_1 _09225_ (.A1(_03959_),
    .A2(_03966_),
    .B1(_03960_),
    .X(_03967_));
 sky130_fd_sc_hd__or2b_1 _09226_ (.A(_03957_),
    .B_N(_03749_),
    .X(_03968_));
 sky130_fd_sc_hd__a221o_1 _09227_ (.A1(_03895_),
    .A2(_03958_),
    .B1(_03967_),
    .B2(_03927_),
    .C1(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__o211a_1 _09228_ (.A1(_03749_),
    .A2(_03966_),
    .B1(_03969_),
    .C1(_03739_),
    .X(_03970_));
 sky130_fd_sc_hd__nor2_1 _09229_ (.A(_03779_),
    .B(_03784_),
    .Y(_03971_));
 sky130_fd_sc_hd__or2_1 _09230_ (.A(_03894_),
    .B(_03948_),
    .X(_03972_));
 sky130_fd_sc_hd__a32o_1 _09231_ (.A1(_03862_),
    .A2(_03864_),
    .A3(_03882_),
    .B1(_03966_),
    .B2(_03786_),
    .X(_03973_));
 sky130_fd_sc_hd__a221o_1 _09232_ (.A1(_03895_),
    .A2(_03971_),
    .B1(_03972_),
    .B2(_03822_),
    .C1(_03973_),
    .X(_03974_));
 sky130_fd_sc_hd__or2_1 _09233_ (.A(_03970_),
    .B(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__a22o_1 _09234_ (.A1(_03837_),
    .A2(_03966_),
    .B1(_03975_),
    .B2(_03888_),
    .X(_00052_));
 sky130_fd_sc_hd__or2_1 _09235_ (.A(_03786_),
    .B(_03837_),
    .X(_03976_));
 sky130_fd_sc_hd__a22o_2 _09236_ (.A1(_03754_),
    .A2(_03759_),
    .B1(_03760_),
    .B2(_03753_),
    .X(_03977_));
 sky130_fd_sc_hd__mux2_1 _09237_ (.A0(\mem_rdata_q[27] ),
    .A1(_03977_),
    .S(_03227_),
    .X(_03978_));
 sky130_fd_sc_hd__a31o_2 _09238_ (.A1(_03728_),
    .A2(_03806_),
    .A3(_03808_),
    .B1(_03809_),
    .X(_03979_));
 sky130_fd_sc_hd__a21o_1 _09239_ (.A1(_03959_),
    .A2(_03978_),
    .B1(_03960_),
    .X(_03980_));
 sky130_fd_sc_hd__a2bb2o_1 _09240_ (.A1_N(_03979_),
    .A2_N(_03902_),
    .B1(_03927_),
    .B2(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__a211o_1 _09241_ (.A1(_03878_),
    .A2(_03844_),
    .B1(_03968_),
    .C1(_03981_),
    .X(_03982_));
 sky130_fd_sc_hd__o211a_1 _09242_ (.A1(_03749_),
    .A2(_03978_),
    .B1(_03982_),
    .C1(_03739_),
    .X(_03983_));
 sky130_fd_sc_hd__a32o_1 _09243_ (.A1(_03891_),
    .A2(_03862_),
    .A3(_03810_),
    .B1(_03867_),
    .B2(_03844_),
    .X(_03984_));
 sky130_fd_sc_hd__and3_1 _09244_ (.A(_03748_),
    .B(_03790_),
    .C(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__a311o_1 _09245_ (.A1(_03879_),
    .A2(_03867_),
    .A3(_03923_),
    .B1(_03983_),
    .C1(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__a22o_1 _09246_ (.A1(_03976_),
    .A2(_03978_),
    .B1(_03986_),
    .B2(_03888_),
    .X(_00053_));
 sky130_fd_sc_hd__a22o_2 _09247_ (.A1(_03754_),
    .A2(_03733_),
    .B1(_03731_),
    .B2(_03753_),
    .X(_03987_));
 sky130_fd_sc_hd__mux2_1 _09248_ (.A0(\mem_rdata_q[28] ),
    .A1(_03987_),
    .S(_03757_),
    .X(_03988_));
 sky130_fd_sc_hd__and2b_1 _09249_ (.A_N(_03902_),
    .B(_03885_),
    .X(_03989_));
 sky130_fd_sc_hd__a21o_1 _09250_ (.A1(_03959_),
    .A2(_03988_),
    .B1(_03960_),
    .X(_03990_));
 sky130_fd_sc_hd__a22o_1 _09251_ (.A1(_03737_),
    .A2(_03844_),
    .B1(_03927_),
    .B2(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__o31a_1 _09252_ (.A1(_03957_),
    .A2(_03989_),
    .A3(_03991_),
    .B1(_03932_),
    .X(_03992_));
 sky130_fd_sc_hd__a221o_1 _09253_ (.A1(_03826_),
    .A2(_03894_),
    .B1(_03988_),
    .B2(_03786_),
    .C1(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__a22o_1 _09254_ (.A1(_03838_),
    .A2(_03988_),
    .B1(_03993_),
    .B2(_03888_),
    .X(_00054_));
 sky130_fd_sc_hd__a22o_2 _09255_ (.A1(_03754_),
    .A2(_03744_),
    .B1(_03745_),
    .B2(_03753_),
    .X(_03994_));
 sky130_fd_sc_hd__mux2_1 _09256_ (.A0(\mem_rdata_q[29] ),
    .A1(_03994_),
    .S(_03757_),
    .X(_03995_));
 sky130_fd_sc_hd__or2_1 _09257_ (.A(_03891_),
    .B(_03862_),
    .X(_03996_));
 sky130_fd_sc_hd__o21a_1 _09258_ (.A1(_03775_),
    .A2(_03995_),
    .B1(_03763_),
    .X(_03997_));
 sky130_fd_sc_hd__o211a_1 _09259_ (.A1(_03996_),
    .A2(_03997_),
    .B1(_03737_),
    .C1(_03932_),
    .X(_03998_));
 sky130_fd_sc_hd__a21o_1 _09260_ (.A1(_03892_),
    .A2(_03894_),
    .B1(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__a22o_1 _09261_ (.A1(_03840_),
    .A2(_03995_),
    .B1(_03999_),
    .B2(_03888_),
    .X(_00055_));
 sky130_fd_sc_hd__a22o_2 _09262_ (.A1(_03753_),
    .A2(_03740_),
    .B1(_03741_),
    .B2(_03850_),
    .X(_04000_));
 sky130_fd_sc_hd__mux2_1 _09263_ (.A0(\mem_rdata_q[30] ),
    .A1(_04000_),
    .S(_03757_),
    .X(_04001_));
 sky130_fd_sc_hd__a21bo_1 _09264_ (.A1(_03737_),
    .A2(_04001_),
    .B1_N(_03763_),
    .X(_04002_));
 sky130_fd_sc_hd__inv_2 _09265_ (.A(_03942_),
    .Y(_04003_));
 sky130_fd_sc_hd__a211o_1 _09266_ (.A1(_03892_),
    .A2(_04002_),
    .B1(_03960_),
    .C1(_04003_),
    .X(_04004_));
 sky130_fd_sc_hd__a22o_1 _09267_ (.A1(_03737_),
    .A2(_03996_),
    .B1(_04004_),
    .B2(_03853_),
    .X(_04005_));
 sky130_fd_sc_hd__a22o_1 _09268_ (.A1(_03840_),
    .A2(_04001_),
    .B1(_04005_),
    .B2(_03751_),
    .X(_00056_));
 sky130_fd_sc_hd__or3_4 _09269_ (.A(\cpu_state[3] ),
    .B(\cpu_state[6] ),
    .C(_03410_),
    .X(_04006_));
 sky130_fd_sc_hd__clkbuf_4 _09270_ (.A(_04006_),
    .X(_04007_));
 sky130_fd_sc_hd__clkbuf_4 _09271_ (.A(_04007_),
    .X(_04008_));
 sky130_fd_sc_hd__buf_4 _09272_ (.A(_03252_),
    .X(_04009_));
 sky130_fd_sc_hd__clkbuf_4 _09273_ (.A(_04009_),
    .X(_04010_));
 sky130_fd_sc_hd__clkbuf_4 _09274_ (.A(instr_rdinstr),
    .X(_04011_));
 sky130_fd_sc_hd__clkbuf_4 _09275_ (.A(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__clkbuf_4 _09276_ (.A(_03253_),
    .X(_04013_));
 sky130_fd_sc_hd__buf_4 _09277_ (.A(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__clkbuf_4 _09278_ (.A(instr_rdinstrh),
    .X(_04015_));
 sky130_fd_sc_hd__buf_4 _09279_ (.A(_04015_),
    .X(_04016_));
 sky130_fd_sc_hd__clkbuf_4 _09280_ (.A(instr_rdcycleh),
    .X(_04017_));
 sky130_fd_sc_hd__buf_4 _09281_ (.A(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__a22o_1 _09282_ (.A1(\count_instr[32] ),
    .A2(_04016_),
    .B1(_04018_),
    .B2(\count_cycle[32] ),
    .X(_04019_));
 sky130_fd_sc_hd__a221o_1 _09283_ (.A1(\count_instr[0] ),
    .A2(_04012_),
    .B1(\count_cycle[0] ),
    .B2(_04014_),
    .C1(_04019_),
    .X(_04020_));
 sky130_fd_sc_hd__clkbuf_4 _09284_ (.A(instr_maskirq),
    .X(_04021_));
 sky130_fd_sc_hd__clkbuf_8 _09285_ (.A(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__clkbuf_4 _09286_ (.A(instr_timer),
    .X(_04023_));
 sky130_fd_sc_hd__clkbuf_4 _09287_ (.A(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__nor3_2 _09288_ (.A(instr_timer),
    .B(instr_maskirq),
    .C(instr_retirq),
    .Y(_04025_));
 sky130_fd_sc_hd__clkbuf_4 _09289_ (.A(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__clkbuf_4 _09290_ (.A(_04026_),
    .X(_04027_));
 sky130_fd_sc_hd__a221o_1 _09291_ (.A1(\irq_mask[0] ),
    .A2(_04022_),
    .B1(\timer[0] ),
    .B2(_04024_),
    .C1(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__o211a_1 _09292_ (.A1(_04010_),
    .A2(_04020_),
    .B1(_04028_),
    .C1(_03303_),
    .X(_04029_));
 sky130_fd_sc_hd__nand2_4 _09293_ (.A(_03242_),
    .B(\mem_wordsize[2] ),
    .Y(_04030_));
 sky130_fd_sc_hd__or2b_1 _09294_ (.A(\mem_wordsize[2] ),
    .B_N(\mem_wordsize[1] ),
    .X(_04031_));
 sky130_fd_sc_hd__a21bo_1 _09295_ (.A1(_04030_),
    .A2(_04031_),
    .B1_N(_03243_),
    .X(_04032_));
 sky130_fd_sc_hd__buf_4 _09296_ (.A(_04032_),
    .X(net258));
 sky130_fd_sc_hd__inv_2 _09297_ (.A(net67),
    .Y(_04033_));
 sky130_fd_sc_hd__o21a_2 _09298_ (.A1(\mem_wordsize[2] ),
    .A2(\mem_wordsize[1] ),
    .B1(_03242_),
    .X(_04034_));
 sky130_fd_sc_hd__o21a_2 _09299_ (.A1(_04033_),
    .A2(\mem_wordsize[2] ),
    .B1(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__clkbuf_4 _09300_ (.A(net67),
    .X(_04036_));
 sky130_fd_sc_hd__clkbuf_4 _09301_ (.A(_04036_),
    .X(_04037_));
 sky130_fd_sc_hd__clkbuf_4 _09302_ (.A(\mem_wordsize[1] ),
    .X(_04038_));
 sky130_fd_sc_hd__clkbuf_4 _09303_ (.A(_03242_),
    .X(_04039_));
 sky130_fd_sc_hd__buf_4 _09304_ (.A(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__mux2_1 _09305_ (.A0(net63),
    .A1(net49),
    .S(_04040_),
    .X(_04041_));
 sky130_fd_sc_hd__and3_1 _09306_ (.A(_04037_),
    .B(_04038_),
    .C(_04041_),
    .X(_04042_));
 sky130_fd_sc_hd__a221o_1 _09307_ (.A1(net33),
    .A2(net258),
    .B1(_04035_),
    .B2(net40),
    .C1(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__or2_1 _09308_ (.A(\reg_next_pc[0] ),
    .B(\decoded_imm[0] ),
    .X(_04044_));
 sky130_fd_sc_hd__nand2_1 _09309_ (.A(\reg_next_pc[0] ),
    .B(\decoded_imm[0] ),
    .Y(_04045_));
 sky130_fd_sc_hd__buf_4 _09310_ (.A(_03312_),
    .X(_04046_));
 sky130_fd_sc_hd__a32o_1 _09311_ (.A1(\cpu_state[3] ),
    .A2(_04044_),
    .A3(_04045_),
    .B1(_04037_),
    .B2(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__nor3_2 _09312_ (.A(\cpu_state[3] ),
    .B(\cpu_state[6] ),
    .C(_03410_),
    .Y(_04048_));
 sky130_fd_sc_hd__buf_4 _09313_ (.A(_04048_),
    .X(_04049_));
 sky130_fd_sc_hd__a211o_2 _09314_ (.A1(_03226_),
    .A2(_04043_),
    .B1(_04047_),
    .C1(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__o22a_1 _09315_ (.A1(\irq_pending[0] ),
    .A2(_04008_),
    .B1(_04029_),
    .B2(_04050_),
    .X(_08369_));
 sky130_fd_sc_hd__inv_2 _09316_ (.A(instr_retirq),
    .Y(_04051_));
 sky130_fd_sc_hd__buf_4 _09317_ (.A(_00072_),
    .X(_04052_));
 sky130_fd_sc_hd__clkbuf_8 _09318_ (.A(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__clkbuf_8 _09319_ (.A(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__clkbuf_8 _09320_ (.A(_00069_),
    .X(_04055_));
 sky130_fd_sc_hd__buf_6 _09321_ (.A(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__buf_8 _09322_ (.A(_04056_),
    .X(_04057_));
 sky130_fd_sc_hd__clkbuf_8 _09323_ (.A(_00070_),
    .X(_04058_));
 sky130_fd_sc_hd__clkbuf_8 _09324_ (.A(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__clkbuf_8 _09325_ (.A(_04059_),
    .X(_04060_));
 sky130_fd_sc_hd__mux4_1 _09326_ (.A0(\cpuregs.regs[28][1] ),
    .A1(\cpuregs.regs[29][1] ),
    .A2(\cpuregs.regs[30][1] ),
    .A3(\cpuregs.regs[31][1] ),
    .S0(_04057_),
    .S1(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__mux4_1 _09327_ (.A0(\cpuregs.regs[24][1] ),
    .A1(\cpuregs.regs[25][1] ),
    .A2(\cpuregs.regs[26][1] ),
    .A3(\cpuregs.regs[27][1] ),
    .S0(_04057_),
    .S1(_04060_),
    .X(_04062_));
 sky130_fd_sc_hd__clkinv_4 _09328_ (.A(_00071_),
    .Y(_04063_));
 sky130_fd_sc_hd__buf_8 _09329_ (.A(_04063_),
    .X(_04064_));
 sky130_fd_sc_hd__buf_8 _09330_ (.A(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__mux2_1 _09331_ (.A0(_04061_),
    .A1(_04062_),
    .S(_04065_),
    .X(_04066_));
 sky130_fd_sc_hd__nand2_1 _09332_ (.A(_04054_),
    .B(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__inv_6 _09333_ (.A(_00072_),
    .Y(_04068_));
 sky130_fd_sc_hd__buf_6 _09334_ (.A(_04068_),
    .X(_04069_));
 sky130_fd_sc_hd__buf_4 _09335_ (.A(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__clkbuf_8 _09336_ (.A(_00069_),
    .X(_04071_));
 sky130_fd_sc_hd__buf_6 _09337_ (.A(_04071_),
    .X(_04072_));
 sky130_fd_sc_hd__buf_4 _09338_ (.A(_00070_),
    .X(_04073_));
 sky130_fd_sc_hd__clkbuf_8 _09339_ (.A(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__mux4_1 _09340_ (.A0(\cpuregs.regs[20][1] ),
    .A1(\cpuregs.regs[21][1] ),
    .A2(\cpuregs.regs[22][1] ),
    .A3(\cpuregs.regs[23][1] ),
    .S0(_04072_),
    .S1(_04074_),
    .X(_04075_));
 sky130_fd_sc_hd__mux4_1 _09341_ (.A0(\cpuregs.regs[16][1] ),
    .A1(\cpuregs.regs[17][1] ),
    .A2(\cpuregs.regs[18][1] ),
    .A3(\cpuregs.regs[19][1] ),
    .S0(_04072_),
    .S1(_04074_),
    .X(_04076_));
 sky130_fd_sc_hd__buf_6 _09342_ (.A(_04063_),
    .X(_04077_));
 sky130_fd_sc_hd__buf_6 _09343_ (.A(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__mux2_1 _09344_ (.A0(_04075_),
    .A1(_04076_),
    .S(_04078_),
    .X(_04079_));
 sky130_fd_sc_hd__inv_2 _09345_ (.A(_00073_),
    .Y(_04080_));
 sky130_fd_sc_hd__clkbuf_8 _09346_ (.A(_04080_),
    .X(_04081_));
 sky130_fd_sc_hd__clkbuf_8 _09347_ (.A(_04081_),
    .X(_04082_));
 sky130_fd_sc_hd__a21oi_1 _09348_ (.A1(_04070_),
    .A2(_04079_),
    .B1(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__buf_8 _09349_ (.A(_00069_),
    .X(_04084_));
 sky130_fd_sc_hd__buf_8 _09350_ (.A(_04084_),
    .X(_04085_));
 sky130_fd_sc_hd__buf_6 _09351_ (.A(_00070_),
    .X(_04086_));
 sky130_fd_sc_hd__buf_6 _09352_ (.A(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__mux4_1 _09353_ (.A0(\cpuregs.regs[4][1] ),
    .A1(\cpuregs.regs[5][1] ),
    .A2(\cpuregs.regs[6][1] ),
    .A3(\cpuregs.regs[7][1] ),
    .S0(_04085_),
    .S1(_04087_),
    .X(_04088_));
 sky130_fd_sc_hd__mux4_1 _09354_ (.A0(\cpuregs.regs[0][1] ),
    .A1(\cpuregs.regs[1][1] ),
    .A2(\cpuregs.regs[2][1] ),
    .A3(\cpuregs.regs[3][1] ),
    .S0(_04085_),
    .S1(_04087_),
    .X(_04089_));
 sky130_fd_sc_hd__mux2_1 _09355_ (.A0(_04088_),
    .A1(_04089_),
    .S(_04078_),
    .X(_04090_));
 sky130_fd_sc_hd__clkbuf_8 _09356_ (.A(_04058_),
    .X(_04091_));
 sky130_fd_sc_hd__mux4_1 _09357_ (.A0(\cpuregs.regs[12][1] ),
    .A1(\cpuregs.regs[13][1] ),
    .A2(\cpuregs.regs[14][1] ),
    .A3(\cpuregs.regs[15][1] ),
    .S0(_04056_),
    .S1(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__mux4_1 _09358_ (.A0(\cpuregs.regs[8][1] ),
    .A1(\cpuregs.regs[9][1] ),
    .A2(\cpuregs.regs[10][1] ),
    .A3(\cpuregs.regs[11][1] ),
    .S0(_04056_),
    .S1(_04091_),
    .X(_04093_));
 sky130_fd_sc_hd__mux2_1 _09359_ (.A0(_04092_),
    .A1(_04093_),
    .S(_04064_),
    .X(_04094_));
 sky130_fd_sc_hd__clkbuf_8 _09360_ (.A(_00073_),
    .X(_04095_));
 sky130_fd_sc_hd__a21o_1 _09361_ (.A1(_04053_),
    .A2(_04094_),
    .B1(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__a21oi_1 _09362_ (.A1(_04070_),
    .A2(_04090_),
    .B1(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__or2_1 _09363_ (.A(\cpuregs.raddr1[1] ),
    .B(\cpuregs.raddr1[0] ),
    .X(_04098_));
 sky130_fd_sc_hd__nor4_4 _09364_ (.A(\cpuregs.raddr1[3] ),
    .B(\cpuregs.raddr1[2] ),
    .C(\cpuregs.raddr1[4] ),
    .D(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__buf_6 _09365_ (.A(net300),
    .X(_04100_));
 sky130_fd_sc_hd__a211o_4 _09366_ (.A1(_04067_),
    .A2(_04083_),
    .B1(_04097_),
    .C1(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__nor2_1 _09367_ (.A(_04051_),
    .B(_04101_),
    .Y(_04102_));
 sky130_fd_sc_hd__a221o_1 _09368_ (.A1(\irq_mask[1] ),
    .A2(_04022_),
    .B1(\timer[1] ),
    .B2(_04024_),
    .C1(_04027_),
    .X(_04103_));
 sky130_fd_sc_hd__buf_4 _09369_ (.A(instr_rdinstrh),
    .X(_04104_));
 sky130_fd_sc_hd__clkbuf_4 _09370_ (.A(instr_rdcycleh),
    .X(_04105_));
 sky130_fd_sc_hd__a22o_1 _09371_ (.A1(\count_instr[33] ),
    .A2(_04104_),
    .B1(_04105_),
    .B2(\count_cycle[33] ),
    .X(_04106_));
 sky130_fd_sc_hd__a211o_1 _09372_ (.A1(\count_instr[1] ),
    .A2(_04012_),
    .B1(_04009_),
    .C1(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__a21o_1 _09373_ (.A1(\count_cycle[1] ),
    .A2(_04014_),
    .B1(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__o211a_1 _09374_ (.A1(_04102_),
    .A2(_04103_),
    .B1(_04108_),
    .C1(_03303_),
    .X(_04109_));
 sky130_fd_sc_hd__mux2_1 _09375_ (.A0(net64),
    .A1(net50),
    .S(_04040_),
    .X(_04110_));
 sky130_fd_sc_hd__and3_1 _09376_ (.A(_04037_),
    .B(_04038_),
    .C(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__a221o_1 _09377_ (.A1(net44),
    .A2(net258),
    .B1(_04035_),
    .B2(net41),
    .C1(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__nand2_1 _09378_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .Y(_04113_));
 sky130_fd_sc_hd__or2_1 _09379_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .X(_04114_));
 sky130_fd_sc_hd__and3b_1 _09380_ (.A_N(_04045_),
    .B(_04113_),
    .C(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__inv_2 _09381_ (.A(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__a21bo_1 _09382_ (.A1(_04113_),
    .A2(_04114_),
    .B1_N(_04045_),
    .X(_04117_));
 sky130_fd_sc_hd__and2_1 _09383_ (.A(_04040_),
    .B(_03312_),
    .X(_04118_));
 sky130_fd_sc_hd__a31o_1 _09384_ (.A1(_03384_),
    .A2(_04116_),
    .A3(_04117_),
    .B1(_04118_),
    .X(_04119_));
 sky130_fd_sc_hd__a211o_1 _09385_ (.A1(_03226_),
    .A2(_04112_),
    .B1(_04119_),
    .C1(_04049_),
    .X(_04120_));
 sky130_fd_sc_hd__o22a_1 _09386_ (.A1(\irq_pending[1] ),
    .A2(_04008_),
    .B1(_04109_),
    .B2(_04120_),
    .X(_08380_));
 sky130_fd_sc_hd__buf_6 _09387_ (.A(_04077_),
    .X(_04121_));
 sky130_fd_sc_hd__mux4_1 _09388_ (.A0(\cpuregs.regs[20][2] ),
    .A1(\cpuregs.regs[21][2] ),
    .A2(\cpuregs.regs[22][2] ),
    .A3(\cpuregs.regs[23][2] ),
    .S0(_04072_),
    .S1(_04074_),
    .X(_04122_));
 sky130_fd_sc_hd__buf_6 _09389_ (.A(_00069_),
    .X(_04123_));
 sky130_fd_sc_hd__clkbuf_8 _09390_ (.A(_00070_),
    .X(_04124_));
 sky130_fd_sc_hd__mux4_1 _09391_ (.A0(\cpuregs.regs[16][2] ),
    .A1(\cpuregs.regs[17][2] ),
    .A2(\cpuregs.regs[18][2] ),
    .A3(\cpuregs.regs[19][2] ),
    .S0(_04123_),
    .S1(_04124_),
    .X(_04125_));
 sky130_fd_sc_hd__or2_1 _09392_ (.A(_00071_),
    .B(_04125_),
    .X(_04126_));
 sky130_fd_sc_hd__o211a_1 _09393_ (.A1(_04121_),
    .A2(_04122_),
    .B1(_04126_),
    .C1(_04068_),
    .X(_04127_));
 sky130_fd_sc_hd__mux4_1 _09394_ (.A0(\cpuregs.regs[24][2] ),
    .A1(\cpuregs.regs[25][2] ),
    .A2(\cpuregs.regs[26][2] ),
    .A3(\cpuregs.regs[27][2] ),
    .S0(_04071_),
    .S1(_04073_),
    .X(_04128_));
 sky130_fd_sc_hd__mux4_1 _09395_ (.A0(\cpuregs.regs[28][2] ),
    .A1(\cpuregs.regs[29][2] ),
    .A2(\cpuregs.regs[30][2] ),
    .A3(\cpuregs.regs[31][2] ),
    .S0(_04071_),
    .S1(_04073_),
    .X(_04129_));
 sky130_fd_sc_hd__mux2_1 _09396_ (.A0(_04128_),
    .A1(_04129_),
    .S(_00071_),
    .X(_04130_));
 sky130_fd_sc_hd__a21o_1 _09397_ (.A1(_04052_),
    .A2(_04130_),
    .B1(_04080_),
    .X(_04131_));
 sky130_fd_sc_hd__or4_1 _09398_ (.A(\cpuregs.raddr1[3] ),
    .B(\cpuregs.raddr1[2] ),
    .C(\cpuregs.raddr1[4] ),
    .D(_04098_),
    .X(_04132_));
 sky130_fd_sc_hd__buf_8 _09399_ (.A(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__mux4_1 _09400_ (.A0(\cpuregs.regs[0][2] ),
    .A1(\cpuregs.regs[1][2] ),
    .A2(\cpuregs.regs[2][2] ),
    .A3(\cpuregs.regs[3][2] ),
    .S0(_04123_),
    .S1(_04124_),
    .X(_04134_));
 sky130_fd_sc_hd__or2_1 _09401_ (.A(_00071_),
    .B(_04134_),
    .X(_04135_));
 sky130_fd_sc_hd__mux4_1 _09402_ (.A0(\cpuregs.regs[4][2] ),
    .A1(\cpuregs.regs[5][2] ),
    .A2(\cpuregs.regs[6][2] ),
    .A3(\cpuregs.regs[7][2] ),
    .S0(_04071_),
    .S1(_04073_),
    .X(_04136_));
 sky130_fd_sc_hd__o21a_1 _09403_ (.A1(_04064_),
    .A2(_04136_),
    .B1(_04068_),
    .X(_04137_));
 sky130_fd_sc_hd__mux4_1 _09404_ (.A0(\cpuregs.regs[12][2] ),
    .A1(\cpuregs.regs[13][2] ),
    .A2(\cpuregs.regs[14][2] ),
    .A3(\cpuregs.regs[15][2] ),
    .S0(_04123_),
    .S1(_04124_),
    .X(_04138_));
 sky130_fd_sc_hd__mux4_1 _09405_ (.A0(\cpuregs.regs[8][2] ),
    .A1(\cpuregs.regs[9][2] ),
    .A2(\cpuregs.regs[10][2] ),
    .A3(\cpuregs.regs[11][2] ),
    .S0(_04123_),
    .S1(_04058_),
    .X(_04139_));
 sky130_fd_sc_hd__mux2_1 _09406_ (.A0(_04138_),
    .A1(_04139_),
    .S(_04077_),
    .X(_04140_));
 sky130_fd_sc_hd__a221o_1 _09407_ (.A1(_04135_),
    .A2(_04137_),
    .B1(_04140_),
    .B2(_04052_),
    .C1(_00073_),
    .X(_04141_));
 sky130_fd_sc_hd__o211ai_4 _09408_ (.A1(_04127_),
    .A2(_04131_),
    .B1(_04133_),
    .C1(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__nor2_1 _09409_ (.A(_04051_),
    .B(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__a221o_1 _09410_ (.A1(\irq_mask[2] ),
    .A2(_04022_),
    .B1(\timer[2] ),
    .B2(_04024_),
    .C1(_04027_),
    .X(_04144_));
 sky130_fd_sc_hd__clkbuf_4 _09411_ (.A(_04011_),
    .X(_04145_));
 sky130_fd_sc_hd__a22o_1 _09412_ (.A1(\count_instr[34] ),
    .A2(_04015_),
    .B1(_04017_),
    .B2(\count_cycle[34] ),
    .X(_04146_));
 sky130_fd_sc_hd__a211o_1 _09413_ (.A1(\count_instr[2] ),
    .A2(_04145_),
    .B1(_04009_),
    .C1(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__a21o_1 _09414_ (.A1(\count_cycle[2] ),
    .A2(_04014_),
    .B1(_04147_),
    .X(_04148_));
 sky130_fd_sc_hd__clkbuf_4 _09415_ (.A(_03301_),
    .X(_04149_));
 sky130_fd_sc_hd__clkbuf_4 _09416_ (.A(_04149_),
    .X(_04150_));
 sky130_fd_sc_hd__o211a_1 _09417_ (.A1(_04143_),
    .A2(_04144_),
    .B1(_04148_),
    .C1(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__nand2_1 _09418_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .Y(_04152_));
 sky130_fd_sc_hd__or2_1 _09419_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .X(_04153_));
 sky130_fd_sc_hd__nor2_1 _09420_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .Y(_04154_));
 sky130_fd_sc_hd__o21ai_2 _09421_ (.A1(_04045_),
    .A2(_04154_),
    .B1(_04113_),
    .Y(_04155_));
 sky130_fd_sc_hd__buf_4 _09422_ (.A(_03317_),
    .X(_04156_));
 sky130_fd_sc_hd__a31o_1 _09423_ (.A1(_04152_),
    .A2(_04153_),
    .A3(_04155_),
    .B1(_04156_),
    .X(_04157_));
 sky130_fd_sc_hd__a21o_1 _09424_ (.A1(_04152_),
    .A2(_04153_),
    .B1(_04155_),
    .X(_04158_));
 sky130_fd_sc_hd__and2b_1 _09425_ (.A_N(_04157_),
    .B(_04158_),
    .X(_04159_));
 sky130_fd_sc_hd__clkbuf_4 _09426_ (.A(net89),
    .X(_04160_));
 sky130_fd_sc_hd__mux2_1 _09427_ (.A0(net34),
    .A1(net51),
    .S(_04039_),
    .X(_04161_));
 sky130_fd_sc_hd__and3_1 _09428_ (.A(_04037_),
    .B(_04038_),
    .C(_04161_),
    .X(_04162_));
 sky130_fd_sc_hd__a221o_1 _09429_ (.A1(net55),
    .A2(net258),
    .B1(_04035_),
    .B2(net42),
    .C1(_04162_),
    .X(_04163_));
 sky130_fd_sc_hd__a221o_1 _09430_ (.A1(_03680_),
    .A2(_04160_),
    .B1(_04163_),
    .B2(_03226_),
    .C1(_04049_),
    .X(_04164_));
 sky130_fd_sc_hd__o32a_2 _09431_ (.A1(_04151_),
    .A2(_04159_),
    .A3(_04164_),
    .B1(_04008_),
    .B2(\irq_pending[2] ),
    .X(_08391_));
 sky130_fd_sc_hd__clkbuf_4 _09432_ (.A(_03253_),
    .X(_04165_));
 sky130_fd_sc_hd__a22o_1 _09433_ (.A1(\count_instr[35] ),
    .A2(_04104_),
    .B1(_04145_),
    .B2(\count_instr[3] ),
    .X(_04166_));
 sky130_fd_sc_hd__a221o_1 _09434_ (.A1(_04018_),
    .A2(\count_cycle[35] ),
    .B1(_04165_),
    .B2(\count_cycle[3] ),
    .C1(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__buf_4 _09435_ (.A(instr_retirq),
    .X(_04168_));
 sky130_fd_sc_hd__mux4_1 _09436_ (.A0(\cpuregs.regs[28][3] ),
    .A1(\cpuregs.regs[29][3] ),
    .A2(\cpuregs.regs[30][3] ),
    .A3(\cpuregs.regs[31][3] ),
    .S0(_04056_),
    .S1(_04091_),
    .X(_04169_));
 sky130_fd_sc_hd__mux4_1 _09437_ (.A0(\cpuregs.regs[24][3] ),
    .A1(\cpuregs.regs[25][3] ),
    .A2(\cpuregs.regs[26][3] ),
    .A3(\cpuregs.regs[27][3] ),
    .S0(_04056_),
    .S1(_04086_),
    .X(_04170_));
 sky130_fd_sc_hd__mux2_1 _09438_ (.A0(_04169_),
    .A1(_04170_),
    .S(_04064_),
    .X(_04171_));
 sky130_fd_sc_hd__nand2_1 _09439_ (.A(_04053_),
    .B(_04171_),
    .Y(_04172_));
 sky130_fd_sc_hd__mux4_1 _09440_ (.A0(\cpuregs.regs[20][3] ),
    .A1(\cpuregs.regs[21][3] ),
    .A2(\cpuregs.regs[22][3] ),
    .A3(\cpuregs.regs[23][3] ),
    .S0(_04071_),
    .S1(_04073_),
    .X(_04173_));
 sky130_fd_sc_hd__mux4_1 _09441_ (.A0(\cpuregs.regs[16][3] ),
    .A1(\cpuregs.regs[17][3] ),
    .A2(\cpuregs.regs[18][3] ),
    .A3(\cpuregs.regs[19][3] ),
    .S0(_04071_),
    .S1(_04073_),
    .X(_04174_));
 sky130_fd_sc_hd__mux2_1 _09442_ (.A0(_04173_),
    .A1(_04174_),
    .S(_04077_),
    .X(_04175_));
 sky130_fd_sc_hd__a21oi_1 _09443_ (.A1(_04069_),
    .A2(_04175_),
    .B1(_04081_),
    .Y(_04176_));
 sky130_fd_sc_hd__mux4_1 _09444_ (.A0(\cpuregs.regs[4][3] ),
    .A1(\cpuregs.regs[5][3] ),
    .A2(\cpuregs.regs[6][3] ),
    .A3(\cpuregs.regs[7][3] ),
    .S0(_04084_),
    .S1(_04086_),
    .X(_04177_));
 sky130_fd_sc_hd__mux4_1 _09445_ (.A0(\cpuregs.regs[0][3] ),
    .A1(\cpuregs.regs[1][3] ),
    .A2(\cpuregs.regs[2][3] ),
    .A3(\cpuregs.regs[3][3] ),
    .S0(_04084_),
    .S1(_04086_),
    .X(_04178_));
 sky130_fd_sc_hd__mux2_1 _09446_ (.A0(_04177_),
    .A1(_04178_),
    .S(_04077_),
    .X(_04179_));
 sky130_fd_sc_hd__mux4_1 _09447_ (.A0(\cpuregs.regs[12][3] ),
    .A1(\cpuregs.regs[13][3] ),
    .A2(\cpuregs.regs[14][3] ),
    .A3(\cpuregs.regs[15][3] ),
    .S0(_04055_),
    .S1(_04058_),
    .X(_04180_));
 sky130_fd_sc_hd__mux4_1 _09448_ (.A0(\cpuregs.regs[8][3] ),
    .A1(\cpuregs.regs[9][3] ),
    .A2(\cpuregs.regs[10][3] ),
    .A3(\cpuregs.regs[11][3] ),
    .S0(_04055_),
    .S1(_04058_),
    .X(_04181_));
 sky130_fd_sc_hd__mux2_1 _09449_ (.A0(_04180_),
    .A1(_04181_),
    .S(_04063_),
    .X(_04182_));
 sky130_fd_sc_hd__a21o_1 _09450_ (.A1(_04052_),
    .A2(_04182_),
    .B1(_00073_),
    .X(_04183_));
 sky130_fd_sc_hd__a21oi_1 _09451_ (.A1(_04069_),
    .A2(_04179_),
    .B1(_04183_),
    .Y(_04184_));
 sky130_fd_sc_hd__a211o_4 _09452_ (.A1(_04172_),
    .A2(_04176_),
    .B1(_04099_),
    .C1(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__inv_2 _09453_ (.A(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hd__clkbuf_4 _09454_ (.A(instr_timer),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_4 _09455_ (.A(_04025_),
    .X(_04188_));
 sky130_fd_sc_hd__a221o_1 _09456_ (.A1(\irq_mask[3] ),
    .A2(_04021_),
    .B1(\timer[3] ),
    .B2(_04187_),
    .C1(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__a21o_1 _09457_ (.A1(_04168_),
    .A2(_04186_),
    .B1(_04189_),
    .X(_04190_));
 sky130_fd_sc_hd__o211a_1 _09458_ (.A1(_04010_),
    .A2(_04167_),
    .B1(_04190_),
    .C1(_04150_),
    .X(_04191_));
 sky130_fd_sc_hd__nand2_1 _09459_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .Y(_04192_));
 sky130_fd_sc_hd__or2_1 _09460_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .X(_04193_));
 sky130_fd_sc_hd__a21bo_1 _09461_ (.A1(_04153_),
    .A2(_04155_),
    .B1_N(_04152_),
    .X(_04194_));
 sky130_fd_sc_hd__a31o_1 _09462_ (.A1(_04192_),
    .A2(_04193_),
    .A3(_04194_),
    .B1(_04156_),
    .X(_04195_));
 sky130_fd_sc_hd__a21o_1 _09463_ (.A1(_04192_),
    .A2(_04193_),
    .B1(_04194_),
    .X(_04196_));
 sky130_fd_sc_hd__and2b_1 _09464_ (.A_N(_04195_),
    .B(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__clkbuf_4 _09465_ (.A(net92),
    .X(_04198_));
 sky130_fd_sc_hd__mux2_1 _09466_ (.A0(net35),
    .A1(net52),
    .S(_04039_),
    .X(_04199_));
 sky130_fd_sc_hd__and3_1 _09467_ (.A(_04036_),
    .B(\mem_wordsize[1] ),
    .C(_04199_),
    .X(_04200_));
 sky130_fd_sc_hd__a221o_1 _09468_ (.A1(net58),
    .A2(net258),
    .B1(_04035_),
    .B2(net43),
    .C1(_04200_),
    .X(_04201_));
 sky130_fd_sc_hd__clkbuf_4 _09469_ (.A(_04048_),
    .X(_04202_));
 sky130_fd_sc_hd__a221o_1 _09470_ (.A1(_03680_),
    .A2(_04198_),
    .B1(_04201_),
    .B2(_03226_),
    .C1(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__o32a_2 _09471_ (.A1(_04191_),
    .A2(_04197_),
    .A3(_04203_),
    .B1(_04008_),
    .B2(\irq_pending[3] ),
    .X(_08394_));
 sky130_fd_sc_hd__a22o_1 _09472_ (.A1(\count_instr[36] ),
    .A2(_04104_),
    .B1(_04145_),
    .B2(\count_instr[4] ),
    .X(_04204_));
 sky130_fd_sc_hd__a221o_1 _09473_ (.A1(_04018_),
    .A2(\count_cycle[36] ),
    .B1(_04165_),
    .B2(\count_cycle[4] ),
    .C1(_04204_),
    .X(_04205_));
 sky130_fd_sc_hd__clkbuf_8 _09474_ (.A(_04053_),
    .X(_04206_));
 sky130_fd_sc_hd__buf_6 _09475_ (.A(_04072_),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_8 _09476_ (.A(_04074_),
    .X(_04208_));
 sky130_fd_sc_hd__mux4_1 _09477_ (.A0(\cpuregs.regs[28][4] ),
    .A1(\cpuregs.regs[29][4] ),
    .A2(\cpuregs.regs[30][4] ),
    .A3(\cpuregs.regs[31][4] ),
    .S0(_04207_),
    .S1(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__mux4_1 _09478_ (.A0(\cpuregs.regs[24][4] ),
    .A1(\cpuregs.regs[25][4] ),
    .A2(\cpuregs.regs[26][4] ),
    .A3(\cpuregs.regs[27][4] ),
    .S0(_04207_),
    .S1(_04208_),
    .X(_04210_));
 sky130_fd_sc_hd__buf_8 _09479_ (.A(_04078_),
    .X(_04211_));
 sky130_fd_sc_hd__mux2_1 _09480_ (.A0(_04209_),
    .A1(_04210_),
    .S(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__nand2_1 _09481_ (.A(_04206_),
    .B(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__clkbuf_8 _09482_ (.A(_04068_),
    .X(_04214_));
 sky130_fd_sc_hd__buf_4 _09483_ (.A(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__buf_6 _09484_ (.A(_04055_),
    .X(_04216_));
 sky130_fd_sc_hd__buf_6 _09485_ (.A(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__buf_4 _09486_ (.A(_04124_),
    .X(_04218_));
 sky130_fd_sc_hd__clkbuf_8 _09487_ (.A(_04218_),
    .X(_04219_));
 sky130_fd_sc_hd__mux4_1 _09488_ (.A0(\cpuregs.regs[20][4] ),
    .A1(\cpuregs.regs[21][4] ),
    .A2(\cpuregs.regs[22][4] ),
    .A3(\cpuregs.regs[23][4] ),
    .S0(_04217_),
    .S1(_04219_),
    .X(_04220_));
 sky130_fd_sc_hd__mux4_1 _09489_ (.A0(\cpuregs.regs[16][4] ),
    .A1(\cpuregs.regs[17][4] ),
    .A2(\cpuregs.regs[18][4] ),
    .A3(\cpuregs.regs[19][4] ),
    .S0(_04217_),
    .S1(_04219_),
    .X(_04221_));
 sky130_fd_sc_hd__buf_6 _09490_ (.A(_04063_),
    .X(_04222_));
 sky130_fd_sc_hd__buf_6 _09491_ (.A(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__mux2_1 _09492_ (.A0(_04220_),
    .A1(_04221_),
    .S(_04223_),
    .X(_04224_));
 sky130_fd_sc_hd__clkbuf_8 _09493_ (.A(_04081_),
    .X(_04225_));
 sky130_fd_sc_hd__a21oi_1 _09494_ (.A1(_04215_),
    .A2(_04224_),
    .B1(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__buf_8 _09495_ (.A(net301),
    .X(_04227_));
 sky130_fd_sc_hd__mux4_1 _09496_ (.A0(\cpuregs.regs[4][4] ),
    .A1(\cpuregs.regs[5][4] ),
    .A2(\cpuregs.regs[6][4] ),
    .A3(\cpuregs.regs[7][4] ),
    .S0(_04207_),
    .S1(_04208_),
    .X(_04228_));
 sky130_fd_sc_hd__mux4_1 _09497_ (.A0(\cpuregs.regs[0][4] ),
    .A1(\cpuregs.regs[1][4] ),
    .A2(\cpuregs.regs[2][4] ),
    .A3(\cpuregs.regs[3][4] ),
    .S0(_04207_),
    .S1(_04208_),
    .X(_04229_));
 sky130_fd_sc_hd__mux2_1 _09498_ (.A0(_04228_),
    .A1(_04229_),
    .S(_04211_),
    .X(_04230_));
 sky130_fd_sc_hd__buf_6 _09499_ (.A(_04052_),
    .X(_04231_));
 sky130_fd_sc_hd__buf_6 _09500_ (.A(_04084_),
    .X(_04232_));
 sky130_fd_sc_hd__clkbuf_8 _09501_ (.A(_04091_),
    .X(_04233_));
 sky130_fd_sc_hd__mux4_1 _09502_ (.A0(\cpuregs.regs[12][4] ),
    .A1(\cpuregs.regs[13][4] ),
    .A2(\cpuregs.regs[14][4] ),
    .A3(\cpuregs.regs[15][4] ),
    .S0(_04232_),
    .S1(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__mux4_1 _09503_ (.A0(\cpuregs.regs[8][4] ),
    .A1(\cpuregs.regs[9][4] ),
    .A2(\cpuregs.regs[10][4] ),
    .A3(\cpuregs.regs[11][4] ),
    .S0(_04232_),
    .S1(_04233_),
    .X(_04235_));
 sky130_fd_sc_hd__mux2_1 _09504_ (.A0(_04234_),
    .A1(_04235_),
    .S(_04121_),
    .X(_04236_));
 sky130_fd_sc_hd__buf_6 _09505_ (.A(_00073_),
    .X(_04237_));
 sky130_fd_sc_hd__a21o_1 _09506_ (.A1(_04231_),
    .A2(_04236_),
    .B1(_04237_),
    .X(_04238_));
 sky130_fd_sc_hd__a21oi_1 _09507_ (.A1(_04215_),
    .A2(_04230_),
    .B1(_04238_),
    .Y(_04239_));
 sky130_fd_sc_hd__a211o_4 _09508_ (.A1(_04213_),
    .A2(_04226_),
    .B1(_04227_),
    .C1(_04239_),
    .X(_04240_));
 sky130_fd_sc_hd__inv_2 _09509_ (.A(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__a221o_1 _09510_ (.A1(\irq_mask[4] ),
    .A2(_04021_),
    .B1(\timer[4] ),
    .B2(_04187_),
    .C1(_04188_),
    .X(_04242_));
 sky130_fd_sc_hd__a21o_1 _09511_ (.A1(_04168_),
    .A2(_04241_),
    .B1(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__o211a_1 _09512_ (.A1(_04010_),
    .A2(_04205_),
    .B1(_04243_),
    .C1(_04150_),
    .X(_04244_));
 sky130_fd_sc_hd__nand2_1 _09513_ (.A(\reg_pc[4] ),
    .B(\decoded_imm[4] ),
    .Y(_04245_));
 sky130_fd_sc_hd__or2_1 _09514_ (.A(\reg_pc[4] ),
    .B(\decoded_imm[4] ),
    .X(_04246_));
 sky130_fd_sc_hd__a21bo_1 _09515_ (.A1(_04193_),
    .A2(_04194_),
    .B1_N(_04192_),
    .X(_04247_));
 sky130_fd_sc_hd__and3_1 _09516_ (.A(_04245_),
    .B(_04246_),
    .C(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__a21o_1 _09517_ (.A1(_04245_),
    .A2(_04246_),
    .B1(_04247_),
    .X(_04249_));
 sky130_fd_sc_hd__and3b_1 _09518_ (.A_N(_04248_),
    .B(_04249_),
    .C(_03384_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_4 _09519_ (.A(net93),
    .X(_04251_));
 sky130_fd_sc_hd__mux2_1 _09520_ (.A0(net36),
    .A1(net53),
    .S(_04039_),
    .X(_04252_));
 sky130_fd_sc_hd__and3_1 _09521_ (.A(_04036_),
    .B(\mem_wordsize[1] ),
    .C(_04252_),
    .X(_04253_));
 sky130_fd_sc_hd__a221o_1 _09522_ (.A1(net59),
    .A2(net258),
    .B1(_04035_),
    .B2(net45),
    .C1(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__a221o_2 _09523_ (.A1(_03680_),
    .A2(_04251_),
    .B1(_04254_),
    .B2(_03226_),
    .C1(_04202_),
    .X(_04255_));
 sky130_fd_sc_hd__o32a_2 _09524_ (.A1(_04244_),
    .A2(_04250_),
    .A3(_04255_),
    .B1(_04008_),
    .B2(\irq_pending[4] ),
    .X(_08395_));
 sky130_fd_sc_hd__inv_2 _09525_ (.A(_04245_),
    .Y(_04256_));
 sky130_fd_sc_hd__nor2_1 _09526_ (.A(_04256_),
    .B(_04248_),
    .Y(_04257_));
 sky130_fd_sc_hd__nor2_1 _09527_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .Y(_04258_));
 sky130_fd_sc_hd__and2_1 _09528_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .X(_04259_));
 sky130_fd_sc_hd__nor2_1 _09529_ (.A(_04258_),
    .B(_04259_),
    .Y(_04260_));
 sky130_fd_sc_hd__xnor2_1 _09530_ (.A(_04257_),
    .B(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__clkbuf_4 _09531_ (.A(_03524_),
    .X(_04262_));
 sky130_fd_sc_hd__mux2_1 _09532_ (.A0(net37),
    .A1(net54),
    .S(_04039_),
    .X(_04263_));
 sky130_fd_sc_hd__and3_1 _09533_ (.A(_04036_),
    .B(\mem_wordsize[1] ),
    .C(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__a221o_2 _09534_ (.A1(net60),
    .A2(net258),
    .B1(_04035_),
    .B2(net46),
    .C1(_04264_),
    .X(_04265_));
 sky130_fd_sc_hd__buf_2 _09535_ (.A(_04048_),
    .X(_04266_));
 sky130_fd_sc_hd__a221o_1 _09536_ (.A1(_03637_),
    .A2(_04262_),
    .B1(_04265_),
    .B2(_03225_),
    .C1(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_4 _09537_ (.A(_04009_),
    .X(_04268_));
 sky130_fd_sc_hd__a22o_1 _09538_ (.A1(\count_instr[5] ),
    .A2(_04011_),
    .B1(_04017_),
    .B2(\count_cycle[37] ),
    .X(_04269_));
 sky130_fd_sc_hd__a221o_1 _09539_ (.A1(\count_instr[37] ),
    .A2(_04016_),
    .B1(\count_cycle[5] ),
    .B2(_04013_),
    .C1(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__buf_4 _09540_ (.A(instr_retirq),
    .X(_04271_));
 sky130_fd_sc_hd__clkbuf_8 _09541_ (.A(_04054_),
    .X(_04272_));
 sky130_fd_sc_hd__buf_8 _09542_ (.A(_04055_),
    .X(_04273_));
 sky130_fd_sc_hd__clkbuf_8 _09543_ (.A(_04273_),
    .X(_04274_));
 sky130_fd_sc_hd__clkbuf_8 _09544_ (.A(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__buf_4 _09545_ (.A(_04058_),
    .X(_04276_));
 sky130_fd_sc_hd__buf_4 _09546_ (.A(_04276_),
    .X(_04277_));
 sky130_fd_sc_hd__buf_4 _09547_ (.A(_04277_),
    .X(_04278_));
 sky130_fd_sc_hd__mux4_1 _09548_ (.A0(\cpuregs.regs[12][5] ),
    .A1(\cpuregs.regs[13][5] ),
    .A2(\cpuregs.regs[14][5] ),
    .A3(\cpuregs.regs[15][5] ),
    .S0(_04275_),
    .S1(_04278_),
    .X(_04279_));
 sky130_fd_sc_hd__buf_6 _09549_ (.A(_04055_),
    .X(_04280_));
 sky130_fd_sc_hd__buf_6 _09550_ (.A(_04280_),
    .X(_04281_));
 sky130_fd_sc_hd__buf_6 _09551_ (.A(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__clkbuf_8 _09552_ (.A(_04058_),
    .X(_04283_));
 sky130_fd_sc_hd__buf_6 _09553_ (.A(_04283_),
    .X(_04284_));
 sky130_fd_sc_hd__clkbuf_8 _09554_ (.A(_04284_),
    .X(_04285_));
 sky130_fd_sc_hd__mux4_1 _09555_ (.A0(\cpuregs.regs[8][5] ),
    .A1(\cpuregs.regs[9][5] ),
    .A2(\cpuregs.regs[10][5] ),
    .A3(\cpuregs.regs[11][5] ),
    .S0(_04282_),
    .S1(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__clkbuf_8 _09556_ (.A(_04065_),
    .X(_04287_));
 sky130_fd_sc_hd__mux2_1 _09557_ (.A0(_04279_),
    .A1(_04286_),
    .S(_04287_),
    .X(_04288_));
 sky130_fd_sc_hd__clkbuf_8 _09558_ (.A(_04214_),
    .X(_04289_));
 sky130_fd_sc_hd__buf_6 _09559_ (.A(_04055_),
    .X(_04290_));
 sky130_fd_sc_hd__clkbuf_8 _09560_ (.A(_04290_),
    .X(_04291_));
 sky130_fd_sc_hd__buf_4 _09561_ (.A(_04276_),
    .X(_04292_));
 sky130_fd_sc_hd__mux4_1 _09562_ (.A0(\cpuregs.regs[4][5] ),
    .A1(\cpuregs.regs[5][5] ),
    .A2(\cpuregs.regs[6][5] ),
    .A3(\cpuregs.regs[7][5] ),
    .S0(_04291_),
    .S1(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__mux4_1 _09563_ (.A0(\cpuregs.regs[0][5] ),
    .A1(\cpuregs.regs[1][5] ),
    .A2(\cpuregs.regs[2][5] ),
    .A3(\cpuregs.regs[3][5] ),
    .S0(_04291_),
    .S1(_04292_),
    .X(_04294_));
 sky130_fd_sc_hd__mux2_1 _09564_ (.A0(_04293_),
    .A1(_04294_),
    .S(_04223_),
    .X(_04295_));
 sky130_fd_sc_hd__buf_6 _09565_ (.A(_04237_),
    .X(_04296_));
 sky130_fd_sc_hd__a21o_1 _09566_ (.A1(_04289_),
    .A2(_04295_),
    .B1(_04296_),
    .X(_04297_));
 sky130_fd_sc_hd__a21oi_2 _09567_ (.A1(_04272_),
    .A2(_04288_),
    .B1(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__mux4_1 _09568_ (.A0(\cpuregs.regs[28][5] ),
    .A1(\cpuregs.regs[29][5] ),
    .A2(\cpuregs.regs[30][5] ),
    .A3(\cpuregs.regs[31][5] ),
    .S0(_04275_),
    .S1(_04278_),
    .X(_04299_));
 sky130_fd_sc_hd__mux4_1 _09569_ (.A0(\cpuregs.regs[24][5] ),
    .A1(\cpuregs.regs[25][5] ),
    .A2(\cpuregs.regs[26][5] ),
    .A3(\cpuregs.regs[27][5] ),
    .S0(_04275_),
    .S1(_04278_),
    .X(_04300_));
 sky130_fd_sc_hd__mux2_1 _09570_ (.A0(_04299_),
    .A1(_04300_),
    .S(_04287_),
    .X(_04301_));
 sky130_fd_sc_hd__mux4_1 _09571_ (.A0(\cpuregs.regs[20][5] ),
    .A1(\cpuregs.regs[21][5] ),
    .A2(\cpuregs.regs[22][5] ),
    .A3(\cpuregs.regs[23][5] ),
    .S0(_04217_),
    .S1(_04219_),
    .X(_04302_));
 sky130_fd_sc_hd__mux4_1 _09572_ (.A0(\cpuregs.regs[16][5] ),
    .A1(\cpuregs.regs[17][5] ),
    .A2(\cpuregs.regs[18][5] ),
    .A3(\cpuregs.regs[19][5] ),
    .S0(_04217_),
    .S1(_04219_),
    .X(_04303_));
 sky130_fd_sc_hd__mux2_1 _09573_ (.A0(_04302_),
    .A1(_04303_),
    .S(_04223_),
    .X(_04304_));
 sky130_fd_sc_hd__a21o_1 _09574_ (.A1(_04289_),
    .A2(_04304_),
    .B1(_04225_),
    .X(_04305_));
 sky130_fd_sc_hd__a21oi_2 _09575_ (.A1(_04272_),
    .A2(_04301_),
    .B1(_04305_),
    .Y(_04306_));
 sky130_fd_sc_hd__nor3_4 _09576_ (.A(_04227_),
    .B(_04298_),
    .C(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__clkbuf_4 _09577_ (.A(instr_maskirq),
    .X(_04308_));
 sky130_fd_sc_hd__a221o_1 _09578_ (.A1(\irq_mask[5] ),
    .A2(_04308_),
    .B1(\timer[5] ),
    .B2(_04023_),
    .C1(_04026_),
    .X(_04309_));
 sky130_fd_sc_hd__a21o_1 _09579_ (.A1(_04271_),
    .A2(_04307_),
    .B1(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__o211a_1 _09580_ (.A1(_04268_),
    .A2(_04270_),
    .B1(_04310_),
    .C1(_03302_),
    .X(_04311_));
 sky130_fd_sc_hd__a211o_1 _09581_ (.A1(_03385_),
    .A2(_04261_),
    .B1(_04267_),
    .C1(_04311_),
    .X(_04312_));
 sky130_fd_sc_hd__o21a_1 _09582_ (.A1(\irq_pending[5] ),
    .A2(_04008_),
    .B1(_04312_),
    .X(_08396_));
 sky130_fd_sc_hd__mux4_1 _09583_ (.A0(\cpuregs.regs[20][6] ),
    .A1(\cpuregs.regs[21][6] ),
    .A2(\cpuregs.regs[22][6] ),
    .A3(\cpuregs.regs[23][6] ),
    .S0(_04217_),
    .S1(_04219_),
    .X(_04313_));
 sky130_fd_sc_hd__mux4_1 _09584_ (.A0(\cpuregs.regs[16][6] ),
    .A1(\cpuregs.regs[17][6] ),
    .A2(\cpuregs.regs[18][6] ),
    .A3(\cpuregs.regs[19][6] ),
    .S0(_04217_),
    .S1(_04219_),
    .X(_04314_));
 sky130_fd_sc_hd__mux2_1 _09585_ (.A0(_04313_),
    .A1(_04314_),
    .S(_04223_),
    .X(_04315_));
 sky130_fd_sc_hd__nand2_1 _09586_ (.A(_04215_),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__buf_4 _09587_ (.A(_04283_),
    .X(_04317_));
 sky130_fd_sc_hd__mux4_1 _09588_ (.A0(\cpuregs.regs[28][6] ),
    .A1(\cpuregs.regs[29][6] ),
    .A2(\cpuregs.regs[30][6] ),
    .A3(\cpuregs.regs[31][6] ),
    .S0(_04274_),
    .S1(_04317_),
    .X(_04318_));
 sky130_fd_sc_hd__mux4_1 _09589_ (.A0(\cpuregs.regs[24][6] ),
    .A1(\cpuregs.regs[25][6] ),
    .A2(\cpuregs.regs[26][6] ),
    .A3(\cpuregs.regs[27][6] ),
    .S0(_04274_),
    .S1(_04317_),
    .X(_04319_));
 sky130_fd_sc_hd__buf_6 _09590_ (.A(_04063_),
    .X(_04320_));
 sky130_fd_sc_hd__clkbuf_8 _09591_ (.A(_04320_),
    .X(_04321_));
 sky130_fd_sc_hd__mux2_1 _09592_ (.A0(_04318_),
    .A1(_04319_),
    .S(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__a21oi_1 _09593_ (.A1(_04206_),
    .A2(_04322_),
    .B1(_04225_),
    .Y(_04323_));
 sky130_fd_sc_hd__mux4_1 _09594_ (.A0(\cpuregs.regs[4][6] ),
    .A1(\cpuregs.regs[5][6] ),
    .A2(\cpuregs.regs[6][6] ),
    .A3(\cpuregs.regs[7][6] ),
    .S0(_04291_),
    .S1(_04292_),
    .X(_04324_));
 sky130_fd_sc_hd__clkbuf_8 _09595_ (.A(_04273_),
    .X(_04325_));
 sky130_fd_sc_hd__mux4_1 _09596_ (.A0(\cpuregs.regs[0][6] ),
    .A1(\cpuregs.regs[1][6] ),
    .A2(\cpuregs.regs[2][6] ),
    .A3(\cpuregs.regs[3][6] ),
    .S0(_04325_),
    .S1(_04277_),
    .X(_04326_));
 sky130_fd_sc_hd__mux2_1 _09597_ (.A0(_04324_),
    .A1(_04326_),
    .S(_04223_),
    .X(_04327_));
 sky130_fd_sc_hd__buf_4 _09598_ (.A(_04052_),
    .X(_04328_));
 sky130_fd_sc_hd__clkbuf_8 _09599_ (.A(_04123_),
    .X(_04329_));
 sky130_fd_sc_hd__mux4_1 _09600_ (.A0(\cpuregs.regs[12][6] ),
    .A1(\cpuregs.regs[13][6] ),
    .A2(\cpuregs.regs[14][6] ),
    .A3(\cpuregs.regs[15][6] ),
    .S0(_04329_),
    .S1(_04218_),
    .X(_04330_));
 sky130_fd_sc_hd__mux4_1 _09601_ (.A0(\cpuregs.regs[8][6] ),
    .A1(\cpuregs.regs[9][6] ),
    .A2(\cpuregs.regs[10][6] ),
    .A3(\cpuregs.regs[11][6] ),
    .S0(_04329_),
    .S1(_04218_),
    .X(_04331_));
 sky130_fd_sc_hd__mux2_1 _09602_ (.A0(_04330_),
    .A1(_04331_),
    .S(_04222_),
    .X(_04332_));
 sky130_fd_sc_hd__a21o_1 _09603_ (.A1(_04328_),
    .A2(_04332_),
    .B1(_04237_),
    .X(_04333_));
 sky130_fd_sc_hd__a21oi_1 _09604_ (.A1(_04289_),
    .A2(_04327_),
    .B1(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__a211o_4 _09605_ (.A1(_04316_),
    .A2(_04323_),
    .B1(_04100_),
    .C1(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__nor2_1 _09606_ (.A(_04051_),
    .B(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__a221o_1 _09607_ (.A1(\irq_mask[6] ),
    .A2(_04021_),
    .B1(\timer[6] ),
    .B2(_04187_),
    .C1(_04188_),
    .X(_04337_));
 sky130_fd_sc_hd__a22o_1 _09608_ (.A1(\count_instr[38] ),
    .A2(_04015_),
    .B1(instr_rdinstr),
    .B2(\count_instr[6] ),
    .X(_04338_));
 sky130_fd_sc_hd__a211o_1 _09609_ (.A1(_04105_),
    .A2(\count_cycle[38] ),
    .B1(_04009_),
    .C1(_04338_),
    .X(_04339_));
 sky130_fd_sc_hd__a21o_1 _09610_ (.A1(\count_cycle[6] ),
    .A2(_04165_),
    .B1(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__o211a_1 _09611_ (.A1(_04336_),
    .A2(_04337_),
    .B1(_04340_),
    .C1(_04149_),
    .X(_04341_));
 sky130_fd_sc_hd__clkbuf_4 _09612_ (.A(net95),
    .X(_04342_));
 sky130_fd_sc_hd__mux2_1 _09613_ (.A0(net38),
    .A1(net56),
    .S(_04039_),
    .X(_04343_));
 sky130_fd_sc_hd__and3_1 _09614_ (.A(_04036_),
    .B(\mem_wordsize[1] ),
    .C(_04343_),
    .X(_04344_));
 sky130_fd_sc_hd__a221o_2 _09615_ (.A1(net61),
    .A2(net258),
    .B1(_04035_),
    .B2(net47),
    .C1(_04344_),
    .X(_04345_));
 sky130_fd_sc_hd__a22o_1 _09616_ (.A1(_04046_),
    .A2(_04342_),
    .B1(_04345_),
    .B2(_03225_),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_1 _09617_ (.A(\reg_pc[6] ),
    .B(\decoded_imm[6] ),
    .Y(_04347_));
 sky130_fd_sc_hd__or2_1 _09618_ (.A(\reg_pc[6] ),
    .B(\decoded_imm[6] ),
    .X(_04348_));
 sky130_fd_sc_hd__nand2_1 _09619_ (.A(_04347_),
    .B(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__a211o_1 _09620_ (.A1(_04246_),
    .A2(_04247_),
    .B1(_04259_),
    .C1(_04256_),
    .X(_04350_));
 sky130_fd_sc_hd__or3b_2 _09621_ (.A(_04258_),
    .B(_04349_),
    .C_N(_04350_),
    .X(_04351_));
 sky130_fd_sc_hd__or2_1 _09622_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .X(_04352_));
 sky130_fd_sc_hd__a21bo_1 _09623_ (.A1(_04352_),
    .A2(_04350_),
    .B1_N(_04349_),
    .X(_04353_));
 sky130_fd_sc_hd__a32o_1 _09624_ (.A1(\cpu_state[3] ),
    .A2(_04351_),
    .A3(_04353_),
    .B1(\irq_pending[6] ),
    .B2(_04266_),
    .X(_04354_));
 sky130_fd_sc_hd__or3_1 _09625_ (.A(_04341_),
    .B(_04346_),
    .C(_04354_),
    .X(_04355_));
 sky130_fd_sc_hd__clkbuf_1 _09626_ (.A(_04355_),
    .X(_08397_));
 sky130_fd_sc_hd__and2_1 _09627_ (.A(\reg_pc[7] ),
    .B(\decoded_imm[7] ),
    .X(_04356_));
 sky130_fd_sc_hd__nor2_1 _09628_ (.A(\reg_pc[7] ),
    .B(\decoded_imm[7] ),
    .Y(_04357_));
 sky130_fd_sc_hd__o211a_1 _09629_ (.A1(_04356_),
    .A2(_04357_),
    .B1(_04347_),
    .C1(_04351_),
    .X(_04358_));
 sky130_fd_sc_hd__a211oi_2 _09630_ (.A1(_04347_),
    .A2(_04351_),
    .B1(_04356_),
    .C1(_04357_),
    .Y(_04359_));
 sky130_fd_sc_hd__clkbuf_4 _09631_ (.A(_03518_),
    .X(_04360_));
 sky130_fd_sc_hd__or2b_1 _09632_ (.A(net57),
    .B_N(_03242_),
    .X(_04361_));
 sky130_fd_sc_hd__o2111a_1 _09633_ (.A1(_03242_),
    .A2(net39),
    .B1(_04361_),
    .C1(net67),
    .D1(\mem_wordsize[1] ),
    .X(_04362_));
 sky130_fd_sc_hd__a221o_2 _09634_ (.A1(net62),
    .A2(net258),
    .B1(_04035_),
    .B2(net48),
    .C1(_04362_),
    .X(_04363_));
 sky130_fd_sc_hd__mux4_1 _09635_ (.A0(\cpuregs.regs[4][7] ),
    .A1(\cpuregs.regs[5][7] ),
    .A2(\cpuregs.regs[6][7] ),
    .A3(\cpuregs.regs[7][7] ),
    .S0(_04274_),
    .S1(_04317_),
    .X(_04364_));
 sky130_fd_sc_hd__mux4_1 _09636_ (.A0(\cpuregs.regs[0][7] ),
    .A1(\cpuregs.regs[1][7] ),
    .A2(\cpuregs.regs[2][7] ),
    .A3(\cpuregs.regs[3][7] ),
    .S0(_04274_),
    .S1(_04317_),
    .X(_04365_));
 sky130_fd_sc_hd__mux2_1 _09637_ (.A0(_04364_),
    .A1(_04365_),
    .S(_04321_),
    .X(_04366_));
 sky130_fd_sc_hd__mux4_1 _09638_ (.A0(\cpuregs.regs[8][7] ),
    .A1(\cpuregs.regs[9][7] ),
    .A2(\cpuregs.regs[10][7] ),
    .A3(\cpuregs.regs[11][7] ),
    .S0(_04290_),
    .S1(_04276_),
    .X(_04367_));
 sky130_fd_sc_hd__mux4_1 _09639_ (.A0(\cpuregs.regs[12][7] ),
    .A1(\cpuregs.regs[13][7] ),
    .A2(\cpuregs.regs[14][7] ),
    .A3(\cpuregs.regs[15][7] ),
    .S0(_04290_),
    .S1(_04276_),
    .X(_04368_));
 sky130_fd_sc_hd__buf_6 _09640_ (.A(_00071_),
    .X(_04369_));
 sky130_fd_sc_hd__mux2_1 _09641_ (.A0(_04367_),
    .A1(_04368_),
    .S(_04369_),
    .X(_04370_));
 sky130_fd_sc_hd__a21o_1 _09642_ (.A1(_04328_),
    .A2(_04370_),
    .B1(_04237_),
    .X(_04371_));
 sky130_fd_sc_hd__a21oi_1 _09643_ (.A1(_04289_),
    .A2(_04366_),
    .B1(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__mux4_1 _09644_ (.A0(\cpuregs.regs[28][7] ),
    .A1(\cpuregs.regs[29][7] ),
    .A2(\cpuregs.regs[30][7] ),
    .A3(\cpuregs.regs[31][7] ),
    .S0(_04325_),
    .S1(_04277_),
    .X(_04373_));
 sky130_fd_sc_hd__mux4_1 _09645_ (.A0(\cpuregs.regs[24][7] ),
    .A1(\cpuregs.regs[25][7] ),
    .A2(\cpuregs.regs[26][7] ),
    .A3(\cpuregs.regs[27][7] ),
    .S0(_04325_),
    .S1(_04317_),
    .X(_04374_));
 sky130_fd_sc_hd__mux2_1 _09646_ (.A0(_04373_),
    .A1(_04374_),
    .S(_04321_),
    .X(_04375_));
 sky130_fd_sc_hd__clkbuf_8 _09647_ (.A(_04124_),
    .X(_04376_));
 sky130_fd_sc_hd__mux4_1 _09648_ (.A0(\cpuregs.regs[20][7] ),
    .A1(\cpuregs.regs[21][7] ),
    .A2(\cpuregs.regs[22][7] ),
    .A3(\cpuregs.regs[23][7] ),
    .S0(_04216_),
    .S1(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__mux4_1 _09649_ (.A0(\cpuregs.regs[16][7] ),
    .A1(\cpuregs.regs[17][7] ),
    .A2(\cpuregs.regs[18][7] ),
    .A3(\cpuregs.regs[19][7] ),
    .S0(_04216_),
    .S1(_04376_),
    .X(_04378_));
 sky130_fd_sc_hd__mux2_1 _09650_ (.A0(_04377_),
    .A1(_04378_),
    .S(_04222_),
    .X(_04379_));
 sky130_fd_sc_hd__a21o_1 _09651_ (.A1(_04214_),
    .A2(_04379_),
    .B1(_04081_),
    .X(_04380_));
 sky130_fd_sc_hd__a21oi_1 _09652_ (.A1(_04206_),
    .A2(_04375_),
    .B1(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__or3_4 _09653_ (.A(_04100_),
    .B(_04372_),
    .C(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__nor2_1 _09654_ (.A(_04051_),
    .B(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__a221o_1 _09655_ (.A1(\irq_mask[7] ),
    .A2(_04308_),
    .B1(\timer[7] ),
    .B2(_04023_),
    .C1(_04026_),
    .X(_04384_));
 sky130_fd_sc_hd__a22o_1 _09656_ (.A1(\count_instr[39] ),
    .A2(instr_rdinstrh),
    .B1(instr_rdinstr),
    .B2(\count_instr[7] ),
    .X(_04385_));
 sky130_fd_sc_hd__a211o_1 _09657_ (.A1(instr_rdcycleh),
    .A2(\count_cycle[39] ),
    .B1(_03252_),
    .C1(_04385_),
    .X(_04386_));
 sky130_fd_sc_hd__a21o_1 _09658_ (.A1(\count_cycle[7] ),
    .A2(_04013_),
    .B1(_04386_),
    .X(_04387_));
 sky130_fd_sc_hd__o211a_2 _09659_ (.A1(_04383_),
    .A2(_04384_),
    .B1(_04387_),
    .C1(_03301_),
    .X(_04388_));
 sky130_fd_sc_hd__a221o_2 _09660_ (.A1(_03680_),
    .A2(_04360_),
    .B1(_04363_),
    .B2(_03225_),
    .C1(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__a21oi_2 _09661_ (.A1(\irq_pending[7] ),
    .A2(_04049_),
    .B1(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__o31ai_1 _09662_ (.A1(_04156_),
    .A2(_04358_),
    .A3(_04359_),
    .B1(_04390_),
    .Y(_08398_));
 sky130_fd_sc_hd__clkbuf_4 _09663_ (.A(_03385_),
    .X(_04391_));
 sky130_fd_sc_hd__nand2_1 _09664_ (.A(\reg_pc[8] ),
    .B(\decoded_imm[8] ),
    .Y(_04392_));
 sky130_fd_sc_hd__or2_1 _09665_ (.A(\reg_pc[8] ),
    .B(\decoded_imm[8] ),
    .X(_04393_));
 sky130_fd_sc_hd__a211o_1 _09666_ (.A1(_04392_),
    .A2(_04393_),
    .B1(_04356_),
    .C1(_04359_),
    .X(_04394_));
 sky130_fd_sc_hd__o211ai_2 _09667_ (.A1(_04356_),
    .A2(_04359_),
    .B1(_04392_),
    .C1(_04393_),
    .Y(_04395_));
 sky130_fd_sc_hd__a22o_1 _09668_ (.A1(\count_instr[40] ),
    .A2(_04104_),
    .B1(_04011_),
    .B2(\count_instr[8] ),
    .X(_04396_));
 sky130_fd_sc_hd__a221o_1 _09669_ (.A1(_04105_),
    .A2(\count_cycle[40] ),
    .B1(_04013_),
    .B2(\count_cycle[8] ),
    .C1(_04396_),
    .X(_04397_));
 sky130_fd_sc_hd__mux4_1 _09670_ (.A0(\cpuregs.regs[4][8] ),
    .A1(\cpuregs.regs[5][8] ),
    .A2(\cpuregs.regs[6][8] ),
    .A3(\cpuregs.regs[7][8] ),
    .S0(_04072_),
    .S1(_04074_),
    .X(_04398_));
 sky130_fd_sc_hd__mux4_1 _09671_ (.A0(\cpuregs.regs[0][8] ),
    .A1(\cpuregs.regs[1][8] ),
    .A2(\cpuregs.regs[2][8] ),
    .A3(\cpuregs.regs[3][8] ),
    .S0(_04072_),
    .S1(_04074_),
    .X(_04399_));
 sky130_fd_sc_hd__mux2_1 _09672_ (.A0(_04398_),
    .A1(_04399_),
    .S(_04078_),
    .X(_04400_));
 sky130_fd_sc_hd__mux4_1 _09673_ (.A0(\cpuregs.regs[8][8] ),
    .A1(\cpuregs.regs[9][8] ),
    .A2(\cpuregs.regs[10][8] ),
    .A3(\cpuregs.regs[11][8] ),
    .S0(_04056_),
    .S1(_04091_),
    .X(_04401_));
 sky130_fd_sc_hd__mux4_1 _09674_ (.A0(\cpuregs.regs[12][8] ),
    .A1(\cpuregs.regs[13][8] ),
    .A2(\cpuregs.regs[14][8] ),
    .A3(\cpuregs.regs[15][8] ),
    .S0(_04056_),
    .S1(_04091_),
    .X(_04402_));
 sky130_fd_sc_hd__mux2_1 _09675_ (.A0(_04401_),
    .A1(_04402_),
    .S(_00071_),
    .X(_04403_));
 sky130_fd_sc_hd__a21o_1 _09676_ (.A1(_04053_),
    .A2(_04403_),
    .B1(_04095_),
    .X(_04404_));
 sky130_fd_sc_hd__a21oi_1 _09677_ (.A1(_04070_),
    .A2(_04400_),
    .B1(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__mux4_1 _09678_ (.A0(\cpuregs.regs[28][8] ),
    .A1(\cpuregs.regs[29][8] ),
    .A2(\cpuregs.regs[30][8] ),
    .A3(\cpuregs.regs[31][8] ),
    .S0(_04085_),
    .S1(_04087_),
    .X(_04406_));
 sky130_fd_sc_hd__mux4_1 _09679_ (.A0(\cpuregs.regs[24][8] ),
    .A1(\cpuregs.regs[25][8] ),
    .A2(\cpuregs.regs[26][8] ),
    .A3(\cpuregs.regs[27][8] ),
    .S0(_04085_),
    .S1(_04087_),
    .X(_04407_));
 sky130_fd_sc_hd__mux2_1 _09680_ (.A0(_04406_),
    .A1(_04407_),
    .S(_04078_),
    .X(_04408_));
 sky130_fd_sc_hd__mux4_1 _09681_ (.A0(\cpuregs.regs[20][8] ),
    .A1(\cpuregs.regs[21][8] ),
    .A2(\cpuregs.regs[22][8] ),
    .A3(\cpuregs.regs[23][8] ),
    .S0(_04056_),
    .S1(_04091_),
    .X(_04409_));
 sky130_fd_sc_hd__mux4_1 _09682_ (.A0(\cpuregs.regs[16][8] ),
    .A1(\cpuregs.regs[17][8] ),
    .A2(\cpuregs.regs[18][8] ),
    .A3(\cpuregs.regs[19][8] ),
    .S0(_04056_),
    .S1(_04091_),
    .X(_04410_));
 sky130_fd_sc_hd__mux2_1 _09683_ (.A0(_04409_),
    .A1(_04410_),
    .S(_04064_),
    .X(_04411_));
 sky130_fd_sc_hd__a21o_1 _09684_ (.A1(_04069_),
    .A2(_04411_),
    .B1(_04081_),
    .X(_04412_));
 sky130_fd_sc_hd__a21oi_1 _09685_ (.A1(_04231_),
    .A2(_04408_),
    .B1(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__or3_4 _09686_ (.A(_04099_),
    .B(_04405_),
    .C(_04413_),
    .X(_04414_));
 sky130_fd_sc_hd__inv_2 _09687_ (.A(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hd__a221o_1 _09688_ (.A1(\irq_mask[8] ),
    .A2(_04308_),
    .B1(\timer[8] ),
    .B2(_04023_),
    .C1(_04026_),
    .X(_04416_));
 sky130_fd_sc_hd__a21o_1 _09689_ (.A1(_04271_),
    .A2(_04415_),
    .B1(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__o211a_1 _09690_ (.A1(_04268_),
    .A2(_04397_),
    .B1(_04417_),
    .C1(_04149_),
    .X(_04418_));
 sky130_fd_sc_hd__buf_4 _09691_ (.A(_03510_),
    .X(_04419_));
 sky130_fd_sc_hd__and2_1 _09692_ (.A(latched_is_lb),
    .B(_04363_),
    .X(_04420_));
 sky130_fd_sc_hd__inv_2 _09693_ (.A(latched_is_lb),
    .Y(_04421_));
 sky130_fd_sc_hd__clkbuf_4 _09694_ (.A(_04031_),
    .X(_04422_));
 sky130_fd_sc_hd__o21a_2 _09695_ (.A1(_04421_),
    .A2(latched_is_lh),
    .B1(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__o221a_1 _09696_ (.A1(net49),
    .A2(_04030_),
    .B1(_04034_),
    .B2(net63),
    .C1(_04423_),
    .X(_04424_));
 sky130_fd_sc_hd__or2_1 _09697_ (.A(_04420_),
    .B(_04424_),
    .X(_04425_));
 sky130_fd_sc_hd__a221o_1 _09698_ (.A1(_04046_),
    .A2(_04419_),
    .B1(_04425_),
    .B2(_03225_),
    .C1(_04266_),
    .X(_04426_));
 sky130_fd_sc_hd__o22a_1 _09699_ (.A1(\irq_pending[8] ),
    .A2(_04007_),
    .B1(_04418_),
    .B2(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__a31o_1 _09700_ (.A1(_04391_),
    .A2(_04394_),
    .A3(_04395_),
    .B1(_04427_),
    .X(_08399_));
 sky130_fd_sc_hd__a22o_1 _09701_ (.A1(\count_instr[9] ),
    .A2(_04145_),
    .B1(_04018_),
    .B2(\count_cycle[41] ),
    .X(_04428_));
 sky130_fd_sc_hd__a221o_1 _09702_ (.A1(\count_instr[41] ),
    .A2(_04016_),
    .B1(\count_cycle[9] ),
    .B2(_04014_),
    .C1(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__clkbuf_8 _09703_ (.A(_04369_),
    .X(_04430_));
 sky130_fd_sc_hd__mux4_1 _09704_ (.A0(\cpuregs.regs[0][9] ),
    .A1(\cpuregs.regs[1][9] ),
    .A2(\cpuregs.regs[2][9] ),
    .A3(\cpuregs.regs[3][9] ),
    .S0(_04325_),
    .S1(_04277_),
    .X(_04431_));
 sky130_fd_sc_hd__or2_1 _09705_ (.A(_04430_),
    .B(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__mux4_1 _09706_ (.A0(\cpuregs.regs[4][9] ),
    .A1(\cpuregs.regs[5][9] ),
    .A2(\cpuregs.regs[6][9] ),
    .A3(\cpuregs.regs[7][9] ),
    .S0(_04291_),
    .S1(_04292_),
    .X(_04433_));
 sky130_fd_sc_hd__o21a_1 _09707_ (.A1(_04211_),
    .A2(_04433_),
    .B1(_04069_),
    .X(_04434_));
 sky130_fd_sc_hd__mux4_1 _09708_ (.A0(\cpuregs.regs[12][9] ),
    .A1(\cpuregs.regs[13][9] ),
    .A2(\cpuregs.regs[14][9] ),
    .A3(\cpuregs.regs[15][9] ),
    .S0(_04274_),
    .S1(_04317_),
    .X(_04435_));
 sky130_fd_sc_hd__mux4_1 _09709_ (.A0(\cpuregs.regs[8][9] ),
    .A1(\cpuregs.regs[9][9] ),
    .A2(\cpuregs.regs[10][9] ),
    .A3(\cpuregs.regs[11][9] ),
    .S0(_04274_),
    .S1(_04317_),
    .X(_04436_));
 sky130_fd_sc_hd__mux2_1 _09710_ (.A0(_04435_),
    .A1(_04436_),
    .S(_04321_),
    .X(_04437_));
 sky130_fd_sc_hd__a221o_1 _09711_ (.A1(_04432_),
    .A2(_04434_),
    .B1(_04437_),
    .B2(_04206_),
    .C1(_04296_),
    .X(_04438_));
 sky130_fd_sc_hd__mux4_1 _09712_ (.A0(\cpuregs.regs[28][9] ),
    .A1(\cpuregs.regs[29][9] ),
    .A2(\cpuregs.regs[30][9] ),
    .A3(\cpuregs.regs[31][9] ),
    .S0(_04217_),
    .S1(_04219_),
    .X(_04439_));
 sky130_fd_sc_hd__mux4_1 _09713_ (.A0(\cpuregs.regs[24][9] ),
    .A1(\cpuregs.regs[25][9] ),
    .A2(\cpuregs.regs[26][9] ),
    .A3(\cpuregs.regs[27][9] ),
    .S0(_04217_),
    .S1(_04219_),
    .X(_04440_));
 sky130_fd_sc_hd__mux2_1 _09714_ (.A0(_04439_),
    .A1(_04440_),
    .S(_04223_),
    .X(_04441_));
 sky130_fd_sc_hd__mux4_1 _09715_ (.A0(\cpuregs.regs[20][9] ),
    .A1(\cpuregs.regs[21][9] ),
    .A2(\cpuregs.regs[22][9] ),
    .A3(\cpuregs.regs[23][9] ),
    .S0(_04072_),
    .S1(_04074_),
    .X(_04442_));
 sky130_fd_sc_hd__mux4_1 _09716_ (.A0(\cpuregs.regs[16][9] ),
    .A1(\cpuregs.regs[17][9] ),
    .A2(\cpuregs.regs[18][9] ),
    .A3(\cpuregs.regs[19][9] ),
    .S0(_04072_),
    .S1(_04074_),
    .X(_04443_));
 sky130_fd_sc_hd__mux2_1 _09717_ (.A0(_04442_),
    .A1(_04443_),
    .S(_04078_),
    .X(_04444_));
 sky130_fd_sc_hd__a21o_1 _09718_ (.A1(_04214_),
    .A2(_04444_),
    .B1(_04081_),
    .X(_04445_));
 sky130_fd_sc_hd__a21o_1 _09719_ (.A1(_04206_),
    .A2(_04441_),
    .B1(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__and3_4 _09720_ (.A(_04133_),
    .B(_04438_),
    .C(_04446_),
    .X(_04447_));
 sky130_fd_sc_hd__clkbuf_4 _09721_ (.A(_04308_),
    .X(_04448_));
 sky130_fd_sc_hd__a221o_1 _09722_ (.A1(\irq_mask[9] ),
    .A2(_04448_),
    .B1(\timer[9] ),
    .B2(_04024_),
    .C1(_04027_),
    .X(_04449_));
 sky130_fd_sc_hd__a21o_1 _09723_ (.A1(_04168_),
    .A2(_04447_),
    .B1(_04449_),
    .X(_04450_));
 sky130_fd_sc_hd__o211a_1 _09724_ (.A1(_04010_),
    .A2(_04429_),
    .B1(_04450_),
    .C1(_04150_),
    .X(_04451_));
 sky130_fd_sc_hd__nor2_1 _09725_ (.A(\reg_pc[9] ),
    .B(\decoded_imm[9] ),
    .Y(_04452_));
 sky130_fd_sc_hd__and2_1 _09726_ (.A(\reg_pc[9] ),
    .B(\decoded_imm[9] ),
    .X(_04453_));
 sky130_fd_sc_hd__a211o_1 _09727_ (.A1(_04392_),
    .A2(_04395_),
    .B1(_04452_),
    .C1(_04453_),
    .X(_04454_));
 sky130_fd_sc_hd__o211ai_1 _09728_ (.A1(_04452_),
    .A2(_04453_),
    .B1(_04392_),
    .C1(_04395_),
    .Y(_04455_));
 sky130_fd_sc_hd__buf_4 _09729_ (.A(net98),
    .X(_04456_));
 sky130_fd_sc_hd__o221a_1 _09730_ (.A1(net50),
    .A2(_04030_),
    .B1(_04034_),
    .B2(net64),
    .C1(_04423_),
    .X(_04457_));
 sky130_fd_sc_hd__or2_1 _09731_ (.A(_04420_),
    .B(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__a221o_1 _09732_ (.A1(_03637_),
    .A2(_04456_),
    .B1(_04458_),
    .B2(_03225_),
    .C1(_04266_),
    .X(_04459_));
 sky130_fd_sc_hd__a31o_1 _09733_ (.A1(_03385_),
    .A2(_04454_),
    .A3(_04455_),
    .B1(_04459_),
    .X(_04460_));
 sky130_fd_sc_hd__o22a_1 _09734_ (.A1(\irq_pending[9] ),
    .A2(_04008_),
    .B1(_04451_),
    .B2(_04460_),
    .X(_08400_));
 sky130_fd_sc_hd__nand2_1 _09735_ (.A(\reg_pc[10] ),
    .B(\decoded_imm[10] ),
    .Y(_04461_));
 sky130_fd_sc_hd__or2_1 _09736_ (.A(\reg_pc[10] ),
    .B(\decoded_imm[10] ),
    .X(_04462_));
 sky130_fd_sc_hd__nand2_1 _09737_ (.A(_04461_),
    .B(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__nand2b_1 _09738_ (.A_N(_04453_),
    .B(_04454_),
    .Y(_04464_));
 sky130_fd_sc_hd__xnor2_1 _09739_ (.A(_04463_),
    .B(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__clkbuf_4 _09740_ (.A(net68),
    .X(_04466_));
 sky130_fd_sc_hd__o221a_1 _09741_ (.A1(net51),
    .A2(_04030_),
    .B1(_04034_),
    .B2(net34),
    .C1(_04423_),
    .X(_04467_));
 sky130_fd_sc_hd__or2_2 _09742_ (.A(_04420_),
    .B(_04467_),
    .X(_04468_));
 sky130_fd_sc_hd__buf_4 _09743_ (.A(_04058_),
    .X(_04469_));
 sky130_fd_sc_hd__buf_4 _09744_ (.A(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__mux4_1 _09745_ (.A0(\cpuregs.regs[24][10] ),
    .A1(\cpuregs.regs[25][10] ),
    .A2(\cpuregs.regs[26][10] ),
    .A3(\cpuregs.regs[27][10] ),
    .S0(_04281_),
    .S1(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__buf_6 _09746_ (.A(_04280_),
    .X(_04472_));
 sky130_fd_sc_hd__clkbuf_8 _09747_ (.A(_04059_),
    .X(_04473_));
 sky130_fd_sc_hd__mux4_1 _09748_ (.A0(\cpuregs.regs[28][10] ),
    .A1(\cpuregs.regs[29][10] ),
    .A2(\cpuregs.regs[30][10] ),
    .A3(\cpuregs.regs[31][10] ),
    .S0(_04472_),
    .S1(_04473_),
    .X(_04474_));
 sky130_fd_sc_hd__mux2_1 _09749_ (.A0(_04471_),
    .A1(_04474_),
    .S(_04430_),
    .X(_04475_));
 sky130_fd_sc_hd__nand2_1 _09750_ (.A(_04054_),
    .B(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__buf_6 _09751_ (.A(_04084_),
    .X(_04477_));
 sky130_fd_sc_hd__buf_4 _09752_ (.A(_04086_),
    .X(_04478_));
 sky130_fd_sc_hd__mux4_1 _09753_ (.A0(\cpuregs.regs[20][10] ),
    .A1(\cpuregs.regs[21][10] ),
    .A2(\cpuregs.regs[22][10] ),
    .A3(\cpuregs.regs[23][10] ),
    .S0(_04477_),
    .S1(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__mux4_1 _09754_ (.A0(\cpuregs.regs[16][10] ),
    .A1(\cpuregs.regs[17][10] ),
    .A2(\cpuregs.regs[18][10] ),
    .A3(\cpuregs.regs[19][10] ),
    .S0(_04085_),
    .S1(_04087_),
    .X(_04480_));
 sky130_fd_sc_hd__mux2_1 _09755_ (.A0(_04479_),
    .A1(_04480_),
    .S(_04078_),
    .X(_04481_));
 sky130_fd_sc_hd__a21oi_1 _09756_ (.A1(_04070_),
    .A2(_04481_),
    .B1(_04082_),
    .Y(_04482_));
 sky130_fd_sc_hd__buf_4 _09757_ (.A(_04069_),
    .X(_04483_));
 sky130_fd_sc_hd__mux4_1 _09758_ (.A0(\cpuregs.regs[4][10] ),
    .A1(\cpuregs.regs[5][10] ),
    .A2(\cpuregs.regs[6][10] ),
    .A3(\cpuregs.regs[7][10] ),
    .S0(_04232_),
    .S1(_04233_),
    .X(_04484_));
 sky130_fd_sc_hd__mux4_1 _09759_ (.A0(\cpuregs.regs[0][10] ),
    .A1(\cpuregs.regs[1][10] ),
    .A2(\cpuregs.regs[2][10] ),
    .A3(\cpuregs.regs[3][10] ),
    .S0(_04232_),
    .S1(_04233_),
    .X(_04485_));
 sky130_fd_sc_hd__mux2_1 _09760_ (.A0(_04484_),
    .A1(_04485_),
    .S(_04121_),
    .X(_04486_));
 sky130_fd_sc_hd__buf_6 _09761_ (.A(_04055_),
    .X(_04487_));
 sky130_fd_sc_hd__mux4_1 _09762_ (.A0(\cpuregs.regs[12][10] ),
    .A1(\cpuregs.regs[13][10] ),
    .A2(\cpuregs.regs[14][10] ),
    .A3(\cpuregs.regs[15][10] ),
    .S0(_04487_),
    .S1(_04469_),
    .X(_04488_));
 sky130_fd_sc_hd__mux4_1 _09763_ (.A0(\cpuregs.regs[8][10] ),
    .A1(\cpuregs.regs[9][10] ),
    .A2(\cpuregs.regs[10][10] ),
    .A3(\cpuregs.regs[11][10] ),
    .S0(_04487_),
    .S1(_04469_),
    .X(_04489_));
 sky130_fd_sc_hd__mux2_1 _09764_ (.A0(_04488_),
    .A1(_04489_),
    .S(_04320_),
    .X(_04490_));
 sky130_fd_sc_hd__a21o_1 _09765_ (.A1(_04053_),
    .A2(_04490_),
    .B1(_04095_),
    .X(_04491_));
 sky130_fd_sc_hd__a21oi_1 _09766_ (.A1(_04483_),
    .A2(_04486_),
    .B1(_04491_),
    .Y(_04492_));
 sky130_fd_sc_hd__a211o_2 _09767_ (.A1(_04476_),
    .A2(_04482_),
    .B1(_04100_),
    .C1(_04492_),
    .X(_04493_));
 sky130_fd_sc_hd__nor2_1 _09768_ (.A(_04051_),
    .B(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hd__a221o_1 _09769_ (.A1(\irq_mask[10] ),
    .A2(_04021_),
    .B1(\timer[10] ),
    .B2(_04023_),
    .C1(_04188_),
    .X(_04495_));
 sky130_fd_sc_hd__a22o_1 _09770_ (.A1(\count_instr[42] ),
    .A2(instr_rdinstrh),
    .B1(instr_rdinstr),
    .B2(\count_instr[10] ),
    .X(_04496_));
 sky130_fd_sc_hd__a211o_1 _09771_ (.A1(_04017_),
    .A2(\count_cycle[42] ),
    .B1(_03252_),
    .C1(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__a21o_1 _09772_ (.A1(\count_cycle[10] ),
    .A2(_04013_),
    .B1(_04497_),
    .X(_04498_));
 sky130_fd_sc_hd__o211a_1 _09773_ (.A1(_04494_),
    .A2(_04495_),
    .B1(_04498_),
    .C1(_04149_),
    .X(_04499_));
 sky130_fd_sc_hd__a221o_1 _09774_ (.A1(_03638_),
    .A2(_04466_),
    .B1(_04468_),
    .B2(_03226_),
    .C1(_04499_),
    .X(_04500_));
 sky130_fd_sc_hd__a221o_1 _09775_ (.A1(\irq_pending[10] ),
    .A2(_04049_),
    .B1(_04465_),
    .B2(_03385_),
    .C1(_04500_),
    .X(_08370_));
 sky130_fd_sc_hd__nor2_1 _09776_ (.A(\reg_pc[11] ),
    .B(\decoded_imm[11] ),
    .Y(_04501_));
 sky130_fd_sc_hd__and2_1 _09777_ (.A(\reg_pc[11] ),
    .B(\decoded_imm[11] ),
    .X(_04502_));
 sky130_fd_sc_hd__a21boi_1 _09778_ (.A1(_04462_),
    .A2(_04464_),
    .B1_N(_04461_),
    .Y(_04503_));
 sky130_fd_sc_hd__or3_1 _09779_ (.A(_04501_),
    .B(_04502_),
    .C(_04503_),
    .X(_04504_));
 sky130_fd_sc_hd__o21ai_1 _09780_ (.A1(_04501_),
    .A2(_04502_),
    .B1(_04503_),
    .Y(_04505_));
 sky130_fd_sc_hd__o221a_1 _09781_ (.A1(net52),
    .A2(_04030_),
    .B1(_04034_),
    .B2(net35),
    .C1(_04423_),
    .X(_04506_));
 sky130_fd_sc_hd__o21a_2 _09782_ (.A1(_04420_),
    .A2(_04506_),
    .B1(_03225_),
    .X(_04507_));
 sky130_fd_sc_hd__mux4_1 _09783_ (.A0(\cpuregs.regs[12][11] ),
    .A1(\cpuregs.regs[13][11] ),
    .A2(\cpuregs.regs[14][11] ),
    .A3(\cpuregs.regs[15][11] ),
    .S0(_04282_),
    .S1(_04285_),
    .X(_04508_));
 sky130_fd_sc_hd__mux4_1 _09784_ (.A0(\cpuregs.regs[8][11] ),
    .A1(\cpuregs.regs[9][11] ),
    .A2(\cpuregs.regs[10][11] ),
    .A3(\cpuregs.regs[11][11] ),
    .S0(_04282_),
    .S1(_04285_),
    .X(_04509_));
 sky130_fd_sc_hd__mux2_1 _09785_ (.A0(_04508_),
    .A1(_04509_),
    .S(_04287_),
    .X(_04510_));
 sky130_fd_sc_hd__mux4_1 _09786_ (.A0(\cpuregs.regs[4][11] ),
    .A1(\cpuregs.regs[5][11] ),
    .A2(\cpuregs.regs[6][11] ),
    .A3(\cpuregs.regs[7][11] ),
    .S0(_04274_),
    .S1(_04317_),
    .X(_04511_));
 sky130_fd_sc_hd__buf_8 _09787_ (.A(_04273_),
    .X(_04512_));
 sky130_fd_sc_hd__clkbuf_8 _09788_ (.A(_04283_),
    .X(_04513_));
 sky130_fd_sc_hd__mux4_1 _09789_ (.A0(\cpuregs.regs[0][11] ),
    .A1(\cpuregs.regs[1][11] ),
    .A2(\cpuregs.regs[2][11] ),
    .A3(\cpuregs.regs[3][11] ),
    .S0(_04512_),
    .S1(_04513_),
    .X(_04514_));
 sky130_fd_sc_hd__mux2_1 _09790_ (.A0(_04511_),
    .A1(_04514_),
    .S(_04321_),
    .X(_04515_));
 sky130_fd_sc_hd__a21o_1 _09791_ (.A1(_04289_),
    .A2(_04515_),
    .B1(_04296_),
    .X(_04516_));
 sky130_fd_sc_hd__a21oi_2 _09792_ (.A1(_04272_),
    .A2(_04510_),
    .B1(_04516_),
    .Y(_04517_));
 sky130_fd_sc_hd__mux4_1 _09793_ (.A0(\cpuregs.regs[28][11] ),
    .A1(\cpuregs.regs[29][11] ),
    .A2(\cpuregs.regs[30][11] ),
    .A3(\cpuregs.regs[31][11] ),
    .S0(_04282_),
    .S1(_04285_),
    .X(_04518_));
 sky130_fd_sc_hd__mux4_1 _09794_ (.A0(\cpuregs.regs[24][11] ),
    .A1(\cpuregs.regs[25][11] ),
    .A2(\cpuregs.regs[26][11] ),
    .A3(\cpuregs.regs[27][11] ),
    .S0(_04282_),
    .S1(_04285_),
    .X(_04519_));
 sky130_fd_sc_hd__mux2_1 _09795_ (.A0(_04518_),
    .A1(_04519_),
    .S(_04287_),
    .X(_04520_));
 sky130_fd_sc_hd__mux4_1 _09796_ (.A0(\cpuregs.regs[20][11] ),
    .A1(\cpuregs.regs[21][11] ),
    .A2(\cpuregs.regs[22][11] ),
    .A3(\cpuregs.regs[23][11] ),
    .S0(_04325_),
    .S1(_04277_),
    .X(_04521_));
 sky130_fd_sc_hd__mux4_1 _09797_ (.A0(\cpuregs.regs[16][11] ),
    .A1(\cpuregs.regs[17][11] ),
    .A2(\cpuregs.regs[18][11] ),
    .A3(\cpuregs.regs[19][11] ),
    .S0(_04325_),
    .S1(_04277_),
    .X(_04522_));
 sky130_fd_sc_hd__mux2_1 _09798_ (.A0(_04521_),
    .A1(_04522_),
    .S(_04321_),
    .X(_04523_));
 sky130_fd_sc_hd__a21o_1 _09799_ (.A1(_04289_),
    .A2(_04523_),
    .B1(_04225_),
    .X(_04524_));
 sky130_fd_sc_hd__a21oi_2 _09800_ (.A1(_04272_),
    .A2(_04520_),
    .B1(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__nor3_4 _09801_ (.A(_04227_),
    .B(_04517_),
    .C(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__a221o_1 _09802_ (.A1(\irq_mask[11] ),
    .A2(_04308_),
    .B1(\timer[11] ),
    .B2(instr_timer),
    .C1(_04025_),
    .X(_04527_));
 sky130_fd_sc_hd__a21o_1 _09803_ (.A1(instr_retirq),
    .A2(_04526_),
    .B1(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__a22o_1 _09804_ (.A1(\count_instr[43] ),
    .A2(instr_rdinstrh),
    .B1(instr_rdcycleh),
    .B2(\count_cycle[43] ),
    .X(_04529_));
 sky130_fd_sc_hd__a211o_1 _09805_ (.A1(\count_instr[11] ),
    .A2(_04011_),
    .B1(_03252_),
    .C1(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__a21o_1 _09806_ (.A1(\count_cycle[11] ),
    .A2(_04165_),
    .B1(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__buf_4 _09807_ (.A(net69),
    .X(_04532_));
 sky130_fd_sc_hd__a32o_1 _09808_ (.A1(_04149_),
    .A2(_04528_),
    .A3(_04531_),
    .B1(_04046_),
    .B2(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__a211o_1 _09809_ (.A1(\irq_pending[11] ),
    .A2(_04049_),
    .B1(_04507_),
    .C1(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__a31o_1 _09810_ (.A1(_04391_),
    .A2(_04504_),
    .A3(_04505_),
    .B1(_04534_),
    .X(_08371_));
 sky130_fd_sc_hd__nand2_1 _09811_ (.A(\reg_pc[12] ),
    .B(\decoded_imm[12] ),
    .Y(_04535_));
 sky130_fd_sc_hd__or2_1 _09812_ (.A(\reg_pc[12] ),
    .B(\decoded_imm[12] ),
    .X(_04536_));
 sky130_fd_sc_hd__nand2_1 _09813_ (.A(_04535_),
    .B(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__nand2_1 _09814_ (.A(\reg_pc[11] ),
    .B(\decoded_imm[11] ),
    .Y(_04538_));
 sky130_fd_sc_hd__o211ai_1 _09815_ (.A1(_04501_),
    .A2(_04503_),
    .B1(_04537_),
    .C1(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__or4b_1 _09816_ (.A(_04463_),
    .B(_04501_),
    .C(_04502_),
    .D_N(_04464_),
    .X(_04540_));
 sky130_fd_sc_hd__or2_1 _09817_ (.A(_04461_),
    .B(_04501_),
    .X(_04541_));
 sky130_fd_sc_hd__a31o_1 _09818_ (.A1(_04538_),
    .A2(_04540_),
    .A3(_04541_),
    .B1(_04537_),
    .X(_04542_));
 sky130_fd_sc_hd__a22o_1 _09819_ (.A1(\count_instr[12] ),
    .A2(_04011_),
    .B1(_04017_),
    .B2(\count_cycle[44] ),
    .X(_04543_));
 sky130_fd_sc_hd__a221o_1 _09820_ (.A1(\count_instr[44] ),
    .A2(_04016_),
    .B1(\count_cycle[12] ),
    .B2(_04013_),
    .C1(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__mux4_1 _09821_ (.A0(\cpuregs.regs[8][12] ),
    .A1(\cpuregs.regs[9][12] ),
    .A2(\cpuregs.regs[10][12] ),
    .A3(\cpuregs.regs[11][12] ),
    .S0(_04085_),
    .S1(_04087_),
    .X(_04545_));
 sky130_fd_sc_hd__mux4_1 _09822_ (.A0(\cpuregs.regs[12][12] ),
    .A1(\cpuregs.regs[13][12] ),
    .A2(\cpuregs.regs[14][12] ),
    .A3(\cpuregs.regs[15][12] ),
    .S0(_04085_),
    .S1(_04087_),
    .X(_04546_));
 sky130_fd_sc_hd__mux2_1 _09823_ (.A0(_04545_),
    .A1(_04546_),
    .S(_04369_),
    .X(_04547_));
 sky130_fd_sc_hd__nand2_1 _09824_ (.A(_04231_),
    .B(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__mux4_1 _09825_ (.A0(\cpuregs.regs[4][12] ),
    .A1(\cpuregs.regs[5][12] ),
    .A2(\cpuregs.regs[6][12] ),
    .A3(\cpuregs.regs[7][12] ),
    .S0(_04216_),
    .S1(_04376_),
    .X(_04549_));
 sky130_fd_sc_hd__mux4_1 _09826_ (.A0(\cpuregs.regs[0][12] ),
    .A1(\cpuregs.regs[1][12] ),
    .A2(\cpuregs.regs[2][12] ),
    .A3(\cpuregs.regs[3][12] ),
    .S0(_04216_),
    .S1(_04376_),
    .X(_04550_));
 sky130_fd_sc_hd__mux2_1 _09827_ (.A0(_04549_),
    .A1(_04550_),
    .S(_04222_),
    .X(_04551_));
 sky130_fd_sc_hd__a21oi_1 _09828_ (.A1(_04214_),
    .A2(_04551_),
    .B1(_04237_),
    .Y(_04552_));
 sky130_fd_sc_hd__mux4_1 _09829_ (.A0(\cpuregs.regs[24][12] ),
    .A1(\cpuregs.regs[25][12] ),
    .A2(\cpuregs.regs[26][12] ),
    .A3(\cpuregs.regs[27][12] ),
    .S0(_04329_),
    .S1(_04218_),
    .X(_04553_));
 sky130_fd_sc_hd__mux4_1 _09830_ (.A0(\cpuregs.regs[28][12] ),
    .A1(\cpuregs.regs[29][12] ),
    .A2(\cpuregs.regs[30][12] ),
    .A3(\cpuregs.regs[31][12] ),
    .S0(_04329_),
    .S1(_04376_),
    .X(_04554_));
 sky130_fd_sc_hd__mux2_1 _09831_ (.A0(_04553_),
    .A1(_04554_),
    .S(_04369_),
    .X(_04555_));
 sky130_fd_sc_hd__mux4_1 _09832_ (.A0(\cpuregs.regs[20][12] ),
    .A1(\cpuregs.regs[21][12] ),
    .A2(\cpuregs.regs[22][12] ),
    .A3(\cpuregs.regs[23][12] ),
    .S0(_04084_),
    .S1(_04086_),
    .X(_04556_));
 sky130_fd_sc_hd__mux4_1 _09833_ (.A0(\cpuregs.regs[16][12] ),
    .A1(\cpuregs.regs[17][12] ),
    .A2(\cpuregs.regs[18][12] ),
    .A3(\cpuregs.regs[19][12] ),
    .S0(_04071_),
    .S1(_04073_),
    .X(_04557_));
 sky130_fd_sc_hd__mux2_1 _09834_ (.A0(_04556_),
    .A1(_04557_),
    .S(_04077_),
    .X(_04558_));
 sky130_fd_sc_hd__a21o_1 _09835_ (.A1(_04068_),
    .A2(_04558_),
    .B1(_04081_),
    .X(_04559_));
 sky130_fd_sc_hd__a21oi_1 _09836_ (.A1(_04328_),
    .A2(_04555_),
    .B1(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__a211o_4 _09837_ (.A1(_04548_),
    .A2(_04552_),
    .B1(_04560_),
    .C1(net300),
    .X(_04561_));
 sky130_fd_sc_hd__inv_2 _09838_ (.A(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__a221o_1 _09839_ (.A1(\irq_mask[12] ),
    .A2(_04308_),
    .B1(\timer[12] ),
    .B2(instr_timer),
    .C1(_04026_),
    .X(_04563_));
 sky130_fd_sc_hd__a21o_1 _09840_ (.A1(_04271_),
    .A2(_04562_),
    .B1(_04563_),
    .X(_04564_));
 sky130_fd_sc_hd__o211a_1 _09841_ (.A1(_04268_),
    .A2(_04544_),
    .B1(_04564_),
    .C1(_04149_),
    .X(_04565_));
 sky130_fd_sc_hd__clkbuf_4 _09842_ (.A(net70),
    .X(_04566_));
 sky130_fd_sc_hd__o221a_1 _09843_ (.A1(net53),
    .A2(_04030_),
    .B1(_04034_),
    .B2(net36),
    .C1(_04423_),
    .X(_04567_));
 sky130_fd_sc_hd__or2_1 _09844_ (.A(_04420_),
    .B(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__a221o_1 _09845_ (.A1(_03637_),
    .A2(_04566_),
    .B1(_04568_),
    .B2(_03225_),
    .C1(_04266_),
    .X(_04569_));
 sky130_fd_sc_hd__o22a_1 _09846_ (.A1(\irq_pending[12] ),
    .A2(_04007_),
    .B1(_04565_),
    .B2(_04569_),
    .X(_04570_));
 sky130_fd_sc_hd__a31o_1 _09847_ (.A1(_04391_),
    .A2(_04539_),
    .A3(_04542_),
    .B1(_04570_),
    .X(_08372_));
 sky130_fd_sc_hd__a22o_1 _09848_ (.A1(\count_instr[45] ),
    .A2(_04016_),
    .B1(_04012_),
    .B2(\count_instr[13] ),
    .X(_04571_));
 sky130_fd_sc_hd__a221o_1 _09849_ (.A1(_04018_),
    .A2(\count_cycle[45] ),
    .B1(_04014_),
    .B2(\count_cycle[13] ),
    .C1(_04571_),
    .X(_04572_));
 sky130_fd_sc_hd__mux4_1 _09850_ (.A0(\cpuregs.regs[20][13] ),
    .A1(\cpuregs.regs[21][13] ),
    .A2(\cpuregs.regs[22][13] ),
    .A3(\cpuregs.regs[23][13] ),
    .S0(_04512_),
    .S1(_04513_),
    .X(_04573_));
 sky130_fd_sc_hd__mux4_1 _09851_ (.A0(\cpuregs.regs[16][13] ),
    .A1(\cpuregs.regs[17][13] ),
    .A2(\cpuregs.regs[18][13] ),
    .A3(\cpuregs.regs[19][13] ),
    .S0(_04512_),
    .S1(_04513_),
    .X(_04574_));
 sky130_fd_sc_hd__buf_8 _09852_ (.A(_04320_),
    .X(_04575_));
 sky130_fd_sc_hd__mux2_1 _09853_ (.A0(_04573_),
    .A1(_04574_),
    .S(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__nand2_1 _09854_ (.A(_04483_),
    .B(_04576_),
    .Y(_04577_));
 sky130_fd_sc_hd__mux4_1 _09855_ (.A0(\cpuregs.regs[28][13] ),
    .A1(\cpuregs.regs[29][13] ),
    .A2(\cpuregs.regs[30][13] ),
    .A3(\cpuregs.regs[31][13] ),
    .S0(_04512_),
    .S1(_04513_),
    .X(_04578_));
 sky130_fd_sc_hd__buf_8 _09856_ (.A(_04487_),
    .X(_04579_));
 sky130_fd_sc_hd__mux4_1 _09857_ (.A0(\cpuregs.regs[24][13] ),
    .A1(\cpuregs.regs[25][13] ),
    .A2(\cpuregs.regs[26][13] ),
    .A3(\cpuregs.regs[27][13] ),
    .S0(_04579_),
    .S1(_04284_),
    .X(_04580_));
 sky130_fd_sc_hd__mux2_1 _09858_ (.A0(_04578_),
    .A1(_04580_),
    .S(_04575_),
    .X(_04581_));
 sky130_fd_sc_hd__nand2_1 _09859_ (.A(_04206_),
    .B(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__mux4_1 _09860_ (.A0(\cpuregs.regs[0][13] ),
    .A1(\cpuregs.regs[1][13] ),
    .A2(\cpuregs.regs[2][13] ),
    .A3(\cpuregs.regs[3][13] ),
    .S0(_04487_),
    .S1(_04469_),
    .X(_04583_));
 sky130_fd_sc_hd__or2_1 _09861_ (.A(_04369_),
    .B(_04583_),
    .X(_04584_));
 sky130_fd_sc_hd__mux4_1 _09862_ (.A0(\cpuregs.regs[4][13] ),
    .A1(\cpuregs.regs[5][13] ),
    .A2(\cpuregs.regs[6][13] ),
    .A3(\cpuregs.regs[7][13] ),
    .S0(_04273_),
    .S1(_04283_),
    .X(_04585_));
 sky130_fd_sc_hd__o21a_1 _09863_ (.A1(_04320_),
    .A2(_04585_),
    .B1(_04068_),
    .X(_04586_));
 sky130_fd_sc_hd__mux4_1 _09864_ (.A0(\cpuregs.regs[12][13] ),
    .A1(\cpuregs.regs[13][13] ),
    .A2(\cpuregs.regs[14][13] ),
    .A3(\cpuregs.regs[15][13] ),
    .S0(_04280_),
    .S1(_04059_),
    .X(_04587_));
 sky130_fd_sc_hd__mux4_1 _09865_ (.A0(\cpuregs.regs[8][13] ),
    .A1(\cpuregs.regs[9][13] ),
    .A2(\cpuregs.regs[10][13] ),
    .A3(\cpuregs.regs[11][13] ),
    .S0(_04280_),
    .S1(_04091_),
    .X(_04588_));
 sky130_fd_sc_hd__mux2_1 _09866_ (.A0(_04587_),
    .A1(_04588_),
    .S(_04064_),
    .X(_04589_));
 sky130_fd_sc_hd__a221o_1 _09867_ (.A1(_04584_),
    .A2(_04586_),
    .B1(_04589_),
    .B2(_04053_),
    .C1(_04095_),
    .X(_04590_));
 sky130_fd_sc_hd__nand2_1 _09868_ (.A(_04133_),
    .B(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__a31o_2 _09869_ (.A1(_04296_),
    .A2(_04577_),
    .A3(_04582_),
    .B1(_04591_),
    .X(_04592_));
 sky130_fd_sc_hd__inv_2 _09870_ (.A(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__a221o_1 _09871_ (.A1(\irq_mask[13] ),
    .A2(_04448_),
    .B1(\timer[13] ),
    .B2(_04024_),
    .C1(_04027_),
    .X(_04594_));
 sky130_fd_sc_hd__a21o_1 _09872_ (.A1(_04168_),
    .A2(_04593_),
    .B1(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__o211a_1 _09873_ (.A1(_04010_),
    .A2(_04572_),
    .B1(_04595_),
    .C1(_04150_),
    .X(_04596_));
 sky130_fd_sc_hd__nand2_1 _09874_ (.A(\reg_pc[13] ),
    .B(\decoded_imm[13] ),
    .Y(_04597_));
 sky130_fd_sc_hd__or2_1 _09875_ (.A(\reg_pc[13] ),
    .B(\decoded_imm[13] ),
    .X(_04598_));
 sky130_fd_sc_hd__nand2_1 _09876_ (.A(_04597_),
    .B(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__a21o_1 _09877_ (.A1(_04535_),
    .A2(_04542_),
    .B1(_04599_),
    .X(_04600_));
 sky130_fd_sc_hd__nand3_1 _09878_ (.A(_04535_),
    .B(_04542_),
    .C(_04599_),
    .Y(_04601_));
 sky130_fd_sc_hd__clkbuf_4 _09879_ (.A(net71),
    .X(_04602_));
 sky130_fd_sc_hd__o221a_1 _09880_ (.A1(net54),
    .A2(_04030_),
    .B1(_04034_),
    .B2(net37),
    .C1(_04423_),
    .X(_04603_));
 sky130_fd_sc_hd__or2_2 _09881_ (.A(_04420_),
    .B(_04603_),
    .X(_04604_));
 sky130_fd_sc_hd__a221o_1 _09882_ (.A1(_03637_),
    .A2(_04602_),
    .B1(_04604_),
    .B2(_03225_),
    .C1(_04266_),
    .X(_04605_));
 sky130_fd_sc_hd__a31o_1 _09883_ (.A1(_03385_),
    .A2(_04600_),
    .A3(_04601_),
    .B1(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__o22a_1 _09884_ (.A1(\irq_pending[13] ),
    .A2(_04008_),
    .B1(_04596_),
    .B2(_04606_),
    .X(_08373_));
 sky130_fd_sc_hd__xnor2_1 _09885_ (.A(\reg_pc[14] ),
    .B(\decoded_imm[14] ),
    .Y(_04607_));
 sky130_fd_sc_hd__a21oi_1 _09886_ (.A1(_04597_),
    .A2(_04600_),
    .B1(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__a31o_1 _09887_ (.A1(_04597_),
    .A2(_04600_),
    .A3(_04607_),
    .B1(_04156_),
    .X(_04609_));
 sky130_fd_sc_hd__nor2_1 _09888_ (.A(_04608_),
    .B(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__clkbuf_4 _09889_ (.A(net72),
    .X(_04611_));
 sky130_fd_sc_hd__o221a_1 _09890_ (.A1(net56),
    .A2(_04030_),
    .B1(_04034_),
    .B2(net38),
    .C1(_04423_),
    .X(_04612_));
 sky130_fd_sc_hd__or2_2 _09891_ (.A(_04420_),
    .B(_04612_),
    .X(_04613_));
 sky130_fd_sc_hd__mux4_1 _09892_ (.A0(\cpuregs.regs[4][14] ),
    .A1(\cpuregs.regs[5][14] ),
    .A2(\cpuregs.regs[6][14] ),
    .A3(\cpuregs.regs[7][14] ),
    .S0(_04290_),
    .S1(_04276_),
    .X(_04614_));
 sky130_fd_sc_hd__mux4_1 _09893_ (.A0(\cpuregs.regs[0][14] ),
    .A1(\cpuregs.regs[1][14] ),
    .A2(\cpuregs.regs[2][14] ),
    .A3(\cpuregs.regs[3][14] ),
    .S0(_04290_),
    .S1(_04276_),
    .X(_04615_));
 sky130_fd_sc_hd__mux2_1 _09894_ (.A0(_04614_),
    .A1(_04615_),
    .S(_04222_),
    .X(_04616_));
 sky130_fd_sc_hd__nand2_1 _09895_ (.A(_04214_),
    .B(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__mux4_1 _09896_ (.A0(\cpuregs.regs[12][14] ),
    .A1(\cpuregs.regs[13][14] ),
    .A2(\cpuregs.regs[14][14] ),
    .A3(\cpuregs.regs[15][14] ),
    .S0(_04216_),
    .S1(_04376_),
    .X(_04618_));
 sky130_fd_sc_hd__mux4_1 _09897_ (.A0(\cpuregs.regs[8][14] ),
    .A1(\cpuregs.regs[9][14] ),
    .A2(\cpuregs.regs[10][14] ),
    .A3(\cpuregs.regs[11][14] ),
    .S0(_04216_),
    .S1(_04376_),
    .X(_04619_));
 sky130_fd_sc_hd__mux2_1 _09898_ (.A0(_04618_),
    .A1(_04619_),
    .S(_04222_),
    .X(_04620_));
 sky130_fd_sc_hd__nand2_1 _09899_ (.A(_04328_),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__mux4_1 _09900_ (.A0(\cpuregs.regs[20][14] ),
    .A1(\cpuregs.regs[21][14] ),
    .A2(\cpuregs.regs[22][14] ),
    .A3(\cpuregs.regs[23][14] ),
    .S0(_04329_),
    .S1(_04218_),
    .X(_04622_));
 sky130_fd_sc_hd__mux4_1 _09901_ (.A0(\cpuregs.regs[16][14] ),
    .A1(\cpuregs.regs[17][14] ),
    .A2(\cpuregs.regs[18][14] ),
    .A3(\cpuregs.regs[19][14] ),
    .S0(_04329_),
    .S1(_04218_),
    .X(_04623_));
 sky130_fd_sc_hd__mux2_1 _09902_ (.A0(_04622_),
    .A1(_04623_),
    .S(_04078_),
    .X(_04624_));
 sky130_fd_sc_hd__nand2_1 _09903_ (.A(_04070_),
    .B(_04624_),
    .Y(_04625_));
 sky130_fd_sc_hd__mux4_1 _09904_ (.A0(\cpuregs.regs[24][14] ),
    .A1(\cpuregs.regs[25][14] ),
    .A2(\cpuregs.regs[26][14] ),
    .A3(\cpuregs.regs[27][14] ),
    .S0(_04290_),
    .S1(_04276_),
    .X(_04626_));
 sky130_fd_sc_hd__mux4_1 _09905_ (.A0(\cpuregs.regs[28][14] ),
    .A1(\cpuregs.regs[29][14] ),
    .A2(\cpuregs.regs[30][14] ),
    .A3(\cpuregs.regs[31][14] ),
    .S0(_04290_),
    .S1(_04276_),
    .X(_04627_));
 sky130_fd_sc_hd__mux2_1 _09906_ (.A0(_04626_),
    .A1(_04627_),
    .S(_04369_),
    .X(_04628_));
 sky130_fd_sc_hd__a21oi_1 _09907_ (.A1(_04328_),
    .A2(_04628_),
    .B1(_04081_),
    .Y(_04629_));
 sky130_fd_sc_hd__a32o_1 _09908_ (.A1(_04082_),
    .A2(_04617_),
    .A3(_04621_),
    .B1(_04625_),
    .B2(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__or2_4 _09909_ (.A(_04227_),
    .B(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__nor2_1 _09910_ (.A(_04051_),
    .B(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__a221o_1 _09911_ (.A1(\irq_mask[14] ),
    .A2(_04021_),
    .B1(\timer[14] ),
    .B2(_04187_),
    .C1(_04188_),
    .X(_04633_));
 sky130_fd_sc_hd__a22o_1 _09912_ (.A1(\count_instr[46] ),
    .A2(instr_rdinstrh),
    .B1(instr_rdinstr),
    .B2(\count_instr[14] ),
    .X(_04634_));
 sky130_fd_sc_hd__a211o_1 _09913_ (.A1(_04017_),
    .A2(\count_cycle[46] ),
    .B1(_03252_),
    .C1(_04634_),
    .X(_04635_));
 sky130_fd_sc_hd__a21o_1 _09914_ (.A1(\count_cycle[14] ),
    .A2(_04165_),
    .B1(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__o211a_1 _09915_ (.A1(_04632_),
    .A2(_04633_),
    .B1(_04636_),
    .C1(_04149_),
    .X(_04637_));
 sky130_fd_sc_hd__a221o_1 _09916_ (.A1(_03638_),
    .A2(_04611_),
    .B1(_04613_),
    .B2(_03226_),
    .C1(_04637_),
    .X(_04638_));
 sky130_fd_sc_hd__a211o_1 _09917_ (.A1(\irq_pending[14] ),
    .A2(_04049_),
    .B1(_04610_),
    .C1(_04638_),
    .X(_08374_));
 sky130_fd_sc_hd__xnor2_1 _09918_ (.A(\reg_pc[15] ),
    .B(\decoded_imm[15] ),
    .Y(_04639_));
 sky130_fd_sc_hd__a21o_1 _09919_ (.A1(\reg_pc[14] ),
    .A2(\decoded_imm[14] ),
    .B1(_04608_),
    .X(_04640_));
 sky130_fd_sc_hd__xnor2_1 _09920_ (.A(_04639_),
    .B(_04640_),
    .Y(_04641_));
 sky130_fd_sc_hd__clkbuf_4 _09921_ (.A(net73),
    .X(_04642_));
 sky130_fd_sc_hd__mux4_1 _09922_ (.A0(\cpuregs.regs[20][15] ),
    .A1(\cpuregs.regs[21][15] ),
    .A2(\cpuregs.regs[22][15] ),
    .A3(\cpuregs.regs[23][15] ),
    .S0(_04281_),
    .S1(_04470_),
    .X(_04643_));
 sky130_fd_sc_hd__mux4_1 _09923_ (.A0(\cpuregs.regs[16][15] ),
    .A1(\cpuregs.regs[17][15] ),
    .A2(\cpuregs.regs[18][15] ),
    .A3(\cpuregs.regs[19][15] ),
    .S0(_04472_),
    .S1(_04473_),
    .X(_04644_));
 sky130_fd_sc_hd__mux2_1 _09924_ (.A0(_04643_),
    .A1(_04644_),
    .S(_04065_),
    .X(_04645_));
 sky130_fd_sc_hd__nand2_1 _09925_ (.A(_04483_),
    .B(_04645_),
    .Y(_04646_));
 sky130_fd_sc_hd__mux4_1 _09926_ (.A0(\cpuregs.regs[28][15] ),
    .A1(\cpuregs.regs[29][15] ),
    .A2(\cpuregs.regs[30][15] ),
    .A3(\cpuregs.regs[31][15] ),
    .S0(_04477_),
    .S1(_04478_),
    .X(_04647_));
 sky130_fd_sc_hd__mux4_1 _09927_ (.A0(\cpuregs.regs[24][15] ),
    .A1(\cpuregs.regs[25][15] ),
    .A2(\cpuregs.regs[26][15] ),
    .A3(\cpuregs.regs[27][15] ),
    .S0(_04085_),
    .S1(_04087_),
    .X(_04648_));
 sky130_fd_sc_hd__mux2_1 _09928_ (.A0(_04647_),
    .A1(_04648_),
    .S(_04121_),
    .X(_04649_));
 sky130_fd_sc_hd__a21oi_1 _09929_ (.A1(_04231_),
    .A2(_04649_),
    .B1(_04082_),
    .Y(_04650_));
 sky130_fd_sc_hd__mux4_1 _09930_ (.A0(\cpuregs.regs[4][15] ),
    .A1(\cpuregs.regs[5][15] ),
    .A2(\cpuregs.regs[6][15] ),
    .A3(\cpuregs.regs[7][15] ),
    .S0(_04232_),
    .S1(_04233_),
    .X(_04651_));
 sky130_fd_sc_hd__mux4_1 _09931_ (.A0(\cpuregs.regs[0][15] ),
    .A1(\cpuregs.regs[1][15] ),
    .A2(\cpuregs.regs[2][15] ),
    .A3(\cpuregs.regs[3][15] ),
    .S0(_04232_),
    .S1(_04233_),
    .X(_04652_));
 sky130_fd_sc_hd__mux2_1 _09932_ (.A0(_04651_),
    .A1(_04652_),
    .S(_04121_),
    .X(_04653_));
 sky130_fd_sc_hd__mux4_1 _09933_ (.A0(\cpuregs.regs[12][15] ),
    .A1(\cpuregs.regs[13][15] ),
    .A2(\cpuregs.regs[14][15] ),
    .A3(\cpuregs.regs[15][15] ),
    .S0(_04487_),
    .S1(_04469_),
    .X(_04654_));
 sky130_fd_sc_hd__mux4_1 _09934_ (.A0(\cpuregs.regs[8][15] ),
    .A1(\cpuregs.regs[9][15] ),
    .A2(\cpuregs.regs[10][15] ),
    .A3(\cpuregs.regs[11][15] ),
    .S0(_04487_),
    .S1(_04469_),
    .X(_04655_));
 sky130_fd_sc_hd__mux2_1 _09935_ (.A0(_04654_),
    .A1(_04655_),
    .S(_04320_),
    .X(_04656_));
 sky130_fd_sc_hd__a21o_1 _09936_ (.A1(_04053_),
    .A2(_04656_),
    .B1(_04095_),
    .X(_04657_));
 sky130_fd_sc_hd__a21oi_1 _09937_ (.A1(_04483_),
    .A2(_04653_),
    .B1(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__a211o_2 _09938_ (.A1(_04646_),
    .A2(_04650_),
    .B1(_04100_),
    .C1(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__nor2_1 _09939_ (.A(_04051_),
    .B(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hd__a221o_1 _09940_ (.A1(\irq_mask[15] ),
    .A2(_04021_),
    .B1(\timer[15] ),
    .B2(_04023_),
    .C1(_04188_),
    .X(_04661_));
 sky130_fd_sc_hd__a22o_1 _09941_ (.A1(\count_instr[47] ),
    .A2(_04015_),
    .B1(_04017_),
    .B2(\count_cycle[47] ),
    .X(_04662_));
 sky130_fd_sc_hd__a221o_1 _09942_ (.A1(\count_instr[15] ),
    .A2(_04145_),
    .B1(\count_cycle[15] ),
    .B2(_03253_),
    .C1(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__o22a_1 _09943_ (.A1(_04660_),
    .A2(_04661_),
    .B1(_04663_),
    .B2(_04268_),
    .X(_04664_));
 sky130_fd_sc_hd__or2_1 _09944_ (.A(latched_is_lb),
    .B(latched_is_lh),
    .X(_04665_));
 sky130_fd_sc_hd__buf_2 _09945_ (.A(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__buf_2 _09946_ (.A(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__nor2_4 _09947_ (.A(\mem_wordsize[2] ),
    .B(\mem_wordsize[1] ),
    .Y(_04668_));
 sky130_fd_sc_hd__a21o_1 _09948_ (.A1(_03297_),
    .A2(_04361_),
    .B1(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__o21a_1 _09949_ (.A1(net39),
    .A2(_04034_),
    .B1(_04669_),
    .X(_04670_));
 sky130_fd_sc_hd__inv_2 _09950_ (.A(_04666_),
    .Y(_04671_));
 sky130_fd_sc_hd__a211o_1 _09951_ (.A1(latched_is_lh),
    .A2(_04670_),
    .B1(_04671_),
    .C1(_04420_),
    .X(_04672_));
 sky130_fd_sc_hd__and2_2 _09952_ (.A(\cpu_state[6] ),
    .B(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__o21a_1 _09953_ (.A1(_04667_),
    .A2(_04670_),
    .B1(_04673_),
    .X(_04674_));
 sky130_fd_sc_hd__a221o_1 _09954_ (.A1(_03638_),
    .A2(_04642_),
    .B1(_04664_),
    .B2(_03302_),
    .C1(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__a221o_1 _09955_ (.A1(\irq_pending[15] ),
    .A2(_04049_),
    .B1(_04641_),
    .B2(_03385_),
    .C1(_04675_),
    .X(_08375_));
 sky130_fd_sc_hd__or2_1 _09956_ (.A(_04607_),
    .B(_04639_),
    .X(_04676_));
 sky130_fd_sc_hd__or2b_1 _09957_ (.A(_04535_),
    .B_N(_04598_),
    .X(_04677_));
 sky130_fd_sc_hd__a21o_1 _09958_ (.A1(_04597_),
    .A2(_04677_),
    .B1(_04676_),
    .X(_04678_));
 sky130_fd_sc_hd__o211a_1 _09959_ (.A1(\reg_pc[15] ),
    .A2(\decoded_imm[15] ),
    .B1(\decoded_imm[14] ),
    .C1(\reg_pc[14] ),
    .X(_04679_));
 sky130_fd_sc_hd__a21oi_1 _09960_ (.A1(\reg_pc[15] ),
    .A2(\decoded_imm[15] ),
    .B1(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__o311a_1 _09961_ (.A1(_04542_),
    .A2(_04599_),
    .A3(_04676_),
    .B1(_04678_),
    .C1(_04680_),
    .X(_04681_));
 sky130_fd_sc_hd__xnor2_1 _09962_ (.A(\reg_pc[16] ),
    .B(\decoded_imm[16] ),
    .Y(_04682_));
 sky130_fd_sc_hd__nor2_1 _09963_ (.A(_04681_),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__and2_1 _09964_ (.A(_04681_),
    .B(_04682_),
    .X(_04684_));
 sky130_fd_sc_hd__nor2_1 _09965_ (.A(_04683_),
    .B(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__mux4_1 _09966_ (.A0(\cpuregs.regs[28][16] ),
    .A1(\cpuregs.regs[29][16] ),
    .A2(\cpuregs.regs[30][16] ),
    .A3(\cpuregs.regs[31][16] ),
    .S0(_04579_),
    .S1(_04470_),
    .X(_04686_));
 sky130_fd_sc_hd__mux4_1 _09967_ (.A0(\cpuregs.regs[24][16] ),
    .A1(\cpuregs.regs[25][16] ),
    .A2(\cpuregs.regs[26][16] ),
    .A3(\cpuregs.regs[27][16] ),
    .S0(_04281_),
    .S1(_04470_),
    .X(_04687_));
 sky130_fd_sc_hd__mux2_1 _09968_ (.A0(_04686_),
    .A1(_04687_),
    .S(_04575_),
    .X(_04688_));
 sky130_fd_sc_hd__nand2_1 _09969_ (.A(_04054_),
    .B(_04688_),
    .Y(_04689_));
 sky130_fd_sc_hd__mux4_1 _09970_ (.A0(\cpuregs.regs[20][16] ),
    .A1(\cpuregs.regs[21][16] ),
    .A2(\cpuregs.regs[22][16] ),
    .A3(\cpuregs.regs[23][16] ),
    .S0(_04477_),
    .S1(_04478_),
    .X(_04690_));
 sky130_fd_sc_hd__mux4_1 _09971_ (.A0(\cpuregs.regs[16][16] ),
    .A1(\cpuregs.regs[17][16] ),
    .A2(\cpuregs.regs[18][16] ),
    .A3(\cpuregs.regs[19][16] ),
    .S0(_04477_),
    .S1(_04478_),
    .X(_04691_));
 sky130_fd_sc_hd__mux2_1 _09972_ (.A0(_04690_),
    .A1(_04691_),
    .S(_04121_),
    .X(_04692_));
 sky130_fd_sc_hd__a21oi_1 _09973_ (.A1(_04070_),
    .A2(_04692_),
    .B1(_04082_),
    .Y(_04693_));
 sky130_fd_sc_hd__mux4_1 _09974_ (.A0(\cpuregs.regs[8][16] ),
    .A1(\cpuregs.regs[9][16] ),
    .A2(\cpuregs.regs[10][16] ),
    .A3(\cpuregs.regs[11][16] ),
    .S0(_04057_),
    .S1(_04060_),
    .X(_04694_));
 sky130_fd_sc_hd__mux4_1 _09975_ (.A0(\cpuregs.regs[12][16] ),
    .A1(\cpuregs.regs[13][16] ),
    .A2(\cpuregs.regs[14][16] ),
    .A3(\cpuregs.regs[15][16] ),
    .S0(_04232_),
    .S1(_04233_),
    .X(_04695_));
 sky130_fd_sc_hd__mux2_1 _09976_ (.A0(_04694_),
    .A1(_04695_),
    .S(_04369_),
    .X(_04696_));
 sky130_fd_sc_hd__mux4_1 _09977_ (.A0(\cpuregs.regs[4][16] ),
    .A1(\cpuregs.regs[5][16] ),
    .A2(\cpuregs.regs[6][16] ),
    .A3(\cpuregs.regs[7][16] ),
    .S0(_04487_),
    .S1(_04469_),
    .X(_04697_));
 sky130_fd_sc_hd__mux4_1 _09978_ (.A0(\cpuregs.regs[0][16] ),
    .A1(\cpuregs.regs[1][16] ),
    .A2(\cpuregs.regs[2][16] ),
    .A3(\cpuregs.regs[3][16] ),
    .S0(_04487_),
    .S1(_04469_),
    .X(_04698_));
 sky130_fd_sc_hd__mux2_1 _09979_ (.A0(_04697_),
    .A1(_04698_),
    .S(_04320_),
    .X(_04699_));
 sky130_fd_sc_hd__a21o_1 _09980_ (.A1(_04069_),
    .A2(_04699_),
    .B1(_04095_),
    .X(_04700_));
 sky130_fd_sc_hd__a21oi_1 _09981_ (.A1(_04231_),
    .A2(_04696_),
    .B1(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__a211o_4 _09982_ (.A1(_04689_),
    .A2(_04693_),
    .B1(_04100_),
    .C1(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__nor2_1 _09983_ (.A(_04051_),
    .B(_04702_),
    .Y(_04703_));
 sky130_fd_sc_hd__a221o_1 _09984_ (.A1(\irq_mask[16] ),
    .A2(_04022_),
    .B1(\timer[16] ),
    .B2(_04024_),
    .C1(_04027_),
    .X(_04704_));
 sky130_fd_sc_hd__a22o_1 _09985_ (.A1(\count_instr[16] ),
    .A2(_04145_),
    .B1(_04105_),
    .B2(\count_cycle[48] ),
    .X(_04705_));
 sky130_fd_sc_hd__a221o_1 _09986_ (.A1(\count_instr[48] ),
    .A2(_04016_),
    .B1(\count_cycle[16] ),
    .B2(_04014_),
    .C1(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__o22a_1 _09987_ (.A1(_04703_),
    .A2(_04704_),
    .B1(_04706_),
    .B2(_04010_),
    .X(_04707_));
 sky130_fd_sc_hd__clkbuf_4 _09988_ (.A(net74),
    .X(_04708_));
 sky130_fd_sc_hd__nand2_1 _09989_ (.A(_03225_),
    .B(_04672_),
    .Y(_04709_));
 sky130_fd_sc_hd__clkbuf_4 _09990_ (.A(_04668_),
    .X(_04710_));
 sky130_fd_sc_hd__a21oi_1 _09991_ (.A1(net40),
    .A2(_04710_),
    .B1(_04667_),
    .Y(_04711_));
 sky130_fd_sc_hd__nor2_2 _09992_ (.A(_04709_),
    .B(_04711_),
    .Y(_04712_));
 sky130_fd_sc_hd__a221o_1 _09993_ (.A1(_03638_),
    .A2(_04708_),
    .B1(_04202_),
    .B2(\irq_pending[16] ),
    .C1(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__a221o_1 _09994_ (.A1(_03385_),
    .A2(_04685_),
    .B1(_04707_),
    .B2(_03303_),
    .C1(_04713_),
    .X(_08376_));
 sky130_fd_sc_hd__nand2_1 _09995_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .Y(_04714_));
 sky130_fd_sc_hd__or2_1 _09996_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .X(_04715_));
 sky130_fd_sc_hd__and2_1 _09997_ (.A(_04714_),
    .B(_04715_),
    .X(_04716_));
 sky130_fd_sc_hd__a21o_1 _09998_ (.A1(\reg_pc[16] ),
    .A2(\decoded_imm[16] ),
    .B1(_04683_),
    .X(_04717_));
 sky130_fd_sc_hd__nand2_1 _09999_ (.A(_04716_),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__or2_1 _10000_ (.A(_04716_),
    .B(_04717_),
    .X(_04719_));
 sky130_fd_sc_hd__and3_1 _10001_ (.A(_03384_),
    .B(_04718_),
    .C(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__mux4_1 _10002_ (.A0(\cpuregs.regs[20][17] ),
    .A1(\cpuregs.regs[21][17] ),
    .A2(\cpuregs.regs[22][17] ),
    .A3(\cpuregs.regs[23][17] ),
    .S0(_04472_),
    .S1(_04473_),
    .X(_04721_));
 sky130_fd_sc_hd__mux4_1 _10003_ (.A0(\cpuregs.regs[16][17] ),
    .A1(\cpuregs.regs[17][17] ),
    .A2(\cpuregs.regs[18][17] ),
    .A3(\cpuregs.regs[19][17] ),
    .S0(_04057_),
    .S1(_04060_),
    .X(_04722_));
 sky130_fd_sc_hd__mux2_1 _10004_ (.A0(_04721_),
    .A1(_04722_),
    .S(_04065_),
    .X(_04723_));
 sky130_fd_sc_hd__nand2_1 _10005_ (.A(_04483_),
    .B(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__mux4_1 _10006_ (.A0(\cpuregs.regs[28][17] ),
    .A1(\cpuregs.regs[29][17] ),
    .A2(\cpuregs.regs[30][17] ),
    .A3(\cpuregs.regs[31][17] ),
    .S0(_04072_),
    .S1(_04074_),
    .X(_04725_));
 sky130_fd_sc_hd__mux4_1 _10007_ (.A0(\cpuregs.regs[24][17] ),
    .A1(\cpuregs.regs[25][17] ),
    .A2(\cpuregs.regs[26][17] ),
    .A3(\cpuregs.regs[27][17] ),
    .S0(_04072_),
    .S1(_04074_),
    .X(_04726_));
 sky130_fd_sc_hd__mux2_1 _10008_ (.A0(_04725_),
    .A1(_04726_),
    .S(_04078_),
    .X(_04727_));
 sky130_fd_sc_hd__a21oi_1 _10009_ (.A1(_04231_),
    .A2(_04727_),
    .B1(_04082_),
    .Y(_04728_));
 sky130_fd_sc_hd__mux4_1 _10010_ (.A0(\cpuregs.regs[4][17] ),
    .A1(\cpuregs.regs[5][17] ),
    .A2(\cpuregs.regs[6][17] ),
    .A3(\cpuregs.regs[7][17] ),
    .S0(_04477_),
    .S1(_04478_),
    .X(_04729_));
 sky130_fd_sc_hd__mux4_1 _10011_ (.A0(\cpuregs.regs[0][17] ),
    .A1(\cpuregs.regs[1][17] ),
    .A2(\cpuregs.regs[2][17] ),
    .A3(\cpuregs.regs[3][17] ),
    .S0(_04477_),
    .S1(_04478_),
    .X(_04730_));
 sky130_fd_sc_hd__mux2_1 _10012_ (.A0(_04729_),
    .A1(_04730_),
    .S(_04121_),
    .X(_04731_));
 sky130_fd_sc_hd__mux4_1 _10013_ (.A0(\cpuregs.regs[12][17] ),
    .A1(\cpuregs.regs[13][17] ),
    .A2(\cpuregs.regs[14][17] ),
    .A3(\cpuregs.regs[15][17] ),
    .S0(_04280_),
    .S1(_04059_),
    .X(_04732_));
 sky130_fd_sc_hd__mux4_1 _10014_ (.A0(\cpuregs.regs[8][17] ),
    .A1(\cpuregs.regs[9][17] ),
    .A2(\cpuregs.regs[10][17] ),
    .A3(\cpuregs.regs[11][17] ),
    .S0(_04280_),
    .S1(_04059_),
    .X(_04733_));
 sky130_fd_sc_hd__mux2_1 _10015_ (.A0(_04732_),
    .A1(_04733_),
    .S(_04064_),
    .X(_04734_));
 sky130_fd_sc_hd__a21o_1 _10016_ (.A1(_04053_),
    .A2(_04734_),
    .B1(_04095_),
    .X(_04735_));
 sky130_fd_sc_hd__a21oi_1 _10017_ (.A1(_04070_),
    .A2(_04731_),
    .B1(_04735_),
    .Y(_04736_));
 sky130_fd_sc_hd__a211o_4 _10018_ (.A1(_04724_),
    .A2(_04728_),
    .B1(net300),
    .C1(_04736_),
    .X(_04737_));
 sky130_fd_sc_hd__inv_2 _10019_ (.A(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__a221o_1 _10020_ (.A1(\irq_mask[17] ),
    .A2(_04448_),
    .B1(\timer[17] ),
    .B2(_04187_),
    .C1(_04027_),
    .X(_04739_));
 sky130_fd_sc_hd__a21o_1 _10021_ (.A1(_04168_),
    .A2(_04738_),
    .B1(_04739_),
    .X(_04740_));
 sky130_fd_sc_hd__a22o_1 _10022_ (.A1(\count_instr[49] ),
    .A2(_04104_),
    .B1(_04011_),
    .B2(\count_instr[17] ),
    .X(_04741_));
 sky130_fd_sc_hd__a211o_1 _10023_ (.A1(_04018_),
    .A2(\count_cycle[49] ),
    .B1(_04009_),
    .C1(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__a21o_1 _10024_ (.A1(\count_cycle[17] ),
    .A2(_04014_),
    .B1(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__clkbuf_4 _10025_ (.A(net75),
    .X(_04744_));
 sky130_fd_sc_hd__clkbuf_4 _10026_ (.A(_04668_),
    .X(_04745_));
 sky130_fd_sc_hd__a21o_1 _10027_ (.A1(net41),
    .A2(_04745_),
    .B1(_04666_),
    .X(_04746_));
 sky130_fd_sc_hd__a221o_1 _10028_ (.A1(_03637_),
    .A2(_04744_),
    .B1(_04673_),
    .B2(_04746_),
    .C1(_04266_),
    .X(_04747_));
 sky130_fd_sc_hd__a31o_1 _10029_ (.A1(_04150_),
    .A2(_04740_),
    .A3(_04743_),
    .B1(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__o22a_1 _10030_ (.A1(\irq_pending[17] ),
    .A2(_04008_),
    .B1(_04720_),
    .B2(_04748_),
    .X(_08377_));
 sky130_fd_sc_hd__xnor2_1 _10031_ (.A(\reg_pc[18] ),
    .B(\decoded_imm[18] ),
    .Y(_04749_));
 sky130_fd_sc_hd__and3_1 _10032_ (.A(_04714_),
    .B(_04718_),
    .C(_04749_),
    .X(_04750_));
 sky130_fd_sc_hd__a21oi_1 _10033_ (.A1(_04714_),
    .A2(_04718_),
    .B1(_04749_),
    .Y(_04751_));
 sky130_fd_sc_hd__buf_2 _10034_ (.A(_04673_),
    .X(_04752_));
 sky130_fd_sc_hd__a21o_1 _10035_ (.A1(net42),
    .A2(_04710_),
    .B1(_04667_),
    .X(_04753_));
 sky130_fd_sc_hd__clkbuf_4 _10036_ (.A(net76),
    .X(_04754_));
 sky130_fd_sc_hd__a22o_1 _10037_ (.A1(_04046_),
    .A2(_04754_),
    .B1(_04202_),
    .B2(\irq_pending[18] ),
    .X(_04755_));
 sky130_fd_sc_hd__a22o_1 _10038_ (.A1(\count_instr[50] ),
    .A2(_04104_),
    .B1(_04105_),
    .B2(\count_cycle[50] ),
    .X(_04756_));
 sky130_fd_sc_hd__a221o_1 _10039_ (.A1(\count_instr[18] ),
    .A2(_04012_),
    .B1(\count_cycle[18] ),
    .B2(_04165_),
    .C1(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__buf_8 _10040_ (.A(_04232_),
    .X(_04758_));
 sky130_fd_sc_hd__buf_6 _10041_ (.A(_04233_),
    .X(_04759_));
 sky130_fd_sc_hd__mux4_1 _10042_ (.A0(\cpuregs.regs[16][18] ),
    .A1(\cpuregs.regs[17][18] ),
    .A2(\cpuregs.regs[18][18] ),
    .A3(\cpuregs.regs[19][18] ),
    .S0(_04758_),
    .S1(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__mux4_1 _10043_ (.A0(\cpuregs.regs[20][18] ),
    .A1(\cpuregs.regs[21][18] ),
    .A2(\cpuregs.regs[22][18] ),
    .A3(\cpuregs.regs[23][18] ),
    .S0(_04057_),
    .S1(_04060_),
    .X(_04761_));
 sky130_fd_sc_hd__or2_1 _10044_ (.A(_04575_),
    .B(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__o211a_1 _10045_ (.A1(_04430_),
    .A2(_04760_),
    .B1(_04762_),
    .C1(_04070_),
    .X(_04763_));
 sky130_fd_sc_hd__mux4_1 _10046_ (.A0(\cpuregs.regs[28][18] ),
    .A1(\cpuregs.regs[29][18] ),
    .A2(\cpuregs.regs[30][18] ),
    .A3(\cpuregs.regs[31][18] ),
    .S0(_04472_),
    .S1(_04473_),
    .X(_04764_));
 sky130_fd_sc_hd__mux4_1 _10047_ (.A0(\cpuregs.regs[24][18] ),
    .A1(\cpuregs.regs[25][18] ),
    .A2(\cpuregs.regs[26][18] ),
    .A3(\cpuregs.regs[27][18] ),
    .S0(_04472_),
    .S1(_04473_),
    .X(_04765_));
 sky130_fd_sc_hd__mux2_1 _10048_ (.A0(_04764_),
    .A1(_04765_),
    .S(_04065_),
    .X(_04766_));
 sky130_fd_sc_hd__a21o_1 _10049_ (.A1(_04231_),
    .A2(_04766_),
    .B1(_04082_),
    .X(_04767_));
 sky130_fd_sc_hd__mux4_1 _10050_ (.A0(\cpuregs.regs[0][18] ),
    .A1(\cpuregs.regs[1][18] ),
    .A2(\cpuregs.regs[2][18] ),
    .A3(\cpuregs.regs[3][18] ),
    .S0(_04057_),
    .S1(_04060_),
    .X(_04768_));
 sky130_fd_sc_hd__or2_1 _10051_ (.A(_04430_),
    .B(_04768_),
    .X(_04769_));
 sky130_fd_sc_hd__mux4_1 _10052_ (.A0(\cpuregs.regs[4][18] ),
    .A1(\cpuregs.regs[5][18] ),
    .A2(\cpuregs.regs[6][18] ),
    .A3(\cpuregs.regs[7][18] ),
    .S0(_04472_),
    .S1(_04473_),
    .X(_04770_));
 sky130_fd_sc_hd__o21a_1 _10053_ (.A1(_04321_),
    .A2(_04770_),
    .B1(_04069_),
    .X(_04771_));
 sky130_fd_sc_hd__mux4_1 _10054_ (.A0(\cpuregs.regs[12][18] ),
    .A1(\cpuregs.regs[13][18] ),
    .A2(\cpuregs.regs[14][18] ),
    .A3(\cpuregs.regs[15][18] ),
    .S0(_04232_),
    .S1(_04233_),
    .X(_04772_));
 sky130_fd_sc_hd__mux4_1 _10055_ (.A0(\cpuregs.regs[8][18] ),
    .A1(\cpuregs.regs[9][18] ),
    .A2(\cpuregs.regs[10][18] ),
    .A3(\cpuregs.regs[11][18] ),
    .S0(_04477_),
    .S1(_04478_),
    .X(_04773_));
 sky130_fd_sc_hd__mux2_1 _10056_ (.A0(_04772_),
    .A1(_04773_),
    .S(_04121_),
    .X(_04774_));
 sky130_fd_sc_hd__a221o_1 _10057_ (.A1(_04769_),
    .A2(_04771_),
    .B1(_04774_),
    .B2(_04231_),
    .C1(_04237_),
    .X(_04775_));
 sky130_fd_sc_hd__o211ai_4 _10058_ (.A1(_04763_),
    .A2(_04767_),
    .B1(_04133_),
    .C1(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__inv_2 _10059_ (.A(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__a221o_1 _10060_ (.A1(\irq_mask[18] ),
    .A2(_04021_),
    .B1(\timer[18] ),
    .B2(_04023_),
    .C1(_04026_),
    .X(_04778_));
 sky130_fd_sc_hd__a21o_1 _10061_ (.A1(_04271_),
    .A2(_04777_),
    .B1(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__o211a_1 _10062_ (.A1(_04268_),
    .A2(_04757_),
    .B1(_04779_),
    .C1(_03302_),
    .X(_04780_));
 sky130_fd_sc_hd__a211oi_1 _10063_ (.A1(_04752_),
    .A2(_04753_),
    .B1(_04755_),
    .C1(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__o31ai_1 _10064_ (.A1(_04156_),
    .A2(_04750_),
    .A3(_04751_),
    .B1(_04781_),
    .Y(_08378_));
 sky130_fd_sc_hd__nand2_1 _10065_ (.A(\reg_pc[19] ),
    .B(\decoded_imm[19] ),
    .Y(_04782_));
 sky130_fd_sc_hd__or2_1 _10066_ (.A(\reg_pc[19] ),
    .B(\decoded_imm[19] ),
    .X(_04783_));
 sky130_fd_sc_hd__nand2_1 _10067_ (.A(_04782_),
    .B(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__a21o_1 _10068_ (.A1(\reg_pc[18] ),
    .A2(\decoded_imm[18] ),
    .B1(_04751_),
    .X(_04785_));
 sky130_fd_sc_hd__xnor2_1 _10069_ (.A(_04784_),
    .B(_04785_),
    .Y(_04786_));
 sky130_fd_sc_hd__a22o_1 _10070_ (.A1(\count_instr[51] ),
    .A2(_04104_),
    .B1(_04011_),
    .B2(\count_instr[19] ),
    .X(_04787_));
 sky130_fd_sc_hd__a221o_1 _10071_ (.A1(_04018_),
    .A2(\count_cycle[51] ),
    .B1(_04013_),
    .B2(\count_cycle[19] ),
    .C1(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__mux4_1 _10072_ (.A0(\cpuregs.regs[20][19] ),
    .A1(\cpuregs.regs[21][19] ),
    .A2(\cpuregs.regs[22][19] ),
    .A3(\cpuregs.regs[23][19] ),
    .S0(_04512_),
    .S1(_04513_),
    .X(_04789_));
 sky130_fd_sc_hd__mux4_1 _10073_ (.A0(\cpuregs.regs[16][19] ),
    .A1(\cpuregs.regs[17][19] ),
    .A2(\cpuregs.regs[18][19] ),
    .A3(\cpuregs.regs[19][19] ),
    .S0(_04512_),
    .S1(_04513_),
    .X(_04790_));
 sky130_fd_sc_hd__mux2_1 _10074_ (.A0(_04789_),
    .A1(_04790_),
    .S(_04321_),
    .X(_04791_));
 sky130_fd_sc_hd__nand2_1 _10075_ (.A(_04289_),
    .B(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__mux4_1 _10076_ (.A0(\cpuregs.regs[28][19] ),
    .A1(\cpuregs.regs[29][19] ),
    .A2(\cpuregs.regs[30][19] ),
    .A3(\cpuregs.regs[31][19] ),
    .S0(_04579_),
    .S1(_04284_),
    .X(_04793_));
 sky130_fd_sc_hd__mux4_1 _10077_ (.A0(\cpuregs.regs[24][19] ),
    .A1(\cpuregs.regs[25][19] ),
    .A2(\cpuregs.regs[26][19] ),
    .A3(\cpuregs.regs[27][19] ),
    .S0(_04579_),
    .S1(_04284_),
    .X(_04794_));
 sky130_fd_sc_hd__mux2_1 _10078_ (.A0(_04793_),
    .A1(_04794_),
    .S(_04575_),
    .X(_04795_));
 sky130_fd_sc_hd__a21oi_1 _10079_ (.A1(_04054_),
    .A2(_04795_),
    .B1(_04225_),
    .Y(_04796_));
 sky130_fd_sc_hd__mux4_1 _10080_ (.A0(\cpuregs.regs[4][19] ),
    .A1(\cpuregs.regs[5][19] ),
    .A2(\cpuregs.regs[6][19] ),
    .A3(\cpuregs.regs[7][19] ),
    .S0(_04512_),
    .S1(_04513_),
    .X(_04797_));
 sky130_fd_sc_hd__mux4_1 _10081_ (.A0(\cpuregs.regs[0][19] ),
    .A1(\cpuregs.regs[1][19] ),
    .A2(\cpuregs.regs[2][19] ),
    .A3(\cpuregs.regs[3][19] ),
    .S0(_04512_),
    .S1(_04513_),
    .X(_04798_));
 sky130_fd_sc_hd__mux2_1 _10082_ (.A0(_04797_),
    .A1(_04798_),
    .S(_04575_),
    .X(_04799_));
 sky130_fd_sc_hd__mux4_1 _10083_ (.A0(\cpuregs.regs[12][19] ),
    .A1(\cpuregs.regs[13][19] ),
    .A2(\cpuregs.regs[14][19] ),
    .A3(\cpuregs.regs[15][19] ),
    .S0(_04273_),
    .S1(_04283_),
    .X(_04800_));
 sky130_fd_sc_hd__mux4_1 _10084_ (.A0(\cpuregs.regs[8][19] ),
    .A1(\cpuregs.regs[9][19] ),
    .A2(\cpuregs.regs[10][19] ),
    .A3(\cpuregs.regs[11][19] ),
    .S0(_04273_),
    .S1(_04283_),
    .X(_04801_));
 sky130_fd_sc_hd__mux2_1 _10085_ (.A0(_04800_),
    .A1(_04801_),
    .S(_04320_),
    .X(_04802_));
 sky130_fd_sc_hd__a21o_1 _10086_ (.A1(_04328_),
    .A2(_04802_),
    .B1(_04237_),
    .X(_04803_));
 sky130_fd_sc_hd__a21oi_1 _10087_ (.A1(_04483_),
    .A2(_04799_),
    .B1(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__a211o_4 _10088_ (.A1(_04792_),
    .A2(_04796_),
    .B1(_04100_),
    .C1(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__inv_2 _10089_ (.A(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__a221o_1 _10090_ (.A1(\irq_mask[19] ),
    .A2(_04021_),
    .B1(\timer[19] ),
    .B2(_04023_),
    .C1(_04026_),
    .X(_04807_));
 sky130_fd_sc_hd__a21o_1 _10091_ (.A1(_04271_),
    .A2(_04806_),
    .B1(_04807_),
    .X(_04808_));
 sky130_fd_sc_hd__o211a_1 _10092_ (.A1(_04268_),
    .A2(_04788_),
    .B1(_04808_),
    .C1(_03302_),
    .X(_04809_));
 sky130_fd_sc_hd__clkbuf_4 _10093_ (.A(net77),
    .X(_04810_));
 sky130_fd_sc_hd__buf_2 _10094_ (.A(_04668_),
    .X(_04811_));
 sky130_fd_sc_hd__a21o_1 _10095_ (.A1(net43),
    .A2(_04811_),
    .B1(_04667_),
    .X(_04812_));
 sky130_fd_sc_hd__a221o_1 _10096_ (.A1(_04046_),
    .A2(_04810_),
    .B1(_04752_),
    .B2(_04812_),
    .C1(_04202_),
    .X(_04813_));
 sky130_fd_sc_hd__o22a_1 _10097_ (.A1(\irq_pending[19] ),
    .A2(_04007_),
    .B1(_04809_),
    .B2(_04813_),
    .X(_04814_));
 sky130_fd_sc_hd__a21o_1 _10098_ (.A1(_04391_),
    .A2(_04786_),
    .B1(_04814_),
    .X(_08379_));
 sky130_fd_sc_hd__nor2_1 _10099_ (.A(_04749_),
    .B(_04784_),
    .Y(_04815_));
 sky130_fd_sc_hd__and2_1 _10100_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .X(_04816_));
 sky130_fd_sc_hd__a31o_1 _10101_ (.A1(\reg_pc[16] ),
    .A2(\decoded_imm[16] ),
    .A3(_04715_),
    .B1(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__and3_1 _10102_ (.A(\reg_pc[18] ),
    .B(\decoded_imm[18] ),
    .C(_04783_),
    .X(_04818_));
 sky130_fd_sc_hd__a221o_1 _10103_ (.A1(\reg_pc[19] ),
    .A2(\decoded_imm[19] ),
    .B1(_04815_),
    .B2(_04817_),
    .C1(_04818_),
    .X(_04819_));
 sky130_fd_sc_hd__a31oi_1 _10104_ (.A1(_04683_),
    .A2(_04716_),
    .A3(_04815_),
    .B1(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__nand2_1 _10105_ (.A(\reg_pc[20] ),
    .B(\decoded_imm[20] ),
    .Y(_04821_));
 sky130_fd_sc_hd__or2_1 _10106_ (.A(\reg_pc[20] ),
    .B(\decoded_imm[20] ),
    .X(_04822_));
 sky130_fd_sc_hd__nand2_1 _10107_ (.A(_04821_),
    .B(_04822_),
    .Y(_04823_));
 sky130_fd_sc_hd__or2_1 _10108_ (.A(_04820_),
    .B(_04823_),
    .X(_04824_));
 sky130_fd_sc_hd__nand2_1 _10109_ (.A(_04820_),
    .B(_04823_),
    .Y(_04825_));
 sky130_fd_sc_hd__mux4_1 _10110_ (.A0(\cpuregs.regs[12][20] ),
    .A1(\cpuregs.regs[13][20] ),
    .A2(\cpuregs.regs[14][20] ),
    .A3(\cpuregs.regs[15][20] ),
    .S0(_04275_),
    .S1(_04278_),
    .X(_04826_));
 sky130_fd_sc_hd__mux4_1 _10111_ (.A0(\cpuregs.regs[8][20] ),
    .A1(\cpuregs.regs[9][20] ),
    .A2(\cpuregs.regs[10][20] ),
    .A3(\cpuregs.regs[11][20] ),
    .S0(_04275_),
    .S1(_04278_),
    .X(_04827_));
 sky130_fd_sc_hd__mux2_1 _10112_ (.A0(_04826_),
    .A1(_04827_),
    .S(_04287_),
    .X(_04828_));
 sky130_fd_sc_hd__nand2_1 _10113_ (.A(_04272_),
    .B(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__mux4_1 _10114_ (.A0(\cpuregs.regs[4][20] ),
    .A1(\cpuregs.regs[5][20] ),
    .A2(\cpuregs.regs[6][20] ),
    .A3(\cpuregs.regs[7][20] ),
    .S0(_04275_),
    .S1(_04278_),
    .X(_04830_));
 sky130_fd_sc_hd__mux4_1 _10115_ (.A0(\cpuregs.regs[0][20] ),
    .A1(\cpuregs.regs[1][20] ),
    .A2(\cpuregs.regs[2][20] ),
    .A3(\cpuregs.regs[3][20] ),
    .S0(_04275_),
    .S1(_04278_),
    .X(_04831_));
 sky130_fd_sc_hd__mux2_1 _10116_ (.A0(_04830_),
    .A1(_04831_),
    .S(_04287_),
    .X(_04832_));
 sky130_fd_sc_hd__a21oi_2 _10117_ (.A1(_04215_),
    .A2(_04832_),
    .B1(_04296_),
    .Y(_04833_));
 sky130_fd_sc_hd__mux4_1 _10118_ (.A0(\cpuregs.regs[24][20] ),
    .A1(\cpuregs.regs[25][20] ),
    .A2(\cpuregs.regs[26][20] ),
    .A3(\cpuregs.regs[27][20] ),
    .S0(_04275_),
    .S1(_04278_),
    .X(_04834_));
 sky130_fd_sc_hd__mux4_1 _10119_ (.A0(\cpuregs.regs[28][20] ),
    .A1(\cpuregs.regs[29][20] ),
    .A2(\cpuregs.regs[30][20] ),
    .A3(\cpuregs.regs[31][20] ),
    .S0(_04275_),
    .S1(_04278_),
    .X(_04835_));
 sky130_fd_sc_hd__mux2_1 _10120_ (.A0(_04834_),
    .A1(_04835_),
    .S(_04430_),
    .X(_04836_));
 sky130_fd_sc_hd__mux4_1 _10121_ (.A0(\cpuregs.regs[20][20] ),
    .A1(\cpuregs.regs[21][20] ),
    .A2(\cpuregs.regs[22][20] ),
    .A3(\cpuregs.regs[23][20] ),
    .S0(_04282_),
    .S1(_04285_),
    .X(_04837_));
 sky130_fd_sc_hd__mux4_1 _10122_ (.A0(\cpuregs.regs[16][20] ),
    .A1(\cpuregs.regs[17][20] ),
    .A2(\cpuregs.regs[18][20] ),
    .A3(\cpuregs.regs[19][20] ),
    .S0(_04282_),
    .S1(_04285_),
    .X(_04838_));
 sky130_fd_sc_hd__mux2_1 _10123_ (.A0(_04837_),
    .A1(_04838_),
    .S(_04287_),
    .X(_04839_));
 sky130_fd_sc_hd__a21o_1 _10124_ (.A1(_04215_),
    .A2(_04839_),
    .B1(_04225_),
    .X(_04840_));
 sky130_fd_sc_hd__a21oi_1 _10125_ (.A1(_04272_),
    .A2(_04836_),
    .B1(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__a211oi_4 _10126_ (.A1(_04829_),
    .A2(_04833_),
    .B1(_04841_),
    .C1(_04227_),
    .Y(_04842_));
 sky130_fd_sc_hd__a221o_1 _10127_ (.A1(\irq_mask[20] ),
    .A2(_04448_),
    .B1(\timer[20] ),
    .B2(_04024_),
    .C1(_04027_),
    .X(_04843_));
 sky130_fd_sc_hd__a21o_1 _10128_ (.A1(_04168_),
    .A2(_04842_),
    .B1(_04843_),
    .X(_04844_));
 sky130_fd_sc_hd__a22o_1 _10129_ (.A1(\count_instr[52] ),
    .A2(_04104_),
    .B1(_04105_),
    .B2(\count_cycle[52] ),
    .X(_04845_));
 sky130_fd_sc_hd__a211o_1 _10130_ (.A1(\count_instr[20] ),
    .A2(_04012_),
    .B1(_04009_),
    .C1(_04845_),
    .X(_04846_));
 sky130_fd_sc_hd__a21o_1 _10131_ (.A1(\count_cycle[20] ),
    .A2(_04014_),
    .B1(_04846_),
    .X(_04847_));
 sky130_fd_sc_hd__clkbuf_4 _10132_ (.A(net79),
    .X(_04848_));
 sky130_fd_sc_hd__a21oi_1 _10133_ (.A1(net45),
    .A2(_04745_),
    .B1(_04666_),
    .Y(_04849_));
 sky130_fd_sc_hd__nor2_2 _10134_ (.A(_04709_),
    .B(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__a221o_1 _10135_ (.A1(_03637_),
    .A2(_04848_),
    .B1(_04048_),
    .B2(\irq_pending[20] ),
    .C1(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__a31o_1 _10136_ (.A1(_03303_),
    .A2(_04844_),
    .A3(_04847_),
    .B1(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__a31o_1 _10137_ (.A1(_04391_),
    .A2(_04824_),
    .A3(_04825_),
    .B1(_04852_),
    .X(_08381_));
 sky130_fd_sc_hd__a22o_1 _10138_ (.A1(\count_instr[53] ),
    .A2(_04016_),
    .B1(_04012_),
    .B2(\count_instr[21] ),
    .X(_04853_));
 sky130_fd_sc_hd__a221o_1 _10139_ (.A1(_04018_),
    .A2(\count_cycle[53] ),
    .B1(_04014_),
    .B2(\count_cycle[21] ),
    .C1(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__mux4_1 _10140_ (.A0(\cpuregs.regs[8][21] ),
    .A1(\cpuregs.regs[9][21] ),
    .A2(\cpuregs.regs[10][21] ),
    .A3(\cpuregs.regs[11][21] ),
    .S0(_04282_),
    .S1(_04285_),
    .X(_04855_));
 sky130_fd_sc_hd__mux4_1 _10141_ (.A0(\cpuregs.regs[12][21] ),
    .A1(\cpuregs.regs[13][21] ),
    .A2(\cpuregs.regs[14][21] ),
    .A3(\cpuregs.regs[15][21] ),
    .S0(_04282_),
    .S1(_04285_),
    .X(_04856_));
 sky130_fd_sc_hd__mux2_1 _10142_ (.A0(_04855_),
    .A1(_04856_),
    .S(_04430_),
    .X(_04857_));
 sky130_fd_sc_hd__nand2_1 _10143_ (.A(_04272_),
    .B(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__mux4_1 _10144_ (.A0(\cpuregs.regs[4][21] ),
    .A1(\cpuregs.regs[5][21] ),
    .A2(\cpuregs.regs[6][21] ),
    .A3(\cpuregs.regs[7][21] ),
    .S0(_04758_),
    .S1(_04759_),
    .X(_04859_));
 sky130_fd_sc_hd__mux4_1 _10145_ (.A0(\cpuregs.regs[0][21] ),
    .A1(\cpuregs.regs[1][21] ),
    .A2(\cpuregs.regs[2][21] ),
    .A3(\cpuregs.regs[3][21] ),
    .S0(_04758_),
    .S1(_04759_),
    .X(_04860_));
 sky130_fd_sc_hd__mux2_1 _10146_ (.A0(_04859_),
    .A1(_04860_),
    .S(_04211_),
    .X(_04861_));
 sky130_fd_sc_hd__a21oi_1 _10147_ (.A1(_04215_),
    .A2(_04861_),
    .B1(_04296_),
    .Y(_04862_));
 sky130_fd_sc_hd__mux4_1 _10148_ (.A0(\cpuregs.regs[28][21] ),
    .A1(\cpuregs.regs[29][21] ),
    .A2(\cpuregs.regs[30][21] ),
    .A3(\cpuregs.regs[31][21] ),
    .S0(_04758_),
    .S1(_04759_),
    .X(_04863_));
 sky130_fd_sc_hd__mux4_1 _10149_ (.A0(\cpuregs.regs[24][21] ),
    .A1(\cpuregs.regs[25][21] ),
    .A2(\cpuregs.regs[26][21] ),
    .A3(\cpuregs.regs[27][21] ),
    .S0(_04758_),
    .S1(_04759_),
    .X(_04864_));
 sky130_fd_sc_hd__mux2_1 _10150_ (.A0(_04863_),
    .A1(_04864_),
    .S(_04287_),
    .X(_04865_));
 sky130_fd_sc_hd__mux4_1 _10151_ (.A0(\cpuregs.regs[20][21] ),
    .A1(\cpuregs.regs[21][21] ),
    .A2(\cpuregs.regs[22][21] ),
    .A3(\cpuregs.regs[23][21] ),
    .S0(_04579_),
    .S1(_04284_),
    .X(_04866_));
 sky130_fd_sc_hd__mux4_1 _10152_ (.A0(\cpuregs.regs[16][21] ),
    .A1(\cpuregs.regs[17][21] ),
    .A2(\cpuregs.regs[18][21] ),
    .A3(\cpuregs.regs[19][21] ),
    .S0(_04579_),
    .S1(_04284_),
    .X(_04867_));
 sky130_fd_sc_hd__mux2_1 _10153_ (.A0(_04866_),
    .A1(_04867_),
    .S(_04575_),
    .X(_04868_));
 sky130_fd_sc_hd__a21o_1 _10154_ (.A1(_04483_),
    .A2(_04868_),
    .B1(_04082_),
    .X(_04869_));
 sky130_fd_sc_hd__a21oi_1 _10155_ (.A1(_04272_),
    .A2(_04865_),
    .B1(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__a211oi_4 _10156_ (.A1(_04858_),
    .A2(_04862_),
    .B1(_04870_),
    .C1(_04227_),
    .Y(_04871_));
 sky130_fd_sc_hd__a221o_1 _10157_ (.A1(\irq_mask[21] ),
    .A2(_04448_),
    .B1(\timer[21] ),
    .B2(_04024_),
    .C1(_04027_),
    .X(_04872_));
 sky130_fd_sc_hd__a21o_1 _10158_ (.A1(_04168_),
    .A2(_04871_),
    .B1(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__o211a_1 _10159_ (.A1(_04010_),
    .A2(_04854_),
    .B1(_04873_),
    .C1(_04150_),
    .X(_04874_));
 sky130_fd_sc_hd__nand2_1 _10160_ (.A(\reg_pc[21] ),
    .B(\decoded_imm[21] ),
    .Y(_04875_));
 sky130_fd_sc_hd__or2_1 _10161_ (.A(\reg_pc[21] ),
    .B(\decoded_imm[21] ),
    .X(_04876_));
 sky130_fd_sc_hd__nand2_1 _10162_ (.A(_04875_),
    .B(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__a21o_1 _10163_ (.A1(_04821_),
    .A2(_04824_),
    .B1(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__nand3_1 _10164_ (.A(_04821_),
    .B(_04824_),
    .C(_04877_),
    .Y(_04879_));
 sky130_fd_sc_hd__buf_4 _10165_ (.A(net80),
    .X(_04880_));
 sky130_fd_sc_hd__a21o_1 _10166_ (.A1(net46),
    .A2(_04745_),
    .B1(_04666_),
    .X(_04881_));
 sky130_fd_sc_hd__a221o_1 _10167_ (.A1(_03637_),
    .A2(_04880_),
    .B1(_04673_),
    .B2(_04881_),
    .C1(_04048_),
    .X(_04882_));
 sky130_fd_sc_hd__a31o_1 _10168_ (.A1(_03384_),
    .A2(_04878_),
    .A3(_04879_),
    .B1(_04882_),
    .X(_04883_));
 sky130_fd_sc_hd__o22a_1 _10169_ (.A1(\irq_pending[21] ),
    .A2(_04008_),
    .B1(_04874_),
    .B2(_04883_),
    .X(_08382_));
 sky130_fd_sc_hd__nand2_1 _10170_ (.A(\reg_pc[22] ),
    .B(\decoded_imm[22] ),
    .Y(_04884_));
 sky130_fd_sc_hd__or2_1 _10171_ (.A(\reg_pc[22] ),
    .B(\decoded_imm[22] ),
    .X(_04885_));
 sky130_fd_sc_hd__nand2_1 _10172_ (.A(_04884_),
    .B(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__nand3_1 _10173_ (.A(_04875_),
    .B(_04878_),
    .C(_04886_),
    .Y(_04887_));
 sky130_fd_sc_hd__a21o_1 _10174_ (.A1(_04875_),
    .A2(_04878_),
    .B1(_04886_),
    .X(_04888_));
 sky130_fd_sc_hd__a22o_1 _10175_ (.A1(\count_instr[54] ),
    .A2(_04015_),
    .B1(_04017_),
    .B2(\count_cycle[54] ),
    .X(_04889_));
 sky130_fd_sc_hd__a221o_1 _10176_ (.A1(\count_instr[22] ),
    .A2(_04145_),
    .B1(\count_cycle[22] ),
    .B2(_04013_),
    .C1(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__mux4_1 _10177_ (.A0(\cpuregs.regs[20][22] ),
    .A1(\cpuregs.regs[21][22] ),
    .A2(\cpuregs.regs[22][22] ),
    .A3(\cpuregs.regs[23][22] ),
    .S0(_04281_),
    .S1(_04470_),
    .X(_04891_));
 sky130_fd_sc_hd__mux4_1 _10178_ (.A0(\cpuregs.regs[16][22] ),
    .A1(\cpuregs.regs[17][22] ),
    .A2(\cpuregs.regs[18][22] ),
    .A3(\cpuregs.regs[19][22] ),
    .S0(_04281_),
    .S1(_04470_),
    .X(_04892_));
 sky130_fd_sc_hd__mux2_1 _10179_ (.A0(_04891_),
    .A1(_04892_),
    .S(_04065_),
    .X(_04893_));
 sky130_fd_sc_hd__nand2_1 _10180_ (.A(_04483_),
    .B(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__mux4_1 _10181_ (.A0(\cpuregs.regs[28][22] ),
    .A1(\cpuregs.regs[29][22] ),
    .A2(\cpuregs.regs[30][22] ),
    .A3(\cpuregs.regs[31][22] ),
    .S0(_04281_),
    .S1(_04470_),
    .X(_04895_));
 sky130_fd_sc_hd__mux4_1 _10182_ (.A0(\cpuregs.regs[24][22] ),
    .A1(\cpuregs.regs[25][22] ),
    .A2(\cpuregs.regs[26][22] ),
    .A3(\cpuregs.regs[27][22] ),
    .S0(_04281_),
    .S1(_04470_),
    .X(_04896_));
 sky130_fd_sc_hd__mux2_1 _10183_ (.A0(_04895_),
    .A1(_04896_),
    .S(_04065_),
    .X(_04897_));
 sky130_fd_sc_hd__nand2_1 _10184_ (.A(_04054_),
    .B(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__mux4_1 _10185_ (.A0(\cpuregs.regs[0][22] ),
    .A1(\cpuregs.regs[1][22] ),
    .A2(\cpuregs.regs[2][22] ),
    .A3(\cpuregs.regs[3][22] ),
    .S0(_04056_),
    .S1(_04091_),
    .X(_04899_));
 sky130_fd_sc_hd__or2_1 _10186_ (.A(_04369_),
    .B(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__mux4_1 _10187_ (.A0(\cpuregs.regs[4][22] ),
    .A1(\cpuregs.regs[5][22] ),
    .A2(\cpuregs.regs[6][22] ),
    .A3(\cpuregs.regs[7][22] ),
    .S0(_04280_),
    .S1(_04059_),
    .X(_04901_));
 sky130_fd_sc_hd__o21a_1 _10188_ (.A1(_04320_),
    .A2(_04901_),
    .B1(_04068_),
    .X(_04902_));
 sky130_fd_sc_hd__mux4_1 _10189_ (.A0(\cpuregs.regs[12][22] ),
    .A1(\cpuregs.regs[13][22] ),
    .A2(\cpuregs.regs[14][22] ),
    .A3(\cpuregs.regs[15][22] ),
    .S0(_04084_),
    .S1(_04086_),
    .X(_04903_));
 sky130_fd_sc_hd__mux4_1 _10190_ (.A0(\cpuregs.regs[8][22] ),
    .A1(\cpuregs.regs[9][22] ),
    .A2(\cpuregs.regs[10][22] ),
    .A3(\cpuregs.regs[11][22] ),
    .S0(_04084_),
    .S1(_04086_),
    .X(_04904_));
 sky130_fd_sc_hd__mux2_1 _10191_ (.A0(_04903_),
    .A1(_04904_),
    .S(_04064_),
    .X(_04905_));
 sky130_fd_sc_hd__a221o_1 _10192_ (.A1(_04900_),
    .A2(_04902_),
    .B1(_04905_),
    .B2(_04052_),
    .C1(_04095_),
    .X(_04906_));
 sky130_fd_sc_hd__nand2_1 _10193_ (.A(_04133_),
    .B(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__a31o_2 _10194_ (.A1(_04296_),
    .A2(_04894_),
    .A3(_04898_),
    .B1(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__inv_2 _10195_ (.A(_04908_),
    .Y(_04909_));
 sky130_fd_sc_hd__a221o_1 _10196_ (.A1(\irq_mask[22] ),
    .A2(_04308_),
    .B1(\timer[22] ),
    .B2(instr_timer),
    .C1(_04026_),
    .X(_04910_));
 sky130_fd_sc_hd__a21o_1 _10197_ (.A1(_04271_),
    .A2(_04909_),
    .B1(_04910_),
    .X(_04911_));
 sky130_fd_sc_hd__o211a_1 _10198_ (.A1(_04268_),
    .A2(_04890_),
    .B1(_04911_),
    .C1(_04149_),
    .X(_04912_));
 sky130_fd_sc_hd__buf_4 _10199_ (.A(net81),
    .X(_04913_));
 sky130_fd_sc_hd__a21o_1 _10200_ (.A1(net47),
    .A2(_04745_),
    .B1(_04666_),
    .X(_04914_));
 sky130_fd_sc_hd__a221o_1 _10201_ (.A1(_03637_),
    .A2(_04913_),
    .B1(_04673_),
    .B2(_04914_),
    .C1(_04266_),
    .X(_04915_));
 sky130_fd_sc_hd__o22a_1 _10202_ (.A1(\irq_pending[22] ),
    .A2(_04006_),
    .B1(_04912_),
    .B2(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__a31o_1 _10203_ (.A1(_04391_),
    .A2(_04887_),
    .A3(_04888_),
    .B1(_04916_),
    .X(_08383_));
 sky130_fd_sc_hd__nand2_1 _10204_ (.A(\reg_pc[23] ),
    .B(\decoded_imm[23] ),
    .Y(_04917_));
 sky130_fd_sc_hd__or2_1 _10205_ (.A(\reg_pc[23] ),
    .B(\decoded_imm[23] ),
    .X(_04918_));
 sky130_fd_sc_hd__nand2_1 _10206_ (.A(_04917_),
    .B(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__a21o_1 _10207_ (.A1(_04884_),
    .A2(_04888_),
    .B1(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__nand3_1 _10208_ (.A(_04884_),
    .B(_04888_),
    .C(_04919_),
    .Y(_04921_));
 sky130_fd_sc_hd__a22o_1 _10209_ (.A1(\count_instr[55] ),
    .A2(_04015_),
    .B1(_04011_),
    .B2(\count_instr[23] ),
    .X(_04922_));
 sky130_fd_sc_hd__a221o_1 _10210_ (.A1(_04105_),
    .A2(\count_cycle[55] ),
    .B1(_04013_),
    .B2(\count_cycle[23] ),
    .C1(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__mux4_1 _10211_ (.A0(\cpuregs.regs[12][23] ),
    .A1(\cpuregs.regs[13][23] ),
    .A2(\cpuregs.regs[14][23] ),
    .A3(\cpuregs.regs[15][23] ),
    .S0(_04512_),
    .S1(_04513_),
    .X(_04924_));
 sky130_fd_sc_hd__mux4_1 _10212_ (.A0(\cpuregs.regs[8][23] ),
    .A1(\cpuregs.regs[9][23] ),
    .A2(\cpuregs.regs[10][23] ),
    .A3(\cpuregs.regs[11][23] ),
    .S0(_04512_),
    .S1(_04513_),
    .X(_04925_));
 sky130_fd_sc_hd__mux2_1 _10213_ (.A0(_04924_),
    .A1(_04925_),
    .S(_04575_),
    .X(_04926_));
 sky130_fd_sc_hd__nand2_1 _10214_ (.A(_04206_),
    .B(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__mux4_1 _10215_ (.A0(\cpuregs.regs[4][23] ),
    .A1(\cpuregs.regs[5][23] ),
    .A2(\cpuregs.regs[6][23] ),
    .A3(\cpuregs.regs[7][23] ),
    .S0(_04472_),
    .S1(_04473_),
    .X(_04928_));
 sky130_fd_sc_hd__mux4_1 _10216_ (.A0(\cpuregs.regs[0][23] ),
    .A1(\cpuregs.regs[1][23] ),
    .A2(\cpuregs.regs[2][23] ),
    .A3(\cpuregs.regs[3][23] ),
    .S0(_04472_),
    .S1(_04473_),
    .X(_04929_));
 sky130_fd_sc_hd__mux2_1 _10217_ (.A0(_04928_),
    .A1(_04929_),
    .S(_04065_),
    .X(_04930_));
 sky130_fd_sc_hd__a21oi_1 _10218_ (.A1(_04483_),
    .A2(_04930_),
    .B1(_04296_),
    .Y(_04931_));
 sky130_fd_sc_hd__mux4_1 _10219_ (.A0(\cpuregs.regs[24][23] ),
    .A1(\cpuregs.regs[25][23] ),
    .A2(\cpuregs.regs[26][23] ),
    .A3(\cpuregs.regs[27][23] ),
    .S0(_04281_),
    .S1(_04470_),
    .X(_04932_));
 sky130_fd_sc_hd__mux4_1 _10220_ (.A0(\cpuregs.regs[28][23] ),
    .A1(\cpuregs.regs[29][23] ),
    .A2(\cpuregs.regs[30][23] ),
    .A3(\cpuregs.regs[31][23] ),
    .S0(_04281_),
    .S1(_04470_),
    .X(_04933_));
 sky130_fd_sc_hd__mux2_1 _10221_ (.A0(_04932_),
    .A1(_04933_),
    .S(_04430_),
    .X(_04934_));
 sky130_fd_sc_hd__mux4_1 _10222_ (.A0(\cpuregs.regs[20][23] ),
    .A1(\cpuregs.regs[21][23] ),
    .A2(\cpuregs.regs[22][23] ),
    .A3(\cpuregs.regs[23][23] ),
    .S0(_04280_),
    .S1(_04059_),
    .X(_04935_));
 sky130_fd_sc_hd__mux4_1 _10223_ (.A0(\cpuregs.regs[16][23] ),
    .A1(\cpuregs.regs[17][23] ),
    .A2(\cpuregs.regs[18][23] ),
    .A3(\cpuregs.regs[19][23] ),
    .S0(_04280_),
    .S1(_04059_),
    .X(_04936_));
 sky130_fd_sc_hd__mux2_1 _10224_ (.A0(_04935_),
    .A1(_04936_),
    .S(_04064_),
    .X(_04937_));
 sky130_fd_sc_hd__a21oi_1 _10225_ (.A1(_04069_),
    .A2(_04937_),
    .B1(_04081_),
    .Y(_04938_));
 sky130_fd_sc_hd__a21boi_1 _10226_ (.A1(_04054_),
    .A2(_04934_),
    .B1_N(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__a211o_2 _10227_ (.A1(_04927_),
    .A2(_04931_),
    .B1(_04939_),
    .C1(_04100_),
    .X(_04940_));
 sky130_fd_sc_hd__inv_2 _10228_ (.A(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__a221o_1 _10229_ (.A1(\irq_mask[23] ),
    .A2(_04308_),
    .B1(\timer[23] ),
    .B2(instr_timer),
    .C1(_04026_),
    .X(_04942_));
 sky130_fd_sc_hd__a21o_1 _10230_ (.A1(_04271_),
    .A2(_04941_),
    .B1(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__o211a_1 _10231_ (.A1(_04268_),
    .A2(_04923_),
    .B1(_04943_),
    .C1(_04149_),
    .X(_04944_));
 sky130_fd_sc_hd__clkbuf_4 _10232_ (.A(net82),
    .X(_04945_));
 sky130_fd_sc_hd__a21o_1 _10233_ (.A1(net48),
    .A2(_04745_),
    .B1(_04666_),
    .X(_04946_));
 sky130_fd_sc_hd__a221o_1 _10234_ (.A1(_03637_),
    .A2(_04945_),
    .B1(_04673_),
    .B2(_04946_),
    .C1(_04266_),
    .X(_04947_));
 sky130_fd_sc_hd__o22a_1 _10235_ (.A1(\irq_pending[23] ),
    .A2(_04006_),
    .B1(_04944_),
    .B2(_04947_),
    .X(_04948_));
 sky130_fd_sc_hd__a31o_1 _10236_ (.A1(_04391_),
    .A2(_04920_),
    .A3(_04921_),
    .B1(_04948_),
    .X(_08384_));
 sky130_fd_sc_hd__or3_1 _10237_ (.A(_04877_),
    .B(_04886_),
    .C(_04919_),
    .X(_04949_));
 sky130_fd_sc_hd__or2b_1 _10238_ (.A(_04821_),
    .B_N(_04876_),
    .X(_04950_));
 sky130_fd_sc_hd__a211o_1 _10239_ (.A1(_04875_),
    .A2(_04950_),
    .B1(_04919_),
    .C1(_04886_),
    .X(_04951_));
 sky130_fd_sc_hd__nor2_1 _10240_ (.A(\reg_pc[23] ),
    .B(\decoded_imm[23] ),
    .Y(_04952_));
 sky130_fd_sc_hd__o21a_1 _10241_ (.A1(_04884_),
    .A2(_04952_),
    .B1(_04917_),
    .X(_04953_));
 sky130_fd_sc_hd__o211a_1 _10242_ (.A1(_04824_),
    .A2(_04949_),
    .B1(_04951_),
    .C1(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__nand2_1 _10243_ (.A(\reg_pc[24] ),
    .B(\decoded_imm[24] ),
    .Y(_04955_));
 sky130_fd_sc_hd__or2_1 _10244_ (.A(\reg_pc[24] ),
    .B(\decoded_imm[24] ),
    .X(_04956_));
 sky130_fd_sc_hd__nand2_1 _10245_ (.A(_04955_),
    .B(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__xor2_1 _10246_ (.A(_04954_),
    .B(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__clkbuf_4 _10247_ (.A(net83),
    .X(_04959_));
 sky130_fd_sc_hd__a21o_2 _10248_ (.A1(net49),
    .A2(_04811_),
    .B1(_04667_),
    .X(_04960_));
 sky130_fd_sc_hd__a22o_1 _10249_ (.A1(\count_instr[56] ),
    .A2(_04015_),
    .B1(_04017_),
    .B2(\count_cycle[56] ),
    .X(_04961_));
 sky130_fd_sc_hd__a221o_1 _10250_ (.A1(\count_instr[24] ),
    .A2(_04145_),
    .B1(\count_cycle[24] ),
    .B2(_03253_),
    .C1(_04961_),
    .X(_04962_));
 sky130_fd_sc_hd__mux4_1 _10251_ (.A0(\cpuregs.regs[12][24] ),
    .A1(\cpuregs.regs[13][24] ),
    .A2(\cpuregs.regs[14][24] ),
    .A3(\cpuregs.regs[15][24] ),
    .S0(_04217_),
    .S1(_04219_),
    .X(_04963_));
 sky130_fd_sc_hd__mux4_1 _10252_ (.A0(\cpuregs.regs[8][24] ),
    .A1(\cpuregs.regs[9][24] ),
    .A2(\cpuregs.regs[10][24] ),
    .A3(\cpuregs.regs[11][24] ),
    .S0(_04216_),
    .S1(_04376_),
    .X(_04964_));
 sky130_fd_sc_hd__or2_1 _10253_ (.A(_04369_),
    .B(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__o211a_1 _10254_ (.A1(_04211_),
    .A2(_04963_),
    .B1(_04965_),
    .C1(_04328_),
    .X(_04966_));
 sky130_fd_sc_hd__mux4_1 _10255_ (.A0(\cpuregs.regs[4][24] ),
    .A1(\cpuregs.regs[5][24] ),
    .A2(\cpuregs.regs[6][24] ),
    .A3(\cpuregs.regs[7][24] ),
    .S0(_04290_),
    .S1(_04276_),
    .X(_04967_));
 sky130_fd_sc_hd__mux4_1 _10256_ (.A0(\cpuregs.regs[0][24] ),
    .A1(\cpuregs.regs[1][24] ),
    .A2(\cpuregs.regs[2][24] ),
    .A3(\cpuregs.regs[3][24] ),
    .S0(_04290_),
    .S1(_04276_),
    .X(_04968_));
 sky130_fd_sc_hd__mux2_1 _10257_ (.A0(_04967_),
    .A1(_04968_),
    .S(_04222_),
    .X(_04969_));
 sky130_fd_sc_hd__a21o_1 _10258_ (.A1(_04214_),
    .A2(_04969_),
    .B1(_04237_),
    .X(_04970_));
 sky130_fd_sc_hd__mux4_1 _10259_ (.A0(\cpuregs.regs[28][24] ),
    .A1(\cpuregs.regs[29][24] ),
    .A2(\cpuregs.regs[30][24] ),
    .A3(\cpuregs.regs[31][24] ),
    .S0(_04329_),
    .S1(_04218_),
    .X(_04971_));
 sky130_fd_sc_hd__mux4_1 _10260_ (.A0(\cpuregs.regs[24][24] ),
    .A1(\cpuregs.regs[25][24] ),
    .A2(\cpuregs.regs[26][24] ),
    .A3(\cpuregs.regs[27][24] ),
    .S0(_04329_),
    .S1(_04218_),
    .X(_04972_));
 sky130_fd_sc_hd__mux2_1 _10261_ (.A0(_04971_),
    .A1(_04972_),
    .S(_04222_),
    .X(_04973_));
 sky130_fd_sc_hd__mux4_1 _10262_ (.A0(\cpuregs.regs[20][24] ),
    .A1(\cpuregs.regs[21][24] ),
    .A2(\cpuregs.regs[22][24] ),
    .A3(\cpuregs.regs[23][24] ),
    .S0(_04071_),
    .S1(_04073_),
    .X(_04974_));
 sky130_fd_sc_hd__mux4_1 _10263_ (.A0(\cpuregs.regs[16][24] ),
    .A1(\cpuregs.regs[17][24] ),
    .A2(\cpuregs.regs[18][24] ),
    .A3(\cpuregs.regs[19][24] ),
    .S0(_04071_),
    .S1(_04073_),
    .X(_04975_));
 sky130_fd_sc_hd__mux2_1 _10264_ (.A0(_04974_),
    .A1(_04975_),
    .S(_04077_),
    .X(_04976_));
 sky130_fd_sc_hd__a21o_1 _10265_ (.A1(_04068_),
    .A2(_04976_),
    .B1(_04080_),
    .X(_04977_));
 sky130_fd_sc_hd__a21o_1 _10266_ (.A1(_04328_),
    .A2(_04973_),
    .B1(_04977_),
    .X(_04978_));
 sky130_fd_sc_hd__o211a_4 _10267_ (.A1(_04966_),
    .A2(_04970_),
    .B1(_04978_),
    .C1(_04133_),
    .X(_04979_));
 sky130_fd_sc_hd__a221o_1 _10268_ (.A1(\irq_mask[24] ),
    .A2(_04308_),
    .B1(\timer[24] ),
    .B2(instr_timer),
    .C1(_04025_),
    .X(_04980_));
 sky130_fd_sc_hd__a21o_1 _10269_ (.A1(instr_retirq),
    .A2(_04979_),
    .B1(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__o211a_1 _10270_ (.A1(_04268_),
    .A2(_04962_),
    .B1(_04981_),
    .C1(_04149_),
    .X(_04982_));
 sky130_fd_sc_hd__a221o_1 _10271_ (.A1(_03638_),
    .A2(_04959_),
    .B1(_04752_),
    .B2(_04960_),
    .C1(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__a221o_1 _10272_ (.A1(\irq_pending[24] ),
    .A2(_04049_),
    .B1(_04958_),
    .B2(_03385_),
    .C1(_04983_),
    .X(_08385_));
 sky130_fd_sc_hd__o21ai_2 _10273_ (.A1(_04954_),
    .A2(_04957_),
    .B1(_04955_),
    .Y(_04984_));
 sky130_fd_sc_hd__and2_1 _10274_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .X(_04985_));
 sky130_fd_sc_hd__nor2_1 _10275_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .Y(_04986_));
 sky130_fd_sc_hd__nor2_1 _10276_ (.A(_04985_),
    .B(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__or2_1 _10277_ (.A(_04984_),
    .B(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__nand2_1 _10278_ (.A(_04984_),
    .B(_04987_),
    .Y(_04989_));
 sky130_fd_sc_hd__and3_1 _10279_ (.A(_03384_),
    .B(_04988_),
    .C(_04989_),
    .X(_04990_));
 sky130_fd_sc_hd__a22o_1 _10280_ (.A1(\count_instr[57] ),
    .A2(_04016_),
    .B1(_04105_),
    .B2(\count_cycle[57] ),
    .X(_04991_));
 sky130_fd_sc_hd__a221o_1 _10281_ (.A1(\count_instr[25] ),
    .A2(_04012_),
    .B1(\count_cycle[25] ),
    .B2(_04165_),
    .C1(_04991_),
    .X(_04992_));
 sky130_fd_sc_hd__mux4_1 _10282_ (.A0(\cpuregs.regs[20][25] ),
    .A1(\cpuregs.regs[21][25] ),
    .A2(\cpuregs.regs[22][25] ),
    .A3(\cpuregs.regs[23][25] ),
    .S0(_04275_),
    .S1(_04278_),
    .X(_04993_));
 sky130_fd_sc_hd__mux4_1 _10283_ (.A0(\cpuregs.regs[16][25] ),
    .A1(\cpuregs.regs[17][25] ),
    .A2(\cpuregs.regs[18][25] ),
    .A3(\cpuregs.regs[19][25] ),
    .S0(_04291_),
    .S1(_04292_),
    .X(_04994_));
 sky130_fd_sc_hd__or2_1 _10284_ (.A(_04430_),
    .B(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__o211a_1 _10285_ (.A1(_04287_),
    .A2(_04993_),
    .B1(_04995_),
    .C1(_04289_),
    .X(_04996_));
 sky130_fd_sc_hd__mux4_1 _10286_ (.A0(\cpuregs.regs[28][25] ),
    .A1(\cpuregs.regs[29][25] ),
    .A2(\cpuregs.regs[30][25] ),
    .A3(\cpuregs.regs[31][25] ),
    .S0(_04291_),
    .S1(_04292_),
    .X(_04997_));
 sky130_fd_sc_hd__mux4_1 _10287_ (.A0(\cpuregs.regs[24][25] ),
    .A1(\cpuregs.regs[25][25] ),
    .A2(\cpuregs.regs[26][25] ),
    .A3(\cpuregs.regs[27][25] ),
    .S0(_04291_),
    .S1(_04292_),
    .X(_04998_));
 sky130_fd_sc_hd__mux2_1 _10288_ (.A0(_04997_),
    .A1(_04998_),
    .S(_04223_),
    .X(_04999_));
 sky130_fd_sc_hd__a21o_1 _10289_ (.A1(_04206_),
    .A2(_04999_),
    .B1(_04225_),
    .X(_05000_));
 sky130_fd_sc_hd__mux4_1 _10290_ (.A0(\cpuregs.regs[4][25] ),
    .A1(\cpuregs.regs[5][25] ),
    .A2(\cpuregs.regs[6][25] ),
    .A3(\cpuregs.regs[7][25] ),
    .S0(_04291_),
    .S1(_04292_),
    .X(_05001_));
 sky130_fd_sc_hd__or2_1 _10291_ (.A(_04223_),
    .B(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__mux4_1 _10292_ (.A0(\cpuregs.regs[0][25] ),
    .A1(\cpuregs.regs[1][25] ),
    .A2(\cpuregs.regs[2][25] ),
    .A3(\cpuregs.regs[3][25] ),
    .S0(_04217_),
    .S1(_04219_),
    .X(_05003_));
 sky130_fd_sc_hd__o21a_1 _10293_ (.A1(_04430_),
    .A2(_05003_),
    .B1(_04214_),
    .X(_05004_));
 sky130_fd_sc_hd__mux4_1 _10294_ (.A0(\cpuregs.regs[12][25] ),
    .A1(\cpuregs.regs[13][25] ),
    .A2(\cpuregs.regs[14][25] ),
    .A3(\cpuregs.regs[15][25] ),
    .S0(_04325_),
    .S1(_04277_),
    .X(_05005_));
 sky130_fd_sc_hd__mux4_1 _10295_ (.A0(\cpuregs.regs[8][25] ),
    .A1(\cpuregs.regs[9][25] ),
    .A2(\cpuregs.regs[10][25] ),
    .A3(\cpuregs.regs[11][25] ),
    .S0(_04325_),
    .S1(_04277_),
    .X(_05006_));
 sky130_fd_sc_hd__mux2_1 _10296_ (.A0(_05005_),
    .A1(_05006_),
    .S(_04321_),
    .X(_05007_));
 sky130_fd_sc_hd__a221o_1 _10297_ (.A1(_05002_),
    .A2(_05004_),
    .B1(_05007_),
    .B2(_04206_),
    .C1(_04296_),
    .X(_05008_));
 sky130_fd_sc_hd__o211a_4 _10298_ (.A1(_04996_),
    .A2(_05000_),
    .B1(_04133_),
    .C1(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__a221o_1 _10299_ (.A1(\irq_mask[25] ),
    .A2(_04448_),
    .B1(\timer[25] ),
    .B2(_04187_),
    .C1(_04188_),
    .X(_05010_));
 sky130_fd_sc_hd__a21o_1 _10300_ (.A1(_04168_),
    .A2(_05009_),
    .B1(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__o211a_1 _10301_ (.A1(_04010_),
    .A2(_04992_),
    .B1(_05011_),
    .C1(_04150_),
    .X(_05012_));
 sky130_fd_sc_hd__clkbuf_4 _10302_ (.A(net84),
    .X(_05013_));
 sky130_fd_sc_hd__a21o_2 _10303_ (.A1(net50),
    .A2(_04811_),
    .B1(_04667_),
    .X(_05014_));
 sky130_fd_sc_hd__a221o_1 _10304_ (.A1(_03680_),
    .A2(_05013_),
    .B1(_04752_),
    .B2(_05014_),
    .C1(_04202_),
    .X(_05015_));
 sky130_fd_sc_hd__o32a_1 _10305_ (.A1(_04990_),
    .A2(_05012_),
    .A3(_05015_),
    .B1(_04007_),
    .B2(\irq_pending[25] ),
    .X(_08386_));
 sky130_fd_sc_hd__nand2_1 _10306_ (.A(\reg_pc[26] ),
    .B(\decoded_imm[26] ),
    .Y(_05016_));
 sky130_fd_sc_hd__or2_1 _10307_ (.A(\reg_pc[26] ),
    .B(\decoded_imm[26] ),
    .X(_05017_));
 sky130_fd_sc_hd__nand2_1 _10308_ (.A(_05016_),
    .B(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__a21oi_2 _10309_ (.A1(_04984_),
    .A2(_04987_),
    .B1(_04985_),
    .Y(_05019_));
 sky130_fd_sc_hd__xor2_1 _10310_ (.A(_05018_),
    .B(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__mux4_1 _10311_ (.A0(\cpuregs.regs[28][26] ),
    .A1(\cpuregs.regs[29][26] ),
    .A2(\cpuregs.regs[30][26] ),
    .A3(\cpuregs.regs[31][26] ),
    .S0(_04084_),
    .S1(_04086_),
    .X(_05021_));
 sky130_fd_sc_hd__mux4_1 _10312_ (.A0(\cpuregs.regs[24][26] ),
    .A1(\cpuregs.regs[25][26] ),
    .A2(\cpuregs.regs[26][26] ),
    .A3(\cpuregs.regs[27][26] ),
    .S0(_04084_),
    .S1(_04086_),
    .X(_05022_));
 sky130_fd_sc_hd__mux2_1 _10313_ (.A0(_05021_),
    .A1(_05022_),
    .S(_04077_),
    .X(_05023_));
 sky130_fd_sc_hd__nand2_1 _10314_ (.A(_04052_),
    .B(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__mux4_1 _10315_ (.A0(\cpuregs.regs[20][26] ),
    .A1(\cpuregs.regs[21][26] ),
    .A2(\cpuregs.regs[22][26] ),
    .A3(\cpuregs.regs[23][26] ),
    .S0(_04123_),
    .S1(_04124_),
    .X(_05025_));
 sky130_fd_sc_hd__mux4_1 _10316_ (.A0(\cpuregs.regs[16][26] ),
    .A1(\cpuregs.regs[17][26] ),
    .A2(\cpuregs.regs[18][26] ),
    .A3(\cpuregs.regs[19][26] ),
    .S0(_04123_),
    .S1(_04124_),
    .X(_05026_));
 sky130_fd_sc_hd__mux2_1 _10317_ (.A0(_05025_),
    .A1(_05026_),
    .S(_04077_),
    .X(_05027_));
 sky130_fd_sc_hd__a21oi_1 _10318_ (.A1(_04068_),
    .A2(_05027_),
    .B1(_04080_),
    .Y(_05028_));
 sky130_fd_sc_hd__mux4_1 _10319_ (.A0(\cpuregs.regs[8][26] ),
    .A1(\cpuregs.regs[9][26] ),
    .A2(\cpuregs.regs[10][26] ),
    .A3(\cpuregs.regs[11][26] ),
    .S0(_04071_),
    .S1(_04073_),
    .X(_05029_));
 sky130_fd_sc_hd__mux4_1 _10320_ (.A0(\cpuregs.regs[12][26] ),
    .A1(\cpuregs.regs[13][26] ),
    .A2(\cpuregs.regs[14][26] ),
    .A3(\cpuregs.regs[15][26] ),
    .S0(_04123_),
    .S1(_04124_),
    .X(_05030_));
 sky130_fd_sc_hd__mux2_1 _10321_ (.A0(_05029_),
    .A1(_05030_),
    .S(_00071_),
    .X(_05031_));
 sky130_fd_sc_hd__mux4_1 _10322_ (.A0(\cpuregs.regs[4][26] ),
    .A1(\cpuregs.regs[5][26] ),
    .A2(\cpuregs.regs[6][26] ),
    .A3(\cpuregs.regs[7][26] ),
    .S0(_04055_),
    .S1(_04058_),
    .X(_05032_));
 sky130_fd_sc_hd__mux4_1 _10323_ (.A0(\cpuregs.regs[0][26] ),
    .A1(\cpuregs.regs[1][26] ),
    .A2(\cpuregs.regs[2][26] ),
    .A3(\cpuregs.regs[3][26] ),
    .S0(_04055_),
    .S1(_04058_),
    .X(_05033_));
 sky130_fd_sc_hd__mux2_1 _10324_ (.A0(_05032_),
    .A1(_05033_),
    .S(_04063_),
    .X(_05034_));
 sky130_fd_sc_hd__a21o_1 _10325_ (.A1(_04068_),
    .A2(_05034_),
    .B1(_00073_),
    .X(_05035_));
 sky130_fd_sc_hd__a21oi_1 _10326_ (.A1(_04052_),
    .A2(_05031_),
    .B1(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__a211o_4 _10327_ (.A1(_05024_),
    .A2(_05028_),
    .B1(net301),
    .C1(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__nor2_1 _10328_ (.A(_04051_),
    .B(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__a221o_1 _10329_ (.A1(\irq_mask[26] ),
    .A2(_04448_),
    .B1(\timer[26] ),
    .B2(_04187_),
    .C1(_04027_),
    .X(_05039_));
 sky130_fd_sc_hd__a22o_1 _10330_ (.A1(\count_instr[58] ),
    .A2(_04015_),
    .B1(instr_rdcycleh),
    .B2(\count_cycle[58] ),
    .X(_05040_));
 sky130_fd_sc_hd__a211o_1 _10331_ (.A1(\count_instr[26] ),
    .A2(_04145_),
    .B1(_04009_),
    .C1(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__a21o_1 _10332_ (.A1(\count_cycle[26] ),
    .A2(_04165_),
    .B1(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__o211a_1 _10333_ (.A1(_05038_),
    .A2(_05039_),
    .B1(_05042_),
    .C1(_03302_),
    .X(_05043_));
 sky130_fd_sc_hd__clkbuf_4 _10334_ (.A(net85),
    .X(_05044_));
 sky130_fd_sc_hd__a21o_1 _10335_ (.A1(net51),
    .A2(_04811_),
    .B1(_04667_),
    .X(_05045_));
 sky130_fd_sc_hd__a221o_1 _10336_ (.A1(_04046_),
    .A2(_05044_),
    .B1(_04752_),
    .B2(_05045_),
    .C1(_04202_),
    .X(_05046_));
 sky130_fd_sc_hd__o22a_1 _10337_ (.A1(\irq_pending[26] ),
    .A2(_04007_),
    .B1(_05043_),
    .B2(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__a21o_1 _10338_ (.A1(_04391_),
    .A2(_05020_),
    .B1(_05047_),
    .X(_08387_));
 sky130_fd_sc_hd__o21ai_1 _10339_ (.A1(_05018_),
    .A2(_05019_),
    .B1(_05016_),
    .Y(_05048_));
 sky130_fd_sc_hd__nor2_1 _10340_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .Y(_05049_));
 sky130_fd_sc_hd__and2_1 _10341_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .X(_05050_));
 sky130_fd_sc_hd__or2_1 _10342_ (.A(_05049_),
    .B(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__xnor2_1 _10343_ (.A(_05048_),
    .B(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__mux4_1 _10344_ (.A0(\cpuregs.regs[28][27] ),
    .A1(\cpuregs.regs[29][27] ),
    .A2(\cpuregs.regs[30][27] ),
    .A3(\cpuregs.regs[31][27] ),
    .S0(_04758_),
    .S1(_04759_),
    .X(_05053_));
 sky130_fd_sc_hd__mux4_1 _10345_ (.A0(\cpuregs.regs[24][27] ),
    .A1(\cpuregs.regs[25][27] ),
    .A2(\cpuregs.regs[26][27] ),
    .A3(\cpuregs.regs[27][27] ),
    .S0(_04758_),
    .S1(_04759_),
    .X(_05054_));
 sky130_fd_sc_hd__mux2_1 _10346_ (.A0(_05053_),
    .A1(_05054_),
    .S(_04211_),
    .X(_05055_));
 sky130_fd_sc_hd__nand2_1 _10347_ (.A(_04272_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__mux4_1 _10348_ (.A0(\cpuregs.regs[20][27] ),
    .A1(\cpuregs.regs[21][27] ),
    .A2(\cpuregs.regs[22][27] ),
    .A3(\cpuregs.regs[23][27] ),
    .S0(_04207_),
    .S1(_04208_),
    .X(_05057_));
 sky130_fd_sc_hd__mux4_1 _10349_ (.A0(\cpuregs.regs[16][27] ),
    .A1(\cpuregs.regs[17][27] ),
    .A2(\cpuregs.regs[18][27] ),
    .A3(\cpuregs.regs[19][27] ),
    .S0(_04207_),
    .S1(_04208_),
    .X(_05058_));
 sky130_fd_sc_hd__mux2_1 _10350_ (.A0(_05057_),
    .A1(_05058_),
    .S(_04211_),
    .X(_05059_));
 sky130_fd_sc_hd__a21oi_1 _10351_ (.A1(_04215_),
    .A2(_05059_),
    .B1(_04225_),
    .Y(_05060_));
 sky130_fd_sc_hd__mux4_1 _10352_ (.A0(\cpuregs.regs[4][27] ),
    .A1(\cpuregs.regs[5][27] ),
    .A2(\cpuregs.regs[6][27] ),
    .A3(\cpuregs.regs[7][27] ),
    .S0(_04207_),
    .S1(_04208_),
    .X(_05061_));
 sky130_fd_sc_hd__mux4_1 _10353_ (.A0(\cpuregs.regs[0][27] ),
    .A1(\cpuregs.regs[1][27] ),
    .A2(\cpuregs.regs[2][27] ),
    .A3(\cpuregs.regs[3][27] ),
    .S0(_04207_),
    .S1(_04208_),
    .X(_05062_));
 sky130_fd_sc_hd__mux2_1 _10354_ (.A0(_05061_),
    .A1(_05062_),
    .S(_04211_),
    .X(_05063_));
 sky130_fd_sc_hd__mux4_1 _10355_ (.A0(\cpuregs.regs[12][27] ),
    .A1(\cpuregs.regs[13][27] ),
    .A2(\cpuregs.regs[14][27] ),
    .A3(\cpuregs.regs[15][27] ),
    .S0(_04057_),
    .S1(_04060_),
    .X(_05064_));
 sky130_fd_sc_hd__mux4_1 _10356_ (.A0(\cpuregs.regs[8][27] ),
    .A1(\cpuregs.regs[9][27] ),
    .A2(\cpuregs.regs[10][27] ),
    .A3(\cpuregs.regs[11][27] ),
    .S0(_04057_),
    .S1(_04060_),
    .X(_05065_));
 sky130_fd_sc_hd__mux2_1 _10357_ (.A0(_05064_),
    .A1(_05065_),
    .S(_04065_),
    .X(_05066_));
 sky130_fd_sc_hd__a21o_1 _10358_ (.A1(_04231_),
    .A2(_05066_),
    .B1(_04237_),
    .X(_05067_));
 sky130_fd_sc_hd__a21oi_1 _10359_ (.A1(_04215_),
    .A2(_05063_),
    .B1(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__a211o_4 _10360_ (.A1(_05056_),
    .A2(_05060_),
    .B1(_04227_),
    .C1(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__nor2_1 _10361_ (.A(_04051_),
    .B(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__a221o_1 _10362_ (.A1(\irq_mask[27] ),
    .A2(_04448_),
    .B1(\timer[27] ),
    .B2(_04187_),
    .C1(_04188_),
    .X(_05071_));
 sky130_fd_sc_hd__a22o_1 _10363_ (.A1(\count_instr[59] ),
    .A2(_04015_),
    .B1(instr_rdcycleh),
    .B2(\count_cycle[59] ),
    .X(_05072_));
 sky130_fd_sc_hd__a211o_1 _10364_ (.A1(\count_instr[27] ),
    .A2(_04011_),
    .B1(_04009_),
    .C1(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__a21o_1 _10365_ (.A1(\count_cycle[27] ),
    .A2(_04165_),
    .B1(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__o211a_1 _10366_ (.A1(_05070_),
    .A2(_05071_),
    .B1(_05074_),
    .C1(_03302_),
    .X(_05075_));
 sky130_fd_sc_hd__clkbuf_4 _10367_ (.A(net86),
    .X(_05076_));
 sky130_fd_sc_hd__a21o_1 _10368_ (.A1(net52),
    .A2(_04811_),
    .B1(_04666_),
    .X(_05077_));
 sky130_fd_sc_hd__a221o_1 _10369_ (.A1(_04046_),
    .A2(_05076_),
    .B1(_04752_),
    .B2(_05077_),
    .C1(_04202_),
    .X(_05078_));
 sky130_fd_sc_hd__o22a_1 _10370_ (.A1(\irq_pending[27] ),
    .A2(_04007_),
    .B1(_05075_),
    .B2(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__a21o_1 _10371_ (.A1(_04391_),
    .A2(_05052_),
    .B1(_05079_),
    .X(_08388_));
 sky130_fd_sc_hd__nand2_1 _10372_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .Y(_05080_));
 sky130_fd_sc_hd__nor2_1 _10373_ (.A(_05017_),
    .B(_05050_),
    .Y(_05081_));
 sky130_fd_sc_hd__a311o_1 _10374_ (.A1(_05016_),
    .A2(_05019_),
    .A3(_05080_),
    .B1(_05081_),
    .C1(_05049_),
    .X(_05082_));
 sky130_fd_sc_hd__xnor2_1 _10375_ (.A(\reg_pc[28] ),
    .B(\decoded_imm[28] ),
    .Y(_05083_));
 sky130_fd_sc_hd__nor2_1 _10376_ (.A(_05082_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__a21o_1 _10377_ (.A1(_05082_),
    .A2(_05083_),
    .B1(_04156_),
    .X(_05085_));
 sky130_fd_sc_hd__buf_4 _10378_ (.A(net87),
    .X(_05086_));
 sky130_fd_sc_hd__a21o_1 _10379_ (.A1(net53),
    .A2(_04811_),
    .B1(_04667_),
    .X(_05087_));
 sky130_fd_sc_hd__a22o_1 _10380_ (.A1(\count_instr[60] ),
    .A2(_04015_),
    .B1(instr_rdinstr),
    .B2(\count_instr[28] ),
    .X(_05088_));
 sky130_fd_sc_hd__a221o_1 _10381_ (.A1(_04105_),
    .A2(\count_cycle[60] ),
    .B1(_03253_),
    .B2(\count_cycle[28] ),
    .C1(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__mux4_1 _10382_ (.A0(\cpuregs.regs[24][28] ),
    .A1(\cpuregs.regs[25][28] ),
    .A2(\cpuregs.regs[26][28] ),
    .A3(\cpuregs.regs[27][28] ),
    .S0(_04216_),
    .S1(_04376_),
    .X(_05090_));
 sky130_fd_sc_hd__mux4_1 _10383_ (.A0(\cpuregs.regs[28][28] ),
    .A1(\cpuregs.regs[29][28] ),
    .A2(\cpuregs.regs[30][28] ),
    .A3(\cpuregs.regs[31][28] ),
    .S0(_04216_),
    .S1(_04376_),
    .X(_05091_));
 sky130_fd_sc_hd__mux2_1 _10384_ (.A0(_05090_),
    .A1(_05091_),
    .S(_04369_),
    .X(_05092_));
 sky130_fd_sc_hd__nand2_1 _10385_ (.A(_04328_),
    .B(_05092_),
    .Y(_05093_));
 sky130_fd_sc_hd__mux4_1 _10386_ (.A0(\cpuregs.regs[20][28] ),
    .A1(\cpuregs.regs[21][28] ),
    .A2(\cpuregs.regs[22][28] ),
    .A3(\cpuregs.regs[23][28] ),
    .S0(_04273_),
    .S1(_04283_),
    .X(_05094_));
 sky130_fd_sc_hd__mux4_1 _10387_ (.A0(\cpuregs.regs[16][28] ),
    .A1(\cpuregs.regs[17][28] ),
    .A2(\cpuregs.regs[18][28] ),
    .A3(\cpuregs.regs[19][28] ),
    .S0(_04273_),
    .S1(_04283_),
    .X(_05095_));
 sky130_fd_sc_hd__mux2_1 _10388_ (.A0(_05094_),
    .A1(_05095_),
    .S(_04320_),
    .X(_05096_));
 sky130_fd_sc_hd__a21oi_1 _10389_ (.A1(_04214_),
    .A2(_05096_),
    .B1(_04081_),
    .Y(_05097_));
 sky130_fd_sc_hd__mux4_1 _10390_ (.A0(\cpuregs.regs[4][28] ),
    .A1(\cpuregs.regs[5][28] ),
    .A2(\cpuregs.regs[6][28] ),
    .A3(\cpuregs.regs[7][28] ),
    .S0(_04290_),
    .S1(_04283_),
    .X(_05098_));
 sky130_fd_sc_hd__mux4_1 _10391_ (.A0(\cpuregs.regs[0][28] ),
    .A1(\cpuregs.regs[1][28] ),
    .A2(\cpuregs.regs[2][28] ),
    .A3(\cpuregs.regs[3][28] ),
    .S0(_04273_),
    .S1(_04283_),
    .X(_05099_));
 sky130_fd_sc_hd__mux2_1 _10392_ (.A0(_05098_),
    .A1(_05099_),
    .S(_04222_),
    .X(_05100_));
 sky130_fd_sc_hd__mux4_1 _10393_ (.A0(\cpuregs.regs[12][28] ),
    .A1(\cpuregs.regs[13][28] ),
    .A2(\cpuregs.regs[14][28] ),
    .A3(\cpuregs.regs[15][28] ),
    .S0(_04123_),
    .S1(_04124_),
    .X(_05101_));
 sky130_fd_sc_hd__mux4_1 _10394_ (.A0(\cpuregs.regs[8][28] ),
    .A1(\cpuregs.regs[9][28] ),
    .A2(\cpuregs.regs[10][28] ),
    .A3(\cpuregs.regs[11][28] ),
    .S0(_04123_),
    .S1(_04124_),
    .X(_05102_));
 sky130_fd_sc_hd__mux2_1 _10395_ (.A0(_05101_),
    .A1(_05102_),
    .S(_04077_),
    .X(_05103_));
 sky130_fd_sc_hd__a21o_1 _10396_ (.A1(_04052_),
    .A2(_05103_),
    .B1(_00073_),
    .X(_05104_));
 sky130_fd_sc_hd__a21oi_1 _10397_ (.A1(_04214_),
    .A2(_05100_),
    .B1(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__a211o_2 _10398_ (.A1(_05093_),
    .A2(_05097_),
    .B1(net301),
    .C1(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__inv_2 _10399_ (.A(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__a221o_1 _10400_ (.A1(\irq_mask[28] ),
    .A2(instr_maskirq),
    .B1(\timer[28] ),
    .B2(instr_timer),
    .C1(_04025_),
    .X(_05108_));
 sky130_fd_sc_hd__a21o_1 _10401_ (.A1(instr_retirq),
    .A2(_05107_),
    .B1(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__o211a_1 _10402_ (.A1(_04009_),
    .A2(_05089_),
    .B1(_05109_),
    .C1(_03301_),
    .X(_05110_));
 sky130_fd_sc_hd__a221o_1 _10403_ (.A1(_03680_),
    .A2(_05086_),
    .B1(_04752_),
    .B2(_05087_),
    .C1(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__a21oi_1 _10404_ (.A1(\irq_pending[28] ),
    .A2(_04049_),
    .B1(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__o21ai_1 _10405_ (.A1(_05084_),
    .A2(_05085_),
    .B1(_05112_),
    .Y(_08389_));
 sky130_fd_sc_hd__nand2_1 _10406_ (.A(\reg_pc[29] ),
    .B(\decoded_imm[29] ),
    .Y(_05113_));
 sky130_fd_sc_hd__or2_1 _10407_ (.A(\reg_pc[29] ),
    .B(\decoded_imm[29] ),
    .X(_05114_));
 sky130_fd_sc_hd__and2_1 _10408_ (.A(_05113_),
    .B(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__a211o_1 _10409_ (.A1(\reg_pc[28] ),
    .A2(\decoded_imm[28] ),
    .B1(_05084_),
    .C1(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__nand2_1 _10410_ (.A(_05084_),
    .B(_05115_),
    .Y(_05117_));
 sky130_fd_sc_hd__nand3_1 _10411_ (.A(\reg_pc[28] ),
    .B(\decoded_imm[28] ),
    .C(_05115_),
    .Y(_05118_));
 sky130_fd_sc_hd__and4_1 _10412_ (.A(_03384_),
    .B(_05116_),
    .C(_05117_),
    .D(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__a22o_1 _10413_ (.A1(\count_instr[61] ),
    .A2(_04016_),
    .B1(_04145_),
    .B2(\count_instr[29] ),
    .X(_05120_));
 sky130_fd_sc_hd__a221o_1 _10414_ (.A1(_04018_),
    .A2(\count_cycle[61] ),
    .B1(_04014_),
    .B2(\count_cycle[29] ),
    .C1(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__mux4_1 _10415_ (.A0(\cpuregs.regs[28][29] ),
    .A1(\cpuregs.regs[29][29] ),
    .A2(\cpuregs.regs[30][29] ),
    .A3(\cpuregs.regs[31][29] ),
    .S0(_04579_),
    .S1(_04284_),
    .X(_05122_));
 sky130_fd_sc_hd__mux4_1 _10416_ (.A0(\cpuregs.regs[24][29] ),
    .A1(\cpuregs.regs[25][29] ),
    .A2(\cpuregs.regs[26][29] ),
    .A3(\cpuregs.regs[27][29] ),
    .S0(_04579_),
    .S1(_04284_),
    .X(_05123_));
 sky130_fd_sc_hd__mux2_1 _10417_ (.A0(_05122_),
    .A1(_05123_),
    .S(_04575_),
    .X(_05124_));
 sky130_fd_sc_hd__nand2_1 _10418_ (.A(_04054_),
    .B(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__mux4_1 _10419_ (.A0(\cpuregs.regs[20][29] ),
    .A1(\cpuregs.regs[21][29] ),
    .A2(\cpuregs.regs[22][29] ),
    .A3(\cpuregs.regs[23][29] ),
    .S0(_04477_),
    .S1(_04478_),
    .X(_05126_));
 sky130_fd_sc_hd__mux4_1 _10420_ (.A0(\cpuregs.regs[16][29] ),
    .A1(\cpuregs.regs[17][29] ),
    .A2(\cpuregs.regs[18][29] ),
    .A3(\cpuregs.regs[19][29] ),
    .S0(_04477_),
    .S1(_04478_),
    .X(_05127_));
 sky130_fd_sc_hd__mux2_1 _10421_ (.A0(_05126_),
    .A1(_05127_),
    .S(_04121_),
    .X(_05128_));
 sky130_fd_sc_hd__a21oi_1 _10422_ (.A1(_04070_),
    .A2(_05128_),
    .B1(_04082_),
    .Y(_05129_));
 sky130_fd_sc_hd__mux4_1 _10423_ (.A0(\cpuregs.regs[8][29] ),
    .A1(\cpuregs.regs[9][29] ),
    .A2(\cpuregs.regs[10][29] ),
    .A3(\cpuregs.regs[11][29] ),
    .S0(_04057_),
    .S1(_04060_),
    .X(_05130_));
 sky130_fd_sc_hd__mux4_1 _10424_ (.A0(\cpuregs.regs[12][29] ),
    .A1(\cpuregs.regs[13][29] ),
    .A2(\cpuregs.regs[14][29] ),
    .A3(\cpuregs.regs[15][29] ),
    .S0(_04057_),
    .S1(_04060_),
    .X(_05131_));
 sky130_fd_sc_hd__mux2_1 _10425_ (.A0(_05130_),
    .A1(_05131_),
    .S(_04430_),
    .X(_05132_));
 sky130_fd_sc_hd__mux4_1 _10426_ (.A0(\cpuregs.regs[4][29] ),
    .A1(\cpuregs.regs[5][29] ),
    .A2(\cpuregs.regs[6][29] ),
    .A3(\cpuregs.regs[7][29] ),
    .S0(_04273_),
    .S1(_04469_),
    .X(_05133_));
 sky130_fd_sc_hd__mux4_1 _10427_ (.A0(\cpuregs.regs[0][29] ),
    .A1(\cpuregs.regs[1][29] ),
    .A2(\cpuregs.regs[2][29] ),
    .A3(\cpuregs.regs[3][29] ),
    .S0(_04487_),
    .S1(_04469_),
    .X(_05134_));
 sky130_fd_sc_hd__mux2_1 _10428_ (.A0(_05133_),
    .A1(_05134_),
    .S(_04320_),
    .X(_05135_));
 sky130_fd_sc_hd__a21o_1 _10429_ (.A1(_04069_),
    .A2(_05135_),
    .B1(_04095_),
    .X(_05136_));
 sky130_fd_sc_hd__a21oi_1 _10430_ (.A1(_04054_),
    .A2(_05132_),
    .B1(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__a211o_2 _10431_ (.A1(_05125_),
    .A2(_05129_),
    .B1(_04100_),
    .C1(_05137_),
    .X(_05138_));
 sky130_fd_sc_hd__inv_2 _10432_ (.A(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__a221o_1 _10433_ (.A1(\irq_mask[29] ),
    .A2(_04448_),
    .B1(\timer[29] ),
    .B2(_04187_),
    .C1(_04188_),
    .X(_05140_));
 sky130_fd_sc_hd__a21o_1 _10434_ (.A1(_04168_),
    .A2(_05139_),
    .B1(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__o211a_1 _10435_ (.A1(_04010_),
    .A2(_05121_),
    .B1(_05141_),
    .C1(_04150_),
    .X(_05142_));
 sky130_fd_sc_hd__buf_4 _10436_ (.A(net88),
    .X(_05143_));
 sky130_fd_sc_hd__a21o_1 _10437_ (.A1(net54),
    .A2(_04811_),
    .B1(_04667_),
    .X(_05144_));
 sky130_fd_sc_hd__a221o_1 _10438_ (.A1(_03680_),
    .A2(_05143_),
    .B1(_04752_),
    .B2(_05144_),
    .C1(_04202_),
    .X(_05145_));
 sky130_fd_sc_hd__o32a_1 _10439_ (.A1(_05119_),
    .A2(_05142_),
    .A3(_05145_),
    .B1(_04007_),
    .B2(\irq_pending[29] ),
    .X(_08390_));
 sky130_fd_sc_hd__nand2_1 _10440_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .Y(_05146_));
 sky130_fd_sc_hd__or2_1 _10441_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .X(_05147_));
 sky130_fd_sc_hd__nand2_1 _10442_ (.A(_05146_),
    .B(_05147_),
    .Y(_05148_));
 sky130_fd_sc_hd__and3_1 _10443_ (.A(_05113_),
    .B(_05117_),
    .C(_05118_),
    .X(_05149_));
 sky130_fd_sc_hd__xor2_1 _10444_ (.A(_05148_),
    .B(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__a22o_1 _10445_ (.A1(\count_instr[62] ),
    .A2(_04104_),
    .B1(_04017_),
    .B2(\count_cycle[62] ),
    .X(_05151_));
 sky130_fd_sc_hd__a221o_1 _10446_ (.A1(\count_instr[30] ),
    .A2(_04012_),
    .B1(\count_cycle[30] ),
    .B2(_04013_),
    .C1(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__mux4_1 _10447_ (.A0(\cpuregs.regs[20][30] ),
    .A1(\cpuregs.regs[21][30] ),
    .A2(\cpuregs.regs[22][30] ),
    .A3(\cpuregs.regs[23][30] ),
    .S0(_04472_),
    .S1(_04473_),
    .X(_05153_));
 sky130_fd_sc_hd__mux4_1 _10448_ (.A0(\cpuregs.regs[16][30] ),
    .A1(\cpuregs.regs[17][30] ),
    .A2(\cpuregs.regs[18][30] ),
    .A3(\cpuregs.regs[19][30] ),
    .S0(_04472_),
    .S1(_04473_),
    .X(_05154_));
 sky130_fd_sc_hd__mux2_1 _10449_ (.A0(_05153_),
    .A1(_05154_),
    .S(_04065_),
    .X(_05155_));
 sky130_fd_sc_hd__nand2_1 _10450_ (.A(_04483_),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__mux4_1 _10451_ (.A0(\cpuregs.regs[28][30] ),
    .A1(\cpuregs.regs[29][30] ),
    .A2(\cpuregs.regs[30][30] ),
    .A3(\cpuregs.regs[31][30] ),
    .S0(_04085_),
    .S1(_04087_),
    .X(_05157_));
 sky130_fd_sc_hd__mux4_1 _10452_ (.A0(\cpuregs.regs[24][30] ),
    .A1(\cpuregs.regs[25][30] ),
    .A2(\cpuregs.regs[26][30] ),
    .A3(\cpuregs.regs[27][30] ),
    .S0(_04085_),
    .S1(_04087_),
    .X(_05158_));
 sky130_fd_sc_hd__mux2_1 _10453_ (.A0(_05157_),
    .A1(_05158_),
    .S(_04078_),
    .X(_05159_));
 sky130_fd_sc_hd__a21oi_1 _10454_ (.A1(_04231_),
    .A2(_05159_),
    .B1(_04082_),
    .Y(_05160_));
 sky130_fd_sc_hd__mux4_1 _10455_ (.A0(\cpuregs.regs[4][30] ),
    .A1(\cpuregs.regs[5][30] ),
    .A2(\cpuregs.regs[6][30] ),
    .A3(\cpuregs.regs[7][30] ),
    .S0(_04232_),
    .S1(_04233_),
    .X(_05161_));
 sky130_fd_sc_hd__mux4_1 _10456_ (.A0(\cpuregs.regs[0][30] ),
    .A1(\cpuregs.regs[1][30] ),
    .A2(\cpuregs.regs[2][30] ),
    .A3(\cpuregs.regs[3][30] ),
    .S0(_04477_),
    .S1(_04478_),
    .X(_05162_));
 sky130_fd_sc_hd__mux2_1 _10457_ (.A0(_05161_),
    .A1(_05162_),
    .S(_04121_),
    .X(_05163_));
 sky130_fd_sc_hd__mux4_1 _10458_ (.A0(\cpuregs.regs[12][30] ),
    .A1(\cpuregs.regs[13][30] ),
    .A2(\cpuregs.regs[14][30] ),
    .A3(\cpuregs.regs[15][30] ),
    .S0(_04487_),
    .S1(_04059_),
    .X(_05164_));
 sky130_fd_sc_hd__mux4_1 _10459_ (.A0(\cpuregs.regs[8][30] ),
    .A1(\cpuregs.regs[9][30] ),
    .A2(\cpuregs.regs[10][30] ),
    .A3(\cpuregs.regs[11][30] ),
    .S0(_04280_),
    .S1(_04059_),
    .X(_05165_));
 sky130_fd_sc_hd__mux2_1 _10460_ (.A0(_05164_),
    .A1(_05165_),
    .S(_04064_),
    .X(_05166_));
 sky130_fd_sc_hd__a21o_1 _10461_ (.A1(_04053_),
    .A2(_05166_),
    .B1(_04095_),
    .X(_05167_));
 sky130_fd_sc_hd__a21oi_1 _10462_ (.A1(_04070_),
    .A2(_05163_),
    .B1(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__a211o_2 _10463_ (.A1(_05156_),
    .A2(_05160_),
    .B1(net300),
    .C1(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__inv_2 _10464_ (.A(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__a221o_1 _10465_ (.A1(\irq_mask[30] ),
    .A2(_04308_),
    .B1(\timer[30] ),
    .B2(_04023_),
    .C1(_04026_),
    .X(_05171_));
 sky130_fd_sc_hd__a21o_1 _10466_ (.A1(_04271_),
    .A2(_05170_),
    .B1(_05171_),
    .X(_05172_));
 sky130_fd_sc_hd__o211a_1 _10467_ (.A1(_04268_),
    .A2(_05152_),
    .B1(_05172_),
    .C1(_03302_),
    .X(_05173_));
 sky130_fd_sc_hd__clkbuf_4 _10468_ (.A(net90),
    .X(_05174_));
 sky130_fd_sc_hd__a21o_1 _10469_ (.A1(net56),
    .A2(_04745_),
    .B1(_04666_),
    .X(_05175_));
 sky130_fd_sc_hd__a221o_1 _10470_ (.A1(_04046_),
    .A2(_05174_),
    .B1(_04752_),
    .B2(_05175_),
    .C1(_04266_),
    .X(_05176_));
 sky130_fd_sc_hd__o22a_1 _10471_ (.A1(\irq_pending[30] ),
    .A2(_04007_),
    .B1(_05173_),
    .B2(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__a21o_1 _10472_ (.A1(_04391_),
    .A2(_05150_),
    .B1(_05177_),
    .X(_08392_));
 sky130_fd_sc_hd__a31o_1 _10473_ (.A1(_05113_),
    .A2(_05117_),
    .A3(_05118_),
    .B1(_05148_),
    .X(_05178_));
 sky130_fd_sc_hd__xnor2_1 _10474_ (.A(\reg_pc[31] ),
    .B(\decoded_imm[31] ),
    .Y(_05179_));
 sky130_fd_sc_hd__a21oi_1 _10475_ (.A1(_05146_),
    .A2(_05178_),
    .B1(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__a31o_1 _10476_ (.A1(_05146_),
    .A2(_05178_),
    .A3(_05179_),
    .B1(_04156_),
    .X(_05181_));
 sky130_fd_sc_hd__a22o_1 _10477_ (.A1(\count_instr[63] ),
    .A2(_04104_),
    .B1(_04105_),
    .B2(\count_cycle[63] ),
    .X(_05182_));
 sky130_fd_sc_hd__a221o_1 _10478_ (.A1(\count_instr[31] ),
    .A2(_04012_),
    .B1(\count_cycle[31] ),
    .B2(_04165_),
    .C1(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__mux4_1 _10479_ (.A0(\cpuregs.regs[20][31] ),
    .A1(\cpuregs.regs[21][31] ),
    .A2(\cpuregs.regs[22][31] ),
    .A3(\cpuregs.regs[23][31] ),
    .S0(_04291_),
    .S1(_04292_),
    .X(_05184_));
 sky130_fd_sc_hd__mux4_1 _10480_ (.A0(\cpuregs.regs[16][31] ),
    .A1(\cpuregs.regs[17][31] ),
    .A2(\cpuregs.regs[18][31] ),
    .A3(\cpuregs.regs[19][31] ),
    .S0(_04291_),
    .S1(_04292_),
    .X(_05185_));
 sky130_fd_sc_hd__mux2_1 _10481_ (.A0(_05184_),
    .A1(_05185_),
    .S(_04223_),
    .X(_05186_));
 sky130_fd_sc_hd__nand2_1 _10482_ (.A(_04289_),
    .B(_05186_),
    .Y(_05187_));
 sky130_fd_sc_hd__mux4_1 _10483_ (.A0(\cpuregs.regs[28][31] ),
    .A1(\cpuregs.regs[29][31] ),
    .A2(\cpuregs.regs[30][31] ),
    .A3(\cpuregs.regs[31][31] ),
    .S0(_04274_),
    .S1(_04317_),
    .X(_05188_));
 sky130_fd_sc_hd__mux4_1 _10484_ (.A0(\cpuregs.regs[24][31] ),
    .A1(\cpuregs.regs[25][31] ),
    .A2(\cpuregs.regs[26][31] ),
    .A3(\cpuregs.regs[27][31] ),
    .S0(_04274_),
    .S1(_04317_),
    .X(_05189_));
 sky130_fd_sc_hd__mux2_1 _10485_ (.A0(_05188_),
    .A1(_05189_),
    .S(_04321_),
    .X(_05190_));
 sky130_fd_sc_hd__a21oi_1 _10486_ (.A1(_04206_),
    .A2(_05190_),
    .B1(_04225_),
    .Y(_05191_));
 sky130_fd_sc_hd__mux4_1 _10487_ (.A0(\cpuregs.regs[4][31] ),
    .A1(\cpuregs.regs[5][31] ),
    .A2(\cpuregs.regs[6][31] ),
    .A3(\cpuregs.regs[7][31] ),
    .S0(_04325_),
    .S1(_04277_),
    .X(_05192_));
 sky130_fd_sc_hd__mux4_1 _10488_ (.A0(\cpuregs.regs[0][31] ),
    .A1(\cpuregs.regs[1][31] ),
    .A2(\cpuregs.regs[2][31] ),
    .A3(\cpuregs.regs[3][31] ),
    .S0(_04325_),
    .S1(_04277_),
    .X(_05193_));
 sky130_fd_sc_hd__mux2_1 _10489_ (.A0(_05192_),
    .A1(_05193_),
    .S(_04223_),
    .X(_05194_));
 sky130_fd_sc_hd__mux4_1 _10490_ (.A0(\cpuregs.regs[12][31] ),
    .A1(\cpuregs.regs[13][31] ),
    .A2(\cpuregs.regs[14][31] ),
    .A3(\cpuregs.regs[15][31] ),
    .S0(_04329_),
    .S1(_04218_),
    .X(_05195_));
 sky130_fd_sc_hd__mux4_1 _10491_ (.A0(\cpuregs.regs[8][31] ),
    .A1(\cpuregs.regs[9][31] ),
    .A2(\cpuregs.regs[10][31] ),
    .A3(\cpuregs.regs[11][31] ),
    .S0(_04329_),
    .S1(_04218_),
    .X(_05196_));
 sky130_fd_sc_hd__mux2_1 _10492_ (.A0(_05195_),
    .A1(_05196_),
    .S(_04222_),
    .X(_05197_));
 sky130_fd_sc_hd__a21o_1 _10493_ (.A1(_04328_),
    .A2(_05197_),
    .B1(_04237_),
    .X(_05198_));
 sky130_fd_sc_hd__a21oi_1 _10494_ (.A1(_04289_),
    .A2(_05194_),
    .B1(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__a211o_4 _10495_ (.A1(_05187_),
    .A2(_05191_),
    .B1(_04100_),
    .C1(_05199_),
    .X(_05200_));
 sky130_fd_sc_hd__inv_2 _10496_ (.A(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__a221o_1 _10497_ (.A1(\irq_mask[31] ),
    .A2(_04021_),
    .B1(\timer[31] ),
    .B2(_04023_),
    .C1(_04188_),
    .X(_05202_));
 sky130_fd_sc_hd__a21o_1 _10498_ (.A1(_04271_),
    .A2(_05201_),
    .B1(_05202_),
    .X(_05203_));
 sky130_fd_sc_hd__o211a_1 _10499_ (.A1(_04010_),
    .A2(_05183_),
    .B1(_05203_),
    .C1(_03302_),
    .X(_05204_));
 sky130_fd_sc_hd__buf_4 _10500_ (.A(net91),
    .X(_05205_));
 sky130_fd_sc_hd__a21o_1 _10501_ (.A1(net57),
    .A2(_04811_),
    .B1(_04667_),
    .X(_05206_));
 sky130_fd_sc_hd__a221o_1 _10502_ (.A1(_03680_),
    .A2(_05205_),
    .B1(_04752_),
    .B2(_05206_),
    .C1(_04202_),
    .X(_05207_));
 sky130_fd_sc_hd__o22ai_1 _10503_ (.A1(\irq_pending[31] ),
    .A2(_04007_),
    .B1(_05204_),
    .B2(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__o21ai_1 _10504_ (.A1(_05180_),
    .A2(_05181_),
    .B1(_05208_),
    .Y(_08393_));
 sky130_fd_sc_hd__nor4_2 _10505_ (.A(instr_sra),
    .B(instr_srl),
    .C(instr_srai),
    .D(instr_srli),
    .Y(_05209_));
 sky130_fd_sc_hd__nor2_2 _10506_ (.A(instr_sll),
    .B(instr_slli),
    .Y(_05210_));
 sky130_fd_sc_hd__nand2_1 _10507_ (.A(_05209_),
    .B(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__or2_1 _10508_ (.A(instr_and),
    .B(instr_andi),
    .X(_05212_));
 sky130_fd_sc_hd__or2_2 _10509_ (.A(instr_or),
    .B(instr_ori),
    .X(_05213_));
 sky130_fd_sc_hd__or2_1 _10510_ (.A(instr_xor),
    .B(instr_xori),
    .X(_05214_));
 sky130_fd_sc_hd__clkbuf_4 _10511_ (.A(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__or4_1 _10512_ (.A(is_compare),
    .B(_05212_),
    .C(_05213_),
    .D(_05215_),
    .X(_05216_));
 sky130_fd_sc_hd__or2_1 _10513_ (.A(_05211_),
    .B(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__clkbuf_4 _10514_ (.A(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__clkbuf_8 _10515_ (.A(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__clkbuf_4 _10516_ (.A(_05215_),
    .X(_05220_));
 sky130_fd_sc_hd__nor2_4 _10517_ (.A(instr_or),
    .B(instr_ori),
    .Y(_05221_));
 sky130_fd_sc_hd__clkbuf_4 _10518_ (.A(_05212_),
    .X(_05222_));
 sky130_fd_sc_hd__a2bb2o_1 _10519_ (.A1_N(_03610_),
    .A2_N(_05221_),
    .B1(_05222_),
    .B2(_03611_),
    .X(_05223_));
 sky130_fd_sc_hd__a21o_1 _10520_ (.A1(_03612_),
    .A2(_05220_),
    .B1(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__inv_2 _10521_ (.A(_05218_),
    .Y(_05225_));
 sky130_fd_sc_hd__clkbuf_4 _10522_ (.A(net125),
    .X(_05226_));
 sky130_fd_sc_hd__buf_4 _10523_ (.A(_05209_),
    .X(_05227_));
 sky130_fd_sc_hd__nor2_4 _10524_ (.A(_05226_),
    .B(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__clkbuf_4 _10525_ (.A(_03609_),
    .X(_05229_));
 sky130_fd_sc_hd__buf_4 _10526_ (.A(_05229_),
    .X(_05230_));
 sky130_fd_sc_hd__clkbuf_4 _10527_ (.A(net110),
    .X(_05231_));
 sky130_fd_sc_hd__clkbuf_4 _10528_ (.A(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__mux4_1 _10529_ (.A0(_04419_),
    .A1(_04456_),
    .A2(_04466_),
    .A3(_04532_),
    .S0(_05230_),
    .S1(_05232_),
    .X(_05233_));
 sky130_fd_sc_hd__mux4_1 _10530_ (.A0(_04566_),
    .A1(_04602_),
    .A2(_04611_),
    .A3(_04642_),
    .S0(_05230_),
    .S1(_05232_),
    .X(_05234_));
 sky130_fd_sc_hd__clkbuf_4 _10531_ (.A(_05231_),
    .X(_05235_));
 sky130_fd_sc_hd__clkbuf_4 _10532_ (.A(_03609_),
    .X(_05236_));
 sky130_fd_sc_hd__clkbuf_4 _10533_ (.A(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__mux4_1 _10534_ (.A0(_04036_),
    .A1(_04160_),
    .A2(_04039_),
    .A3(_04198_),
    .S0(_05235_),
    .S1(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__buf_4 _10535_ (.A(_05231_),
    .X(_05239_));
 sky130_fd_sc_hd__clkbuf_4 _10536_ (.A(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__mux4_1 _10537_ (.A0(_04251_),
    .A1(_04262_),
    .A2(_04342_),
    .A3(_04360_),
    .S0(_05230_),
    .S1(_05240_),
    .X(_05241_));
 sky130_fd_sc_hd__clkbuf_4 _10538_ (.A(net121),
    .X(_05242_));
 sky130_fd_sc_hd__clkbuf_4 _10539_ (.A(_05242_),
    .X(_05243_));
 sky130_fd_sc_hd__buf_4 _10540_ (.A(_03531_),
    .X(_05244_));
 sky130_fd_sc_hd__mux4_1 _10541_ (.A0(_05233_),
    .A1(_05234_),
    .A2(_05238_),
    .A3(_05241_),
    .S0(_05243_),
    .S1(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__clkbuf_4 _10542_ (.A(_05242_),
    .X(_05246_));
 sky130_fd_sc_hd__or3_1 _10543_ (.A(_04033_),
    .B(_05230_),
    .C(_05235_),
    .X(_05247_));
 sky130_fd_sc_hd__or2_1 _10544_ (.A(_05246_),
    .B(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__inv_2 _10545_ (.A(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__or2_2 _10546_ (.A(_05226_),
    .B(_05210_),
    .X(_05250_));
 sky130_fd_sc_hd__nor2_4 _10547_ (.A(_03530_),
    .B(_05250_),
    .Y(_05251_));
 sky130_fd_sc_hd__a22o_1 _10548_ (.A1(_05228_),
    .A2(_05245_),
    .B1(_05249_),
    .B2(_05251_),
    .X(_05252_));
 sky130_fd_sc_hd__or3_1 _10549_ (.A(_05224_),
    .B(_05225_),
    .C(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__clkbuf_4 _10550_ (.A(_05226_),
    .X(_05254_));
 sky130_fd_sc_hd__clkbuf_8 _10551_ (.A(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__or4_1 _10552_ (.A(instr_sra),
    .B(instr_srl),
    .C(instr_srai),
    .D(instr_srli),
    .X(_05256_));
 sky130_fd_sc_hd__buf_2 _10553_ (.A(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__buf_2 _10554_ (.A(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__clkbuf_4 _10555_ (.A(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__buf_4 _10556_ (.A(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__buf_4 _10557_ (.A(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__mux2_1 _10558_ (.A0(net74),
    .A1(_04744_),
    .S(_05229_),
    .X(_05262_));
 sky130_fd_sc_hd__clkbuf_4 _10559_ (.A(_03609_),
    .X(_05263_));
 sky130_fd_sc_hd__buf_4 _10560_ (.A(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__mux2_1 _10561_ (.A0(_04754_),
    .A1(_04810_),
    .S(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__buf_4 _10562_ (.A(_05235_),
    .X(_05266_));
 sky130_fd_sc_hd__mux2_1 _10563_ (.A0(_05262_),
    .A1(_05265_),
    .S(_05266_),
    .X(_05267_));
 sky130_fd_sc_hd__mux2_1 _10564_ (.A0(_04848_),
    .A1(_04880_),
    .S(_05264_),
    .X(_05268_));
 sky130_fd_sc_hd__mux2_1 _10565_ (.A0(net81),
    .A1(_04945_),
    .S(_05236_),
    .X(_05269_));
 sky130_fd_sc_hd__mux2_1 _10566_ (.A0(_05268_),
    .A1(_05269_),
    .S(_05266_),
    .X(_05270_));
 sky130_fd_sc_hd__mux2_1 _10567_ (.A0(_04959_),
    .A1(_05013_),
    .S(_05236_),
    .X(_05271_));
 sky130_fd_sc_hd__mux2_1 _10568_ (.A0(_05044_),
    .A1(_05076_),
    .S(_05263_),
    .X(_05272_));
 sky130_fd_sc_hd__mux2_1 _10569_ (.A0(_05271_),
    .A1(_05272_),
    .S(_05240_),
    .X(_05273_));
 sky130_fd_sc_hd__mux2_1 _10570_ (.A0(net87),
    .A1(net88),
    .S(_05263_),
    .X(_05274_));
 sky130_fd_sc_hd__mux2_1 _10571_ (.A0(net90),
    .A1(_05205_),
    .S(_05229_),
    .X(_05275_));
 sky130_fd_sc_hd__mux2_1 _10572_ (.A0(_05274_),
    .A1(_05275_),
    .S(_05240_),
    .X(_05276_));
 sky130_fd_sc_hd__buf_4 _10573_ (.A(_05243_),
    .X(_05277_));
 sky130_fd_sc_hd__clkbuf_4 _10574_ (.A(_03530_),
    .X(_05278_));
 sky130_fd_sc_hd__mux4_2 _10575_ (.A0(_05267_),
    .A1(_05270_),
    .A2(_05273_),
    .A3(_05276_),
    .S0(_05277_),
    .S1(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__a32o_1 _10576_ (.A1(_05255_),
    .A2(_05261_),
    .A3(_05279_),
    .B1(is_compare),
    .B2(_03630_),
    .X(_05280_));
 sky130_fd_sc_hd__o22a_1 _10577_ (.A1(_03612_),
    .A2(_05219_),
    .B1(_05253_),
    .B2(_05280_),
    .X(\alu_out[0] ));
 sky130_fd_sc_hd__clkbuf_4 _10578_ (.A(_05251_),
    .X(_05281_));
 sky130_fd_sc_hd__mux2_1 _10579_ (.A0(_03242_),
    .A1(_04036_),
    .S(_03609_),
    .X(_05282_));
 sky130_fd_sc_hd__or2b_1 _10580_ (.A(_05231_),
    .B_N(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__or2_1 _10581_ (.A(_05242_),
    .B(_05283_),
    .X(_05284_));
 sky130_fd_sc_hd__inv_2 _10582_ (.A(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__clkbuf_8 _10583_ (.A(_05266_),
    .X(_05286_));
 sky130_fd_sc_hd__clkbuf_4 _10584_ (.A(_05244_),
    .X(_05287_));
 sky130_fd_sc_hd__clkbuf_4 _10585_ (.A(_05287_),
    .X(_05288_));
 sky130_fd_sc_hd__mux4_1 _10586_ (.A0(net98),
    .A1(net68),
    .A2(net69),
    .A3(net70),
    .S0(_05229_),
    .S1(_05239_),
    .X(_05289_));
 sky130_fd_sc_hd__mux4_1 _10587_ (.A0(net71),
    .A1(net72),
    .A2(net73),
    .A3(_04708_),
    .S0(_05229_),
    .S1(_05239_),
    .X(_05290_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(_05289_),
    .A1(_05290_),
    .S(_05242_),
    .X(_05291_));
 sky130_fd_sc_hd__clkbuf_4 _10589_ (.A(_03530_),
    .X(_05292_));
 sky130_fd_sc_hd__mux4_1 _10590_ (.A0(_04039_),
    .A1(_04198_),
    .A2(_04160_),
    .A3(_04251_),
    .S0(_05239_),
    .S1(_05237_),
    .X(_05293_));
 sky130_fd_sc_hd__mux4_1 _10591_ (.A0(_03524_),
    .A1(net95),
    .A2(_03518_),
    .A3(_03510_),
    .S0(_05264_),
    .S1(_05235_),
    .X(_05294_));
 sky130_fd_sc_hd__clkbuf_4 _10592_ (.A(_05242_),
    .X(_05295_));
 sky130_fd_sc_hd__mux2_1 _10593_ (.A0(_05293_),
    .A1(_05294_),
    .S(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__or2_1 _10594_ (.A(_05292_),
    .B(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__clkbuf_4 _10595_ (.A(_05228_),
    .X(_05298_));
 sky130_fd_sc_hd__o211a_1 _10596_ (.A1(_05288_),
    .A2(_05291_),
    .B1(_05297_),
    .C1(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__or2_2 _10597_ (.A(_03242_),
    .B(_05231_),
    .X(_05300_));
 sky130_fd_sc_hd__clkbuf_4 _10598_ (.A(_05213_),
    .X(_05301_));
 sky130_fd_sc_hd__a22o_1 _10599_ (.A1(_05300_),
    .A2(_05301_),
    .B1(_05220_),
    .B2(_03535_),
    .X(_05302_));
 sky130_fd_sc_hd__a311o_1 _10600_ (.A1(_04040_),
    .A2(_05286_),
    .A3(_05222_),
    .B1(_05299_),
    .C1(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__mux2_1 _10601_ (.A0(_04744_),
    .A1(net76),
    .S(_05229_),
    .X(_05304_));
 sky130_fd_sc_hd__mux2_1 _10602_ (.A0(net77),
    .A1(net79),
    .S(_05263_),
    .X(_05305_));
 sky130_fd_sc_hd__mux2_1 _10603_ (.A0(_05304_),
    .A1(_05305_),
    .S(_05232_),
    .X(_05306_));
 sky130_fd_sc_hd__mux2_1 _10604_ (.A0(_04880_),
    .A1(net81),
    .S(_05263_),
    .X(_05307_));
 sky130_fd_sc_hd__mux2_1 _10605_ (.A0(net82),
    .A1(net83),
    .S(_05263_),
    .X(_05308_));
 sky130_fd_sc_hd__clkbuf_4 _10606_ (.A(_05231_),
    .X(_05309_));
 sky130_fd_sc_hd__mux2_1 _10607_ (.A0(_05307_),
    .A1(_05308_),
    .S(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__mux2_1 _10608_ (.A0(_05306_),
    .A1(_05310_),
    .S(_05246_),
    .X(_05311_));
 sky130_fd_sc_hd__mux2_1 _10609_ (.A0(_05013_),
    .A1(net85),
    .S(_05263_),
    .X(_05312_));
 sky130_fd_sc_hd__mux2_1 _10610_ (.A0(net86),
    .A1(net87),
    .S(_05263_),
    .X(_05313_));
 sky130_fd_sc_hd__mux2_1 _10611_ (.A0(_05312_),
    .A1(_05313_),
    .S(_05309_),
    .X(_05314_));
 sky130_fd_sc_hd__mux2_1 _10612_ (.A0(net88),
    .A1(net90),
    .S(_05263_),
    .X(_05315_));
 sky130_fd_sc_hd__o21ai_2 _10613_ (.A1(instr_sra),
    .A2(instr_srai),
    .B1(_05205_),
    .Y(_05316_));
 sky130_fd_sc_hd__or2b_1 _10614_ (.A(_05263_),
    .B_N(_05205_),
    .X(_05317_));
 sky130_fd_sc_hd__nand2_1 _10615_ (.A(_05316_),
    .B(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__mux2_1 _10616_ (.A0(_05315_),
    .A1(_05318_),
    .S(_05309_),
    .X(_05319_));
 sky130_fd_sc_hd__mux2_1 _10617_ (.A0(_05314_),
    .A1(_05319_),
    .S(_05295_),
    .X(_05320_));
 sky130_fd_sc_hd__mux2_1 _10618_ (.A0(_05311_),
    .A1(_05320_),
    .S(_05292_),
    .X(_05321_));
 sky130_fd_sc_hd__inv_2 _10619_ (.A(instr_sub),
    .Y(_05322_));
 sky130_fd_sc_hd__buf_4 _10620_ (.A(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__clkbuf_8 _10621_ (.A(_05230_),
    .X(_05324_));
 sky130_fd_sc_hd__and2_1 _10622_ (.A(_05323_),
    .B(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__xnor2_1 _10623_ (.A(_03535_),
    .B(_03536_),
    .Y(_05326_));
 sky130_fd_sc_hd__xnor2_1 _10624_ (.A(_05325_),
    .B(_05326_),
    .Y(_05327_));
 sky130_fd_sc_hd__a32o_1 _10625_ (.A1(_05255_),
    .A2(_05261_),
    .A3(_05321_),
    .B1(_05327_),
    .B2(_05225_),
    .X(_05328_));
 sky130_fd_sc_hd__a211o_1 _10626_ (.A1(_05281_),
    .A2(_05285_),
    .B1(_05303_),
    .C1(_05328_),
    .X(\alu_out[1] ));
 sky130_fd_sc_hd__mux2_1 _10627_ (.A0(_05265_),
    .A1(_05268_),
    .S(_05240_),
    .X(_05329_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(_05269_),
    .A1(_05271_),
    .S(_05232_),
    .X(_05330_));
 sky130_fd_sc_hd__clkbuf_4 _10629_ (.A(_05295_),
    .X(_05331_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(_05329_),
    .A1(_05330_),
    .S(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__mux2_1 _10631_ (.A0(_05272_),
    .A1(_05274_),
    .S(_05309_),
    .X(_05333_));
 sky130_fd_sc_hd__o21a_4 _10632_ (.A1(instr_sra),
    .A2(instr_srai),
    .B1(_05205_),
    .X(_05334_));
 sky130_fd_sc_hd__mux2_1 _10633_ (.A0(_05275_),
    .A1(_05334_),
    .S(_05309_),
    .X(_05335_));
 sky130_fd_sc_hd__mux2_1 _10634_ (.A0(_05333_),
    .A1(_05335_),
    .S(_05295_),
    .X(_05336_));
 sky130_fd_sc_hd__mux2_1 _10635_ (.A0(_05332_),
    .A1(_05336_),
    .S(_05278_),
    .X(_05337_));
 sky130_fd_sc_hd__a22o_1 _10636_ (.A1(net67),
    .A2(net99),
    .B1(_05231_),
    .B2(_03242_),
    .X(_05338_));
 sky130_fd_sc_hd__nand2_1 _10637_ (.A(_05300_),
    .B(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__mux2_1 _10638_ (.A0(_03538_),
    .A1(_05339_),
    .S(_05323_),
    .X(_05340_));
 sky130_fd_sc_hd__xor2_1 _10639_ (.A(_03534_),
    .B(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__mux2_1 _10640_ (.A0(net89),
    .A1(_03242_),
    .S(_03609_),
    .X(_05342_));
 sky130_fd_sc_hd__o21ai_1 _10641_ (.A1(_04033_),
    .A2(_05237_),
    .B1(_05232_),
    .Y(_05343_));
 sky130_fd_sc_hd__o21ai_1 _10642_ (.A1(_05240_),
    .A2(_05342_),
    .B1(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__nor2_1 _10643_ (.A(_05331_),
    .B(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__mux4_1 _10644_ (.A0(_04466_),
    .A1(_04532_),
    .A2(_04566_),
    .A3(_04602_),
    .S0(_05264_),
    .S1(_05232_),
    .X(_05346_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(net72),
    .A1(net73),
    .S(_05229_),
    .X(_05347_));
 sky130_fd_sc_hd__mux2_1 _10646_ (.A0(_05347_),
    .A1(_05262_),
    .S(_05235_),
    .X(_05348_));
 sky130_fd_sc_hd__mux2_1 _10647_ (.A0(_05346_),
    .A1(_05348_),
    .S(_05246_),
    .X(_05349_));
 sky130_fd_sc_hd__mux4_1 _10648_ (.A0(_04160_),
    .A1(_04251_),
    .A2(_04198_),
    .A3(_03524_),
    .S0(_05239_),
    .S1(_05237_),
    .X(_05350_));
 sky130_fd_sc_hd__mux4_1 _10649_ (.A0(_04342_),
    .A1(_04419_),
    .A2(_03518_),
    .A3(_04456_),
    .S0(_05239_),
    .S1(_05237_),
    .X(_05351_));
 sky130_fd_sc_hd__mux2_1 _10650_ (.A0(_05350_),
    .A1(_05351_),
    .S(_05246_),
    .X(_05352_));
 sky130_fd_sc_hd__mux2_1 _10651_ (.A0(_05349_),
    .A1(_05352_),
    .S(_05287_),
    .X(_05353_));
 sky130_fd_sc_hd__a22o_1 _10652_ (.A1(_05281_),
    .A2(_05345_),
    .B1(_05353_),
    .B2(_05298_),
    .X(_05354_));
 sky130_fd_sc_hd__and2_1 _10653_ (.A(net121),
    .B(net89),
    .X(_05355_));
 sky130_fd_sc_hd__nor2_2 _10654_ (.A(instr_xor),
    .B(instr_xori),
    .Y(_05356_));
 sky130_fd_sc_hd__clkbuf_4 _10655_ (.A(_05356_),
    .X(_05357_));
 sky130_fd_sc_hd__nor2_1 _10656_ (.A(_03534_),
    .B(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__a221o_1 _10657_ (.A1(_05355_),
    .A2(_05222_),
    .B1(_05301_),
    .B2(_03532_),
    .C1(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__a211o_1 _10658_ (.A1(_05225_),
    .A2(_05341_),
    .B1(_05354_),
    .C1(_05359_),
    .X(_05360_));
 sky130_fd_sc_hd__a31o_1 _10659_ (.A1(_05255_),
    .A2(_05261_),
    .A3(_05337_),
    .B1(_05360_),
    .X(\alu_out[2] ));
 sky130_fd_sc_hd__clkbuf_4 _10660_ (.A(_05225_),
    .X(_05361_));
 sky130_fd_sc_hd__a31o_1 _10661_ (.A1(_05300_),
    .A2(_03532_),
    .A3(_05338_),
    .B1(_05355_),
    .X(_05362_));
 sky130_fd_sc_hd__buf_4 _10662_ (.A(_05323_),
    .X(_05363_));
 sky130_fd_sc_hd__mux2_1 _10663_ (.A0(_03540_),
    .A1(_05362_),
    .S(_05363_),
    .X(_05364_));
 sky130_fd_sc_hd__or2_1 _10664_ (.A(_03608_),
    .B(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__nand2_1 _10665_ (.A(_03608_),
    .B(_05364_),
    .Y(_05366_));
 sky130_fd_sc_hd__buf_4 _10666_ (.A(_05221_),
    .X(_05367_));
 sky130_fd_sc_hd__nor2_1 _10667_ (.A(_03606_),
    .B(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__a221o_1 _10668_ (.A1(_03607_),
    .A2(_05222_),
    .B1(_05220_),
    .B2(_03608_),
    .C1(_05368_),
    .X(_05369_));
 sky130_fd_sc_hd__mux4_2 _10669_ (.A0(_04532_),
    .A1(_04566_),
    .A2(_04602_),
    .A3(_04611_),
    .S0(_05230_),
    .S1(_05240_),
    .X(_05370_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(net73),
    .A1(net74),
    .S(_05229_),
    .X(_05371_));
 sky130_fd_sc_hd__mux2_1 _10671_ (.A0(_05371_),
    .A1(_05304_),
    .S(_05309_),
    .X(_05372_));
 sky130_fd_sc_hd__mux4_1 _10672_ (.A0(_04198_),
    .A1(_04262_),
    .A2(_04251_),
    .A3(_04342_),
    .S0(_05235_),
    .S1(_05324_),
    .X(_05373_));
 sky130_fd_sc_hd__mux4_1 _10673_ (.A0(_04360_),
    .A1(_04456_),
    .A2(_04419_),
    .A3(_04466_),
    .S0(_05235_),
    .S1(_05237_),
    .X(_05374_));
 sky130_fd_sc_hd__mux4_1 _10674_ (.A0(_05370_),
    .A1(_05372_),
    .A2(_05373_),
    .A3(_05374_),
    .S0(_05243_),
    .S1(_05244_),
    .X(_05375_));
 sky130_fd_sc_hd__mux4_1 _10675_ (.A0(_04198_),
    .A1(_04160_),
    .A2(_04039_),
    .A3(_04036_),
    .S0(_05236_),
    .S1(_05239_),
    .X(_05376_));
 sky130_fd_sc_hd__and2b_1 _10676_ (.A_N(_05243_),
    .B(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__a22o_1 _10677_ (.A1(_05228_),
    .A2(_05375_),
    .B1(_05377_),
    .B2(_05251_),
    .X(_05378_));
 sky130_fd_sc_hd__mux2_1 _10678_ (.A0(_05305_),
    .A1(_05307_),
    .S(_05239_),
    .X(_05379_));
 sky130_fd_sc_hd__mux2_1 _10679_ (.A0(_05308_),
    .A1(_05312_),
    .S(_05239_),
    .X(_05380_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(_05379_),
    .A1(_05380_),
    .S(_05242_),
    .X(_05381_));
 sky130_fd_sc_hd__mux2_1 _10681_ (.A0(_05313_),
    .A1(_05315_),
    .S(_05239_),
    .X(_05382_));
 sky130_fd_sc_hd__o21ai_1 _10682_ (.A1(_05232_),
    .A2(_05317_),
    .B1(_05316_),
    .Y(_05383_));
 sky130_fd_sc_hd__mux2_1 _10683_ (.A0(_05382_),
    .A1(_05383_),
    .S(_05242_),
    .X(_05384_));
 sky130_fd_sc_hd__mux2_1 _10684_ (.A0(_05381_),
    .A1(_05384_),
    .S(_03530_),
    .X(_05385_));
 sky130_fd_sc_hd__and3_1 _10685_ (.A(_05254_),
    .B(_05260_),
    .C(_05385_),
    .X(_05386_));
 sky130_fd_sc_hd__or3_1 _10686_ (.A(_05369_),
    .B(_05378_),
    .C(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__a31o_2 _10687_ (.A1(_05361_),
    .A2(_05365_),
    .A3(_05366_),
    .B1(_05387_),
    .X(\alu_out[3] ));
 sky130_fd_sc_hd__a311oi_2 _10688_ (.A1(_05300_),
    .A2(_03532_),
    .A3(_05338_),
    .B1(_05355_),
    .C1(_03607_),
    .Y(_05388_));
 sky130_fd_sc_hd__or2_1 _10689_ (.A(_03606_),
    .B(_05388_),
    .X(_05389_));
 sky130_fd_sc_hd__buf_4 _10690_ (.A(_05323_),
    .X(_05390_));
 sky130_fd_sc_hd__mux2_1 _10691_ (.A0(_03542_),
    .A1(_05389_),
    .S(_05390_),
    .X(_05391_));
 sky130_fd_sc_hd__nand2_1 _10692_ (.A(_03529_),
    .B(_05391_),
    .Y(_05392_));
 sky130_fd_sc_hd__or2_1 _10693_ (.A(_03529_),
    .B(_05391_),
    .X(_05393_));
 sky130_fd_sc_hd__mux4_2 _10694_ (.A0(_05270_),
    .A1(_05273_),
    .A2(_05276_),
    .A3(_05334_),
    .S0(_05277_),
    .S1(_05278_),
    .X(_05394_));
 sky130_fd_sc_hd__clkbuf_4 _10695_ (.A(_05246_),
    .X(_05395_));
 sky130_fd_sc_hd__mux4_1 _10696_ (.A0(_05234_),
    .A1(_05267_),
    .A2(_05241_),
    .A3(_05233_),
    .S0(_05395_),
    .S1(_05287_),
    .X(_05396_));
 sky130_fd_sc_hd__nor2_2 _10697_ (.A(instr_and),
    .B(instr_andi),
    .Y(_05397_));
 sky130_fd_sc_hd__clkbuf_4 _10698_ (.A(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__nor2_2 _10699_ (.A(_05226_),
    .B(_05210_),
    .Y(_05399_));
 sky130_fd_sc_hd__nand2_1 _10700_ (.A(_05244_),
    .B(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(net93),
    .A1(net92),
    .S(_03609_),
    .X(_05401_));
 sky130_fd_sc_hd__mux2_1 _10702_ (.A0(_05401_),
    .A1(_05342_),
    .S(_05231_),
    .X(_05402_));
 sky130_fd_sc_hd__inv_2 _10703_ (.A(_05402_),
    .Y(_05403_));
 sky130_fd_sc_hd__mux2_2 _10704_ (.A0(_05403_),
    .A1(_05247_),
    .S(_05246_),
    .X(_05404_));
 sky130_fd_sc_hd__o22a_1 _10705_ (.A1(_03527_),
    .A2(_05221_),
    .B1(_05356_),
    .B2(_03529_),
    .X(_05405_));
 sky130_fd_sc_hd__o221a_1 _10706_ (.A1(_03528_),
    .A2(_05398_),
    .B1(_05400_),
    .B2(_05404_),
    .C1(_05405_),
    .X(_05406_));
 sky130_fd_sc_hd__a21bo_1 _10707_ (.A1(_05298_),
    .A2(_05396_),
    .B1_N(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__a31o_1 _10708_ (.A1(_05255_),
    .A2(_05261_),
    .A3(_05394_),
    .B1(_05407_),
    .X(_05408_));
 sky130_fd_sc_hd__a31o_1 _10709_ (.A1(_05361_),
    .A2(_05392_),
    .A3(_05393_),
    .B1(_05408_),
    .X(\alu_out[4] ));
 sky130_fd_sc_hd__o21ai_1 _10710_ (.A1(_03527_),
    .A2(_05389_),
    .B1(_03528_),
    .Y(_05409_));
 sky130_fd_sc_hd__mux2_1 _10711_ (.A0(_03544_),
    .A1(_05409_),
    .S(_05390_),
    .X(_05410_));
 sky130_fd_sc_hd__or2_1 _10712_ (.A(_03526_),
    .B(_05410_),
    .X(_05411_));
 sky130_fd_sc_hd__nand2_1 _10713_ (.A(_03526_),
    .B(_05410_),
    .Y(_05412_));
 sky130_fd_sc_hd__buf_6 _10714_ (.A(_05331_),
    .X(_05413_));
 sky130_fd_sc_hd__buf_4 _10715_ (.A(_05292_),
    .X(_05414_));
 sky130_fd_sc_hd__mux4_1 _10716_ (.A0(_05294_),
    .A1(_05289_),
    .A2(_05290_),
    .A3(_05306_),
    .S0(_05413_),
    .S1(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__mux4_2 _10717_ (.A0(_03524_),
    .A1(net93),
    .A2(net92),
    .A3(net89),
    .S0(_03609_),
    .S1(_05231_),
    .X(_05416_));
 sky130_fd_sc_hd__inv_2 _10718_ (.A(_05416_),
    .Y(_05417_));
 sky130_fd_sc_hd__mux2_1 _10719_ (.A0(_05417_),
    .A1(_05283_),
    .S(_05295_),
    .X(_05418_));
 sky130_fd_sc_hd__nor2_1 _10720_ (.A(_05400_),
    .B(_05418_),
    .Y(_05419_));
 sky130_fd_sc_hd__a221o_1 _10721_ (.A1(_03523_),
    .A2(_05301_),
    .B1(_05215_),
    .B2(_03526_),
    .C1(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__a31o_1 _10722_ (.A1(net126),
    .A2(_04262_),
    .A3(_05222_),
    .B1(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__mux2_1 _10723_ (.A0(_05310_),
    .A1(_05314_),
    .S(_05295_),
    .X(_05422_));
 sky130_fd_sc_hd__nand2_1 _10724_ (.A(_05242_),
    .B(_05316_),
    .Y(_05423_));
 sky130_fd_sc_hd__o21a_1 _10725_ (.A1(_05243_),
    .A2(_05319_),
    .B1(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__mux2_1 _10726_ (.A0(_05422_),
    .A1(_05424_),
    .S(_03530_),
    .X(_05425_));
 sky130_fd_sc_hd__and3_1 _10727_ (.A(_05254_),
    .B(_05261_),
    .C(_05425_),
    .X(_05426_));
 sky130_fd_sc_hd__a211o_1 _10728_ (.A1(_05298_),
    .A2(_05415_),
    .B1(_05421_),
    .C1(_05426_),
    .X(_05427_));
 sky130_fd_sc_hd__a31o_1 _10729_ (.A1(_05361_),
    .A2(_05411_),
    .A3(_05412_),
    .B1(_05427_),
    .X(\alu_out[5] ));
 sky130_fd_sc_hd__inv_2 _10730_ (.A(_03523_),
    .Y(_05428_));
 sky130_fd_sc_hd__o311a_1 _10731_ (.A1(_03606_),
    .A2(_03527_),
    .A3(_05388_),
    .B1(_03528_),
    .C1(_03525_),
    .X(_05429_));
 sky130_fd_sc_hd__or2_1 _10732_ (.A(_05428_),
    .B(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__mux2_1 _10733_ (.A0(_03546_),
    .A1(_05430_),
    .S(_05363_),
    .X(_05431_));
 sky130_fd_sc_hd__nor2_1 _10734_ (.A(_03522_),
    .B(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__a21o_1 _10735_ (.A1(_03522_),
    .A2(_05431_),
    .B1(_05218_),
    .X(_05433_));
 sky130_fd_sc_hd__nand2_1 _10736_ (.A(_05226_),
    .B(_05259_),
    .Y(_05434_));
 sky130_fd_sc_hd__and2b_1 _10737_ (.A_N(_05243_),
    .B(_05330_),
    .X(_05435_));
 sky130_fd_sc_hd__a21oi_1 _10738_ (.A1(_05277_),
    .A2(_05333_),
    .B1(_05435_),
    .Y(_05436_));
 sky130_fd_sc_hd__o21a_1 _10739_ (.A1(_05246_),
    .A2(_05335_),
    .B1(_05423_),
    .X(_05437_));
 sky130_fd_sc_hd__inv_2 _10740_ (.A(_05437_),
    .Y(_05438_));
 sky130_fd_sc_hd__mux2_1 _10741_ (.A0(_05436_),
    .A1(_05438_),
    .S(_05278_),
    .X(_05439_));
 sky130_fd_sc_hd__clkbuf_4 _10742_ (.A(_05398_),
    .X(_05440_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(net95),
    .A1(_03524_),
    .S(_03609_),
    .X(_05441_));
 sky130_fd_sc_hd__mux2_1 _10744_ (.A0(_05441_),
    .A1(_05401_),
    .S(_05231_),
    .X(_05442_));
 sky130_fd_sc_hd__inv_2 _10745_ (.A(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hd__mux2_1 _10746_ (.A0(_05443_),
    .A1(_05344_),
    .S(_05246_),
    .X(_05444_));
 sky130_fd_sc_hd__o22a_1 _10747_ (.A1(_03519_),
    .A2(_05367_),
    .B1(_05356_),
    .B2(_03522_),
    .X(_05445_));
 sky130_fd_sc_hd__o221a_1 _10748_ (.A1(_03520_),
    .A2(_05440_),
    .B1(_05400_),
    .B2(_05444_),
    .C1(_05445_),
    .X(_05446_));
 sky130_fd_sc_hd__mux4_1 _10749_ (.A0(_05348_),
    .A1(_05329_),
    .A2(_05351_),
    .A3(_05346_),
    .S0(_05277_),
    .S1(_05288_),
    .X(_05447_));
 sky130_fd_sc_hd__nand2_1 _10750_ (.A(_05298_),
    .B(_05447_),
    .Y(_05448_));
 sky130_fd_sc_hd__o211a_1 _10751_ (.A1(_05434_),
    .A2(_05439_),
    .B1(_05446_),
    .C1(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__o21ai_2 _10752_ (.A1(_05432_),
    .A2(_05433_),
    .B1(_05449_),
    .Y(\alu_out[6] ));
 sky130_fd_sc_hd__a21oi_1 _10753_ (.A1(_03522_),
    .A2(_03546_),
    .B1(_03547_),
    .Y(_05450_));
 sky130_fd_sc_hd__o21ai_1 _10754_ (.A1(_03519_),
    .A2(_05430_),
    .B1(_03520_),
    .Y(_05451_));
 sky130_fd_sc_hd__mux2_1 _10755_ (.A0(_05450_),
    .A1(_05451_),
    .S(_05390_),
    .X(_05452_));
 sky130_fd_sc_hd__or2_1 _10756_ (.A(_03615_),
    .B(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__nand2_1 _10757_ (.A(_03615_),
    .B(_05452_),
    .Y(_05454_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(_05380_),
    .A1(_05382_),
    .S(_05395_),
    .X(_05455_));
 sky130_fd_sc_hd__nand2_1 _10759_ (.A(_05383_),
    .B(_05423_),
    .Y(_05456_));
 sky130_fd_sc_hd__inv_2 _10760_ (.A(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__mux2_1 _10761_ (.A0(_05455_),
    .A1(_05457_),
    .S(_05278_),
    .X(_05458_));
 sky130_fd_sc_hd__mux4_1 _10762_ (.A0(_05372_),
    .A1(_05379_),
    .A2(_05374_),
    .A3(_05370_),
    .S0(_05395_),
    .S1(_05287_),
    .X(_05459_));
 sky130_fd_sc_hd__mux4_1 _10763_ (.A0(_03518_),
    .A1(net95),
    .A2(_03524_),
    .A3(net93),
    .S0(_05236_),
    .S1(_05309_),
    .X(_05460_));
 sky130_fd_sc_hd__mux2_2 _10764_ (.A0(_05460_),
    .A1(_05376_),
    .S(_05242_),
    .X(_05461_));
 sky130_fd_sc_hd__a2bb2o_1 _10765_ (.A1_N(_03613_),
    .A2_N(_05221_),
    .B1(_05215_),
    .B2(_03615_),
    .X(_05462_));
 sky130_fd_sc_hd__a221o_1 _10766_ (.A1(_03614_),
    .A2(_05222_),
    .B1(_05251_),
    .B2(_05461_),
    .C1(_05462_),
    .X(_05463_));
 sky130_fd_sc_hd__a21o_1 _10767_ (.A1(_05298_),
    .A2(_05459_),
    .B1(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__a31o_1 _10768_ (.A1(_05255_),
    .A2(_05261_),
    .A3(_05458_),
    .B1(_05464_),
    .X(_05465_));
 sky130_fd_sc_hd__a31o_1 _10769_ (.A1(_05361_),
    .A2(_05453_),
    .A3(_05454_),
    .B1(_05465_),
    .X(\alu_out[7] ));
 sky130_fd_sc_hd__nand2_1 _10770_ (.A(net128),
    .B(net96),
    .Y(_05466_));
 sky130_fd_sc_hd__o311a_1 _10771_ (.A1(_03519_),
    .A2(_05428_),
    .A3(_05429_),
    .B1(_05466_),
    .C1(_03520_),
    .X(_05467_));
 sky130_fd_sc_hd__or2_1 _10772_ (.A(_03613_),
    .B(_05467_),
    .X(_05468_));
 sky130_fd_sc_hd__mux2_1 _10773_ (.A0(_03549_),
    .A1(_05468_),
    .S(_05363_),
    .X(_05469_));
 sky130_fd_sc_hd__xor2_1 _10774_ (.A(_03512_),
    .B(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__mux4_1 _10775_ (.A0(_05233_),
    .A1(_05234_),
    .A2(_05267_),
    .A3(_05270_),
    .S0(_05413_),
    .S1(_05414_),
    .X(_05471_));
 sky130_fd_sc_hd__nand2_1 _10776_ (.A(_03509_),
    .B(_05301_),
    .Y(_05472_));
 sky130_fd_sc_hd__o221a_1 _10777_ (.A1(_03511_),
    .A2(_05440_),
    .B1(_05357_),
    .B2(_03512_),
    .C1(_05472_),
    .X(_05473_));
 sky130_fd_sc_hd__a21bo_1 _10778_ (.A1(_05298_),
    .A2(_05471_),
    .B1_N(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(_05273_),
    .A1(_05276_),
    .S(_05331_),
    .X(_05475_));
 sky130_fd_sc_hd__nor2_1 _10780_ (.A(_05278_),
    .B(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__nor2_1 _10781_ (.A(_05244_),
    .B(_05334_),
    .Y(_05477_));
 sky130_fd_sc_hd__or2_2 _10782_ (.A(_05434_),
    .B(_05477_),
    .X(_05478_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(_03510_),
    .A1(_03518_),
    .S(_05229_),
    .X(_05479_));
 sky130_fd_sc_hd__mux4_1 _10784_ (.A0(_05479_),
    .A1(_05441_),
    .A2(_05401_),
    .A3(_05342_),
    .S0(_05266_),
    .S1(_05395_),
    .X(_05480_));
 sky130_fd_sc_hd__mux2_1 _10785_ (.A0(_05249_),
    .A1(_05480_),
    .S(_05288_),
    .X(_05481_));
 sky130_fd_sc_hd__a2bb2o_1 _10786_ (.A1_N(_05476_),
    .A2_N(_05478_),
    .B1(_05399_),
    .B2(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__a211o_1 _10787_ (.A1(_05225_),
    .A2(_05470_),
    .B1(_05474_),
    .C1(_05482_),
    .X(\alu_out[8] ));
 sky130_fd_sc_hd__mux4_1 _10788_ (.A0(net98),
    .A1(_03510_),
    .A2(_03518_),
    .A3(net95),
    .S0(_05236_),
    .S1(_05309_),
    .X(_05483_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(_05483_),
    .A1(_05416_),
    .S(_05295_),
    .X(_05484_));
 sky130_fd_sc_hd__mux2_1 _10790_ (.A0(_05285_),
    .A1(_05484_),
    .S(_05244_),
    .X(_05485_));
 sky130_fd_sc_hd__a2bb2o_1 _10791_ (.A1_N(_03514_),
    .A2_N(_05440_),
    .B1(_05399_),
    .B2(_05485_),
    .X(_05486_));
 sky130_fd_sc_hd__nor2_1 _10792_ (.A(_03530_),
    .B(_05320_),
    .Y(_05487_));
 sky130_fd_sc_hd__o21a_1 _10793_ (.A1(_03530_),
    .A2(_05291_),
    .B1(_05228_),
    .X(_05488_));
 sky130_fd_sc_hd__o21ai_1 _10794_ (.A1(_05287_),
    .A2(_05311_),
    .B1(_05488_),
    .Y(_05489_));
 sky130_fd_sc_hd__o221a_1 _10795_ (.A1(_03513_),
    .A2(_05367_),
    .B1(_05357_),
    .B2(_03515_),
    .C1(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__o21ai_1 _10796_ (.A1(_05478_),
    .A2(_05487_),
    .B1(_05490_),
    .Y(_05491_));
 sky130_fd_sc_hd__o21ai_1 _10797_ (.A1(_03512_),
    .A2(_05468_),
    .B1(_03511_),
    .Y(_05492_));
 sky130_fd_sc_hd__a21oi_1 _10798_ (.A1(_03550_),
    .A2(_04419_),
    .B1(_05322_),
    .Y(_05493_));
 sky130_fd_sc_hd__nand2_1 _10799_ (.A(_03512_),
    .B(_03549_),
    .Y(_05494_));
 sky130_fd_sc_hd__a22o_1 _10800_ (.A1(_05323_),
    .A2(_05492_),
    .B1(_05493_),
    .B2(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__xor2_1 _10801_ (.A(_03515_),
    .B(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__nor2_1 _10802_ (.A(_05218_),
    .B(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__or3_2 _10803_ (.A(_05486_),
    .B(_05491_),
    .C(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__buf_1 _10804_ (.A(_05498_),
    .X(\alu_out[9] ));
 sky130_fd_sc_hd__a31oi_1 _10805_ (.A1(_03512_),
    .A2(_03515_),
    .A3(_03549_),
    .B1(_03552_),
    .Y(_05499_));
 sky130_fd_sc_hd__or4_1 _10806_ (.A(_03512_),
    .B(_03515_),
    .C(_03613_),
    .D(_05467_),
    .X(_05500_));
 sky130_fd_sc_hd__a21o_1 _10807_ (.A1(_03511_),
    .A2(_03514_),
    .B1(_03513_),
    .X(_05501_));
 sky130_fd_sc_hd__and2_1 _10808_ (.A(_05500_),
    .B(_05501_),
    .X(_05502_));
 sky130_fd_sc_hd__inv_2 _10809_ (.A(_05502_),
    .Y(_05503_));
 sky130_fd_sc_hd__mux2_1 _10810_ (.A0(_05499_),
    .A1(_05503_),
    .S(_05363_),
    .X(_05504_));
 sky130_fd_sc_hd__xnor2_1 _10811_ (.A(_03507_),
    .B(_05504_),
    .Y(_05505_));
 sky130_fd_sc_hd__o21a_1 _10812_ (.A1(_05278_),
    .A2(_05349_),
    .B1(_05228_),
    .X(_05506_));
 sky130_fd_sc_hd__o21ai_1 _10813_ (.A1(_05288_),
    .A2(_05332_),
    .B1(_05506_),
    .Y(_05507_));
 sky130_fd_sc_hd__nand2_1 _10814_ (.A(_03507_),
    .B(_05220_),
    .Y(_05508_));
 sky130_fd_sc_hd__o221a_1 _10815_ (.A1(_03506_),
    .A2(_05440_),
    .B1(_05367_),
    .B2(_03505_),
    .C1(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__mux2_1 _10816_ (.A0(net68),
    .A1(net98),
    .S(_05229_),
    .X(_05510_));
 sky130_fd_sc_hd__mux2_1 _10817_ (.A0(_05510_),
    .A1(_05479_),
    .S(_05235_),
    .X(_05511_));
 sky130_fd_sc_hd__mux2_1 _10818_ (.A0(_05511_),
    .A1(_05442_),
    .S(_05295_),
    .X(_05512_));
 sky130_fd_sc_hd__mux2_1 _10819_ (.A0(_05345_),
    .A1(_05512_),
    .S(_05287_),
    .X(_05513_));
 sky130_fd_sc_hd__nor2_1 _10820_ (.A(_05292_),
    .B(_05336_),
    .Y(_05514_));
 sky130_fd_sc_hd__o2bb2a_1 _10821_ (.A1_N(_05399_),
    .A2_N(_05513_),
    .B1(_05514_),
    .B2(_05478_),
    .X(_05515_));
 sky130_fd_sc_hd__and3_1 _10822_ (.A(_05507_),
    .B(_05509_),
    .C(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__o21ai_2 _10823_ (.A1(_05219_),
    .A2(_05505_),
    .B1(_05516_),
    .Y(\alu_out[10] ));
 sky130_fd_sc_hd__buf_4 _10824_ (.A(instr_sub),
    .X(_05517_));
 sky130_fd_sc_hd__o21bai_1 _10825_ (.A1(_03507_),
    .A2(_05499_),
    .B1_N(_03553_),
    .Y(_05518_));
 sky130_fd_sc_hd__o211a_1 _10826_ (.A1(_03505_),
    .A2(_05502_),
    .B1(_03506_),
    .C1(_05390_),
    .X(_05519_));
 sky130_fd_sc_hd__a21o_1 _10827_ (.A1(_05517_),
    .A2(_05518_),
    .B1(_05519_),
    .X(_05520_));
 sky130_fd_sc_hd__xor2_2 _10828_ (.A(_03504_),
    .B(_05520_),
    .X(_05521_));
 sky130_fd_sc_hd__a21oi_1 _10829_ (.A1(_03501_),
    .A2(_05220_),
    .B1(_05301_),
    .Y(_05522_));
 sky130_fd_sc_hd__mux2_1 _10830_ (.A0(_05370_),
    .A1(_05372_),
    .S(_05331_),
    .X(_05523_));
 sky130_fd_sc_hd__o21a_1 _10831_ (.A1(_05278_),
    .A2(_05523_),
    .B1(_05228_),
    .X(_05524_));
 sky130_fd_sc_hd__o21ai_1 _10832_ (.A1(_05288_),
    .A2(_05381_),
    .B1(_05524_),
    .Y(_05525_));
 sky130_fd_sc_hd__o221a_1 _10833_ (.A1(_03501_),
    .A2(_05440_),
    .B1(_05522_),
    .B2(_03503_),
    .C1(_05525_),
    .X(_05526_));
 sky130_fd_sc_hd__mux4_1 _10834_ (.A0(net69),
    .A1(net68),
    .A2(net98),
    .A3(_03510_),
    .S0(_05236_),
    .S1(_05309_),
    .X(_05527_));
 sky130_fd_sc_hd__mux2_1 _10835_ (.A0(_05527_),
    .A1(_05460_),
    .S(_05246_),
    .X(_05528_));
 sky130_fd_sc_hd__mux2_1 _10836_ (.A0(_05377_),
    .A1(_05528_),
    .S(_05287_),
    .X(_05529_));
 sky130_fd_sc_hd__nor2_1 _10837_ (.A(_03530_),
    .B(_05384_),
    .Y(_05530_));
 sky130_fd_sc_hd__o2bb2a_1 _10838_ (.A1_N(_05399_),
    .A2_N(_05529_),
    .B1(_05530_),
    .B2(_05478_),
    .X(_05531_));
 sky130_fd_sc_hd__o211ai_4 _10839_ (.A1(_05219_),
    .A2(_05521_),
    .B1(_05526_),
    .C1(_05531_),
    .Y(\alu_out[11] ));
 sky130_fd_sc_hd__o211a_1 _10840_ (.A1(_03503_),
    .A2(_03506_),
    .B1(_05501_),
    .C1(_03501_),
    .X(_05532_));
 sky130_fd_sc_hd__a21o_1 _10841_ (.A1(_03501_),
    .A2(_03505_),
    .B1(_03503_),
    .X(_05533_));
 sky130_fd_sc_hd__a21o_1 _10842_ (.A1(_05500_),
    .A2(_05532_),
    .B1(_05533_),
    .X(_05534_));
 sky130_fd_sc_hd__mux2_1 _10843_ (.A0(_03556_),
    .A1(_05534_),
    .S(_05390_),
    .X(_05535_));
 sky130_fd_sc_hd__nand2_1 _10844_ (.A(_03499_),
    .B(_05535_),
    .Y(_05536_));
 sky130_fd_sc_hd__or2_1 _10845_ (.A(_03499_),
    .B(_05535_),
    .X(_05537_));
 sky130_fd_sc_hd__mux4_2 _10846_ (.A0(_05234_),
    .A1(_05267_),
    .A2(_05270_),
    .A3(_05273_),
    .S0(_05413_),
    .S1(_05414_),
    .X(_05538_));
 sky130_fd_sc_hd__o21a_1 _10847_ (.A1(_05331_),
    .A2(_05276_),
    .B1(_05423_),
    .X(_05539_));
 sky130_fd_sc_hd__nor2_1 _10848_ (.A(_05292_),
    .B(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__o22a_1 _10849_ (.A1(_03498_),
    .A2(_05398_),
    .B1(_05367_),
    .B2(_03497_),
    .X(_05541_));
 sky130_fd_sc_hd__o221a_1 _10850_ (.A1(_03499_),
    .A2(_05357_),
    .B1(_05478_),
    .B2(_05540_),
    .C1(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__mux2_1 _10851_ (.A0(_04566_),
    .A1(_04532_),
    .S(_05264_),
    .X(_05543_));
 sky130_fd_sc_hd__mux4_2 _10852_ (.A0(_05543_),
    .A1(_05510_),
    .A2(_05479_),
    .A3(_05441_),
    .S0(_05266_),
    .S1(_05243_),
    .X(_05544_));
 sky130_fd_sc_hd__nor2_1 _10853_ (.A(_05292_),
    .B(_05544_),
    .Y(_05545_));
 sky130_fd_sc_hd__a211o_1 _10854_ (.A1(_05414_),
    .A2(_05404_),
    .B1(_05545_),
    .C1(_05250_),
    .X(_05546_));
 sky130_fd_sc_hd__nand2_1 _10855_ (.A(_05542_),
    .B(_05546_),
    .Y(_05547_));
 sky130_fd_sc_hd__a21o_1 _10856_ (.A1(_05298_),
    .A2(_05538_),
    .B1(_05547_),
    .X(_05548_));
 sky130_fd_sc_hd__a31o_2 _10857_ (.A1(_05361_),
    .A2(_05536_),
    .A3(_05537_),
    .B1(_05548_),
    .X(\alu_out[12] ));
 sky130_fd_sc_hd__a21oi_1 _10858_ (.A1(_03499_),
    .A2(_03556_),
    .B1(_03557_),
    .Y(_05549_));
 sky130_fd_sc_hd__and2_1 _10859_ (.A(_03498_),
    .B(_05534_),
    .X(_05550_));
 sky130_fd_sc_hd__nor2_1 _10860_ (.A(_03497_),
    .B(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(_05549_),
    .A1(_05551_),
    .S(_05363_),
    .X(_05552_));
 sky130_fd_sc_hd__xor2_1 _10862_ (.A(_03496_),
    .B(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__nor2_1 _10863_ (.A(_05414_),
    .B(_05424_),
    .Y(_05554_));
 sky130_fd_sc_hd__or2_1 _10864_ (.A(_03494_),
    .B(_05367_),
    .X(_05555_));
 sky130_fd_sc_hd__o221a_1 _10865_ (.A1(_03495_),
    .A2(_05440_),
    .B1(_05357_),
    .B2(_03496_),
    .C1(_05555_),
    .X(_05556_));
 sky130_fd_sc_hd__or2_1 _10866_ (.A(_05226_),
    .B(_05227_),
    .X(_05557_));
 sky130_fd_sc_hd__nor2_1 _10867_ (.A(_05288_),
    .B(_05422_),
    .Y(_05558_));
 sky130_fd_sc_hd__mux2_1 _10868_ (.A0(_05290_),
    .A1(_05306_),
    .S(_05331_),
    .X(_05559_));
 sky130_fd_sc_hd__nor2_1 _10869_ (.A(_05278_),
    .B(_05559_),
    .Y(_05560_));
 sky130_fd_sc_hd__mux4_1 _10870_ (.A0(net71),
    .A1(net70),
    .A2(net69),
    .A3(net68),
    .S0(_05264_),
    .S1(_05235_),
    .X(_05561_));
 sky130_fd_sc_hd__mux2_1 _10871_ (.A0(_05561_),
    .A1(_05483_),
    .S(_05295_),
    .X(_05562_));
 sky130_fd_sc_hd__nand2_1 _10872_ (.A(_05287_),
    .B(_05562_),
    .Y(_05563_));
 sky130_fd_sc_hd__o21a_1 _10873_ (.A1(_05287_),
    .A2(_05418_),
    .B1(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__o32a_1 _10874_ (.A1(_05557_),
    .A2(_05558_),
    .A3(_05560_),
    .B1(_05564_),
    .B2(_05250_),
    .X(_05565_));
 sky130_fd_sc_hd__o211a_1 _10875_ (.A1(_05478_),
    .A2(_05554_),
    .B1(_05556_),
    .C1(_05565_),
    .X(_05566_));
 sky130_fd_sc_hd__o21ai_2 _10876_ (.A1(_05219_),
    .A2(_05553_),
    .B1(_05566_),
    .Y(\alu_out[13] ));
 sky130_fd_sc_hd__o31a_1 _10877_ (.A1(_03494_),
    .A2(_03497_),
    .A3(_05550_),
    .B1(_03495_),
    .X(_05567_));
 sky130_fd_sc_hd__mux2_1 _10878_ (.A0(_03560_),
    .A1(_05567_),
    .S(_05363_),
    .X(_05568_));
 sky130_fd_sc_hd__xor2_1 _10879_ (.A(_03493_),
    .B(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__inv_2 _10880_ (.A(_05444_),
    .Y(_05570_));
 sky130_fd_sc_hd__mux2_1 _10881_ (.A0(net72),
    .A1(_04602_),
    .S(_05264_),
    .X(_05571_));
 sky130_fd_sc_hd__mux2_1 _10882_ (.A0(_05571_),
    .A1(_05543_),
    .S(_05240_),
    .X(_05572_));
 sky130_fd_sc_hd__mux2_1 _10883_ (.A0(_05572_),
    .A1(_05511_),
    .S(_05395_),
    .X(_05573_));
 sky130_fd_sc_hd__mux2_1 _10884_ (.A0(_05570_),
    .A1(_05573_),
    .S(_05288_),
    .X(_05574_));
 sky130_fd_sc_hd__nor2_1 _10885_ (.A(_05278_),
    .B(_05437_),
    .Y(_05575_));
 sky130_fd_sc_hd__o22a_1 _10886_ (.A1(_03492_),
    .A2(_05398_),
    .B1(_05367_),
    .B2(_03491_),
    .X(_05576_));
 sky130_fd_sc_hd__o221a_1 _10887_ (.A1(_03493_),
    .A2(_05357_),
    .B1(_05478_),
    .B2(_05575_),
    .C1(_05576_),
    .X(_05577_));
 sky130_fd_sc_hd__a21bo_1 _10888_ (.A1(_05399_),
    .A2(_05574_),
    .B1_N(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(_05348_),
    .A1(_05329_),
    .S(_05413_),
    .X(_05579_));
 sky130_fd_sc_hd__nand2_1 _10890_ (.A(_05414_),
    .B(_05436_),
    .Y(_05580_));
 sky130_fd_sc_hd__o211a_1 _10891_ (.A1(_05414_),
    .A2(_05579_),
    .B1(_05580_),
    .C1(_05298_),
    .X(_05581_));
 sky130_fd_sc_hd__a211o_1 _10892_ (.A1(_05225_),
    .A2(_05569_),
    .B1(_05578_),
    .C1(_05581_),
    .X(\alu_out[14] ));
 sky130_fd_sc_hd__o21a_1 _10893_ (.A1(_03491_),
    .A2(_05567_),
    .B1(_03492_),
    .X(_05582_));
 sky130_fd_sc_hd__mux2_1 _10894_ (.A0(_03562_),
    .A1(_05582_),
    .S(_05390_),
    .X(_05583_));
 sky130_fd_sc_hd__nand2_1 _10895_ (.A(_03619_),
    .B(_05583_),
    .Y(_05584_));
 sky130_fd_sc_hd__or2_1 _10896_ (.A(_03619_),
    .B(_05583_),
    .X(_05585_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(_05372_),
    .A1(_05379_),
    .S(_05295_),
    .X(_05586_));
 sky130_fd_sc_hd__or2_1 _10898_ (.A(_05292_),
    .B(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__o211a_1 _10899_ (.A1(_05288_),
    .A2(_05455_),
    .B1(_05587_),
    .C1(_05298_),
    .X(_05588_));
 sky130_fd_sc_hd__mux4_1 _10900_ (.A0(_04642_),
    .A1(net72),
    .A2(net71),
    .A3(net70),
    .S0(_05236_),
    .S1(_05309_),
    .X(_05589_));
 sky130_fd_sc_hd__mux2_1 _10901_ (.A0(_05589_),
    .A1(_05527_),
    .S(_05242_),
    .X(_05590_));
 sky130_fd_sc_hd__mux2_1 _10902_ (.A0(_05461_),
    .A1(_05590_),
    .S(_05244_),
    .X(_05591_));
 sky130_fd_sc_hd__and2_1 _10903_ (.A(_05399_),
    .B(_05591_),
    .X(_05592_));
 sky130_fd_sc_hd__o2bb2a_1 _10904_ (.A1_N(_03617_),
    .A2_N(_05301_),
    .B1(_05356_),
    .B2(_03619_),
    .X(_05593_));
 sky130_fd_sc_hd__o221a_1 _10905_ (.A1(_03618_),
    .A2(_05440_),
    .B1(_05456_),
    .B2(_05478_),
    .C1(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__or3b_1 _10906_ (.A(_05588_),
    .B(_05592_),
    .C_N(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__a31o_1 _10907_ (.A1(_05361_),
    .A2(_05584_),
    .A3(_05585_),
    .B1(_05595_),
    .X(\alu_out[15] ));
 sky130_fd_sc_hd__nand2_1 _10908_ (.A(_05557_),
    .B(_05316_),
    .Y(_05596_));
 sky130_fd_sc_hd__clkbuf_4 _10909_ (.A(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__mux2_1 _10910_ (.A0(_04708_),
    .A1(_04642_),
    .S(_05230_),
    .X(_05598_));
 sky130_fd_sc_hd__mux4_2 _10911_ (.A0(_05598_),
    .A1(_05571_),
    .A2(_05543_),
    .A3(_05510_),
    .S0(_05286_),
    .S1(_05413_),
    .X(_05599_));
 sky130_fd_sc_hd__nor2_2 _10912_ (.A(_05244_),
    .B(_05250_),
    .Y(_05600_));
 sky130_fd_sc_hd__clkbuf_4 _10913_ (.A(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__o21ai_2 _10914_ (.A1(instr_sll),
    .A2(instr_slli),
    .B1(_05226_),
    .Y(_05602_));
 sky130_fd_sc_hd__nor2_2 _10915_ (.A(_05292_),
    .B(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__nor2_1 _10916_ (.A(_03484_),
    .B(_05398_),
    .Y(_05604_));
 sky130_fd_sc_hd__a221o_1 _10917_ (.A1(_03483_),
    .A2(_05213_),
    .B1(_05334_),
    .B2(_05226_),
    .C1(_05604_),
    .X(_05605_));
 sky130_fd_sc_hd__a221o_1 _10918_ (.A1(_03485_),
    .A2(_05220_),
    .B1(_05249_),
    .B2(_05603_),
    .C1(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__a221o_1 _10919_ (.A1(_05281_),
    .A2(_05599_),
    .B1(_05601_),
    .B2(_05480_),
    .C1(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__a21boi_2 _10920_ (.A1(_03618_),
    .A2(_05582_),
    .B1_N(_03617_),
    .Y(_05608_));
 sky130_fd_sc_hd__mux2_1 _10921_ (.A0(_03564_),
    .A1(_05608_),
    .S(_05390_),
    .X(_05609_));
 sky130_fd_sc_hd__a21oi_1 _10922_ (.A1(_03485_),
    .A2(_05609_),
    .B1(_05218_),
    .Y(_05610_));
 sky130_fd_sc_hd__o21a_1 _10923_ (.A1(_03485_),
    .A2(_05609_),
    .B1(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__a211o_1 _10924_ (.A1(_05279_),
    .A2(_05597_),
    .B1(_05607_),
    .C1(_05611_),
    .X(\alu_out[16] ));
 sky130_fd_sc_hd__or2_1 _10925_ (.A(_03485_),
    .B(_03564_),
    .X(_05612_));
 sky130_fd_sc_hd__nand2_1 _10926_ (.A(_03483_),
    .B(_05608_),
    .Y(_05613_));
 sky130_fd_sc_hd__a21oi_1 _10927_ (.A1(_03484_),
    .A2(_05613_),
    .B1(_05517_),
    .Y(_05614_));
 sky130_fd_sc_hd__a31o_1 _10928_ (.A1(_05517_),
    .A2(_05612_),
    .A3(_03565_),
    .B1(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__xor2_1 _10929_ (.A(_03488_),
    .B(_05615_),
    .X(_05616_));
 sky130_fd_sc_hd__mux4_1 _10930_ (.A0(_04744_),
    .A1(_04708_),
    .A2(_04642_),
    .A3(_04611_),
    .S0(_05237_),
    .S1(_05240_),
    .X(_05617_));
 sky130_fd_sc_hd__mux2_1 _10931_ (.A0(_05617_),
    .A1(_05561_),
    .S(_05395_),
    .X(_05618_));
 sky130_fd_sc_hd__o21a_1 _10932_ (.A1(_05255_),
    .A2(_05321_),
    .B1(_05597_),
    .X(_05619_));
 sky130_fd_sc_hd__or2_1 _10933_ (.A(net107),
    .B(net75),
    .X(_05620_));
 sky130_fd_sc_hd__o21a_2 _10934_ (.A1(instr_sll),
    .A2(instr_slli),
    .B1(_05226_),
    .X(_05621_));
 sky130_fd_sc_hd__nand2_1 _10935_ (.A(_05244_),
    .B(_05621_),
    .Y(_05622_));
 sky130_fd_sc_hd__nor2_1 _10936_ (.A(_05284_),
    .B(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__a221o_1 _10937_ (.A1(_03487_),
    .A2(_05222_),
    .B1(_05215_),
    .B2(_03488_),
    .C1(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__a221o_1 _10938_ (.A1(_05620_),
    .A2(_05301_),
    .B1(_05484_),
    .B2(_05601_),
    .C1(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__a211o_1 _10939_ (.A1(_05281_),
    .A2(_05618_),
    .B1(_05619_),
    .C1(_05625_),
    .X(_05626_));
 sky130_fd_sc_hd__a21o_1 _10940_ (.A1(_05361_),
    .A2(_05616_),
    .B1(_05626_),
    .X(\alu_out[17] ));
 sky130_fd_sc_hd__o21a_1 _10941_ (.A1(_03488_),
    .A2(_05612_),
    .B1(_03568_),
    .X(_05627_));
 sky130_fd_sc_hd__a31o_1 _10942_ (.A1(net106),
    .A2(net74),
    .A3(_05620_),
    .B1(_03487_),
    .X(_05628_));
 sky130_fd_sc_hd__a31o_1 _10943_ (.A1(_03485_),
    .A2(_03488_),
    .A3(_05608_),
    .B1(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__mux2_1 _10944_ (.A0(_05627_),
    .A1(_05629_),
    .S(_05390_),
    .X(_05630_));
 sky130_fd_sc_hd__or2_1 _10945_ (.A(_03482_),
    .B(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__nand2_1 _10946_ (.A(_03482_),
    .B(_05630_),
    .Y(_05632_));
 sky130_fd_sc_hd__mux2_1 _10947_ (.A0(_04754_),
    .A1(_04744_),
    .S(_05230_),
    .X(_05633_));
 sky130_fd_sc_hd__mux2_1 _10948_ (.A0(_05633_),
    .A1(_05598_),
    .S(_05240_),
    .X(_05634_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(_05634_),
    .A1(_05572_),
    .S(_05331_),
    .X(_05635_));
 sky130_fd_sc_hd__a2bb2o_1 _10950_ (.A1_N(_03481_),
    .A2_N(_05397_),
    .B1(_05213_),
    .B2(_03480_),
    .X(_05636_));
 sky130_fd_sc_hd__a221o_1 _10951_ (.A1(_03482_),
    .A2(_05215_),
    .B1(_05334_),
    .B2(_05254_),
    .C1(_05636_),
    .X(_05637_));
 sky130_fd_sc_hd__a221o_1 _10952_ (.A1(_05512_),
    .A2(_05600_),
    .B1(_05603_),
    .B2(_05345_),
    .C1(_05637_),
    .X(_05638_));
 sky130_fd_sc_hd__a221o_1 _10953_ (.A1(_05337_),
    .A2(_05597_),
    .B1(_05635_),
    .B2(_05281_),
    .C1(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__a31o_1 _10954_ (.A1(_05361_),
    .A2(_05631_),
    .A3(_05632_),
    .B1(_05639_),
    .X(\alu_out[18] ));
 sky130_fd_sc_hd__a21boi_1 _10955_ (.A1(_03480_),
    .A2(_05629_),
    .B1_N(_03481_),
    .Y(_05640_));
 sky130_fd_sc_hd__o21ai_1 _10956_ (.A1(_03482_),
    .A2(_05627_),
    .B1(_03569_),
    .Y(_05641_));
 sky130_fd_sc_hd__mux2_1 _10957_ (.A0(_05640_),
    .A1(_05641_),
    .S(_05517_),
    .X(_05642_));
 sky130_fd_sc_hd__xnor2_1 _10958_ (.A(_03479_),
    .B(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__mux4_1 _10959_ (.A0(_04810_),
    .A1(_04754_),
    .A2(_04744_),
    .A3(_04708_),
    .S0(_05237_),
    .S1(_05240_),
    .X(_05644_));
 sky130_fd_sc_hd__mux2_1 _10960_ (.A0(_05644_),
    .A1(_05589_),
    .S(_05331_),
    .X(_05645_));
 sky130_fd_sc_hd__nand2_2 _10961_ (.A(_05226_),
    .B(_05334_),
    .Y(_05646_));
 sky130_fd_sc_hd__o221a_1 _10962_ (.A1(_03477_),
    .A2(_05398_),
    .B1(_05221_),
    .B2(_03476_),
    .C1(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__o21ai_1 _10963_ (.A1(_03478_),
    .A2(_05357_),
    .B1(_05647_),
    .Y(_05648_));
 sky130_fd_sc_hd__a221o_1 _10964_ (.A1(_05377_),
    .A2(_05603_),
    .B1(_05645_),
    .B2(_05251_),
    .C1(_05648_),
    .X(_05649_));
 sky130_fd_sc_hd__a221o_1 _10965_ (.A1(_05385_),
    .A2(_05597_),
    .B1(_05601_),
    .B2(_05528_),
    .C1(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__a21o_1 _10966_ (.A1(_05361_),
    .A2(_05643_),
    .B1(_05650_),
    .X(\alu_out[19] ));
 sky130_fd_sc_hd__a21o_1 _10967_ (.A1(_03477_),
    .A2(_05640_),
    .B1(_03476_),
    .X(_05651_));
 sky130_fd_sc_hd__inv_2 _10968_ (.A(_05651_),
    .Y(_05652_));
 sky130_fd_sc_hd__mux2_1 _10969_ (.A0(_03572_),
    .A1(_05652_),
    .S(_05363_),
    .X(_05653_));
 sky130_fd_sc_hd__xor2_1 _10970_ (.A(_03466_),
    .B(_05653_),
    .X(_05654_));
 sky130_fd_sc_hd__o21a_1 _10971_ (.A1(_05255_),
    .A2(_05394_),
    .B1(_05597_),
    .X(_05655_));
 sky130_fd_sc_hd__o2bb2a_1 _10972_ (.A1_N(_05220_),
    .A2_N(_03466_),
    .B1(_03465_),
    .B2(_05440_),
    .X(_05656_));
 sky130_fd_sc_hd__o21ai_1 _10973_ (.A1(_03464_),
    .A2(_05367_),
    .B1(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__mux2_1 _10974_ (.A0(_04848_),
    .A1(_04810_),
    .S(_05236_),
    .X(_05658_));
 sky130_fd_sc_hd__mux4_1 _10975_ (.A0(_05658_),
    .A1(_05633_),
    .A2(_05598_),
    .A3(_05571_),
    .S0(_05266_),
    .S1(_05395_),
    .X(_05659_));
 sky130_fd_sc_hd__a2bb2o_1 _10976_ (.A1_N(_05404_),
    .A2_N(_05622_),
    .B1(_05659_),
    .B2(_05251_),
    .X(_05660_));
 sky130_fd_sc_hd__a211o_1 _10977_ (.A1(_05544_),
    .A2(_05601_),
    .B1(_05657_),
    .C1(_05660_),
    .X(_05661_));
 sky130_fd_sc_hd__a211o_1 _10978_ (.A1(_05225_),
    .A2(_05654_),
    .B1(_05655_),
    .C1(_05661_),
    .X(\alu_out[20] ));
 sky130_fd_sc_hd__and2_1 _10979_ (.A(_03465_),
    .B(_05651_),
    .X(_05662_));
 sky130_fd_sc_hd__nor2_1 _10980_ (.A(_03466_),
    .B(_03572_),
    .Y(_05663_));
 sky130_fd_sc_hd__a211o_1 _10981_ (.A1(_03573_),
    .A2(_04848_),
    .B1(_05663_),
    .C1(_05323_),
    .X(_05664_));
 sky130_fd_sc_hd__o31a_1 _10982_ (.A1(_05517_),
    .A2(_03464_),
    .A3(_05662_),
    .B1(_05664_),
    .X(_05665_));
 sky130_fd_sc_hd__xnor2_1 _10983_ (.A(_03574_),
    .B(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__mux4_1 _10984_ (.A0(_04880_),
    .A1(_04848_),
    .A2(_04810_),
    .A3(_04754_),
    .S0(_05264_),
    .S1(_05235_),
    .X(_05667_));
 sky130_fd_sc_hd__mux2_1 _10985_ (.A0(_05667_),
    .A1(_05617_),
    .S(_05243_),
    .X(_05668_));
 sky130_fd_sc_hd__o21ai_1 _10986_ (.A1(_03462_),
    .A2(_05398_),
    .B1(_05646_),
    .Y(_05669_));
 sky130_fd_sc_hd__a221o_1 _10987_ (.A1(_03461_),
    .A2(_05301_),
    .B1(_05220_),
    .B2(_03463_),
    .C1(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__a2bb2o_1 _10988_ (.A1_N(_05418_),
    .A2_N(_05622_),
    .B1(_05600_),
    .B2(_05562_),
    .X(_05671_));
 sky130_fd_sc_hd__a211o_1 _10989_ (.A1(_05281_),
    .A2(_05668_),
    .B1(_05670_),
    .C1(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__a21oi_1 _10990_ (.A1(_05425_),
    .A2(_05597_),
    .B1(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__o21ai_1 _10991_ (.A1(_05219_),
    .A2(_05666_),
    .B1(_05673_),
    .Y(\alu_out[21] ));
 sky130_fd_sc_hd__or2b_1 _10992_ (.A(_05255_),
    .B_N(_05439_),
    .X(_05674_));
 sky130_fd_sc_hd__a21oi_1 _10993_ (.A1(_03574_),
    .A2(_05663_),
    .B1(_03577_),
    .Y(_05675_));
 sky130_fd_sc_hd__nor2_1 _10994_ (.A(net112),
    .B(_04880_),
    .Y(_05676_));
 sky130_fd_sc_hd__o31ai_2 _10995_ (.A1(_05676_),
    .A2(_03464_),
    .A3(_05662_),
    .B1(_03462_),
    .Y(_05677_));
 sky130_fd_sc_hd__mux2_1 _10996_ (.A0(_05675_),
    .A1(_05677_),
    .S(_05323_),
    .X(_05678_));
 sky130_fd_sc_hd__nand2_1 _10997_ (.A(_03472_),
    .B(_05678_),
    .Y(_05679_));
 sky130_fd_sc_hd__or2_1 _10998_ (.A(_03472_),
    .B(_05678_),
    .X(_05680_));
 sky130_fd_sc_hd__a21oi_1 _10999_ (.A1(_05679_),
    .A2(_05680_),
    .B1(_05218_),
    .Y(_05681_));
 sky130_fd_sc_hd__mux2_1 _11000_ (.A0(net81),
    .A1(_04880_),
    .S(_05236_),
    .X(_05682_));
 sky130_fd_sc_hd__mux2_1 _11001_ (.A0(_05682_),
    .A1(_05658_),
    .S(_05232_),
    .X(_05683_));
 sky130_fd_sc_hd__mux2_1 _11002_ (.A0(_05683_),
    .A1(_05634_),
    .S(_05395_),
    .X(_05684_));
 sky130_fd_sc_hd__nor2_1 _11003_ (.A(_03471_),
    .B(_05398_),
    .Y(_05685_));
 sky130_fd_sc_hd__a221o_1 _11004_ (.A1(_03470_),
    .A2(_05301_),
    .B1(_05215_),
    .B2(_03473_),
    .C1(_05685_),
    .X(_05686_));
 sky130_fd_sc_hd__a221o_1 _11005_ (.A1(_05573_),
    .A2(_05601_),
    .B1(_05603_),
    .B2(_05570_),
    .C1(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__a21o_1 _11006_ (.A1(_05281_),
    .A2(_05684_),
    .B1(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__a211o_1 _11007_ (.A1(_05597_),
    .A2(_05674_),
    .B1(_05681_),
    .C1(_05688_),
    .X(\alu_out[22] ));
 sky130_fd_sc_hd__mux4_1 _11008_ (.A0(_04945_),
    .A1(_04913_),
    .A2(_04880_),
    .A3(_04848_),
    .S0(_05264_),
    .S1(_05232_),
    .X(_05689_));
 sky130_fd_sc_hd__mux2_1 _11009_ (.A0(_05689_),
    .A1(_05644_),
    .S(_05277_),
    .X(_05690_));
 sky130_fd_sc_hd__a22o_1 _11010_ (.A1(_03467_),
    .A2(_05213_),
    .B1(_05215_),
    .B2(_03469_),
    .X(_05691_));
 sky130_fd_sc_hd__o21ai_1 _11011_ (.A1(_03468_),
    .A2(_05440_),
    .B1(_05646_),
    .Y(_05692_));
 sky130_fd_sc_hd__a211o_1 _11012_ (.A1(_05461_),
    .A2(_05603_),
    .B1(_05691_),
    .C1(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__a221o_1 _11013_ (.A1(_05590_),
    .A2(_05601_),
    .B1(_05690_),
    .B2(_05281_),
    .C1(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__o21ba_1 _11014_ (.A1(instr_sub),
    .A2(_04913_),
    .B1_N(_03578_),
    .X(_05695_));
 sky130_fd_sc_hd__a31o_1 _11015_ (.A1(_05323_),
    .A2(_03470_),
    .A3(_05677_),
    .B1(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__o31ai_1 _11016_ (.A1(_05363_),
    .A2(_03473_),
    .A3(_05675_),
    .B1(_05696_),
    .Y(_05697_));
 sky130_fd_sc_hd__xor2_1 _11017_ (.A(_03469_),
    .B(_05697_),
    .X(_05698_));
 sky130_fd_sc_hd__nor2_1 _11018_ (.A(_05219_),
    .B(_05698_),
    .Y(_05699_));
 sky130_fd_sc_hd__a211o_1 _11019_ (.A1(_05458_),
    .A2(_05597_),
    .B1(_05694_),
    .C1(_05699_),
    .X(\alu_out[23] ));
 sky130_fd_sc_hd__a21oi_4 _11020_ (.A1(_05244_),
    .A2(_05228_),
    .B1(_05334_),
    .Y(_05700_));
 sky130_fd_sc_hd__nor2_1 _11021_ (.A(_05476_),
    .B(_05700_),
    .Y(_05701_));
 sky130_fd_sc_hd__mux2_1 _11022_ (.A0(_04959_),
    .A1(_04945_),
    .S(_05230_),
    .X(_05702_));
 sky130_fd_sc_hd__mux4_1 _11023_ (.A0(_05702_),
    .A1(_05682_),
    .A2(_05658_),
    .A3(_05633_),
    .S0(_05266_),
    .S1(_05395_),
    .X(_05703_));
 sky130_fd_sc_hd__and3_1 _11024_ (.A(_05288_),
    .B(_05399_),
    .C(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__a2bb2o_1 _11025_ (.A1_N(_03457_),
    .A2_N(_05221_),
    .B1(_05215_),
    .B2(_03459_),
    .X(_05705_));
 sky130_fd_sc_hd__a221o_1 _11026_ (.A1(_03458_),
    .A2(_05222_),
    .B1(_05597_),
    .B2(_05254_),
    .C1(_05705_),
    .X(_05706_));
 sky130_fd_sc_hd__a2111o_1 _11027_ (.A1(_05599_),
    .A2(_05601_),
    .B1(_05701_),
    .C1(_05704_),
    .D1(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__a21boi_1 _11028_ (.A1(_03468_),
    .A2(_03471_),
    .B1_N(_03467_),
    .Y(_05708_));
 sky130_fd_sc_hd__a31o_1 _11029_ (.A1(_03469_),
    .A2(_03473_),
    .A3(_05677_),
    .B1(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__mux2_1 _11030_ (.A0(_03581_),
    .A1(_05709_),
    .S(_05390_),
    .X(_05710_));
 sky130_fd_sc_hd__xnor2_1 _11031_ (.A(_03459_),
    .B(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__nor2_1 _11032_ (.A(_05219_),
    .B(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__a211o_1 _11033_ (.A1(_05481_),
    .A2(_05621_),
    .B1(_05707_),
    .C1(_05712_),
    .X(\alu_out[24] ));
 sky130_fd_sc_hd__mux4_1 _11034_ (.A0(_05013_),
    .A1(_04959_),
    .A2(_04945_),
    .A3(net81),
    .S0(_05264_),
    .S1(_05232_),
    .X(_05713_));
 sky130_fd_sc_hd__mux2_1 _11035_ (.A0(_05713_),
    .A1(_05667_),
    .S(_05246_),
    .X(_05714_));
 sky130_fd_sc_hd__and3_1 _11036_ (.A(_05287_),
    .B(_05399_),
    .C(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__a221o_1 _11037_ (.A1(_03456_),
    .A2(_05220_),
    .B1(_05600_),
    .B2(_05618_),
    .C1(_05715_),
    .X(_05716_));
 sky130_fd_sc_hd__o21bai_2 _11038_ (.A1(_05477_),
    .A2(_05487_),
    .B1_N(_05254_),
    .Y(_05717_));
 sky130_fd_sc_hd__a2bb2o_1 _11039_ (.A1_N(_03455_),
    .A2_N(_05367_),
    .B1(_05222_),
    .B2(_03454_),
    .X(_05718_));
 sky130_fd_sc_hd__a221o_1 _11040_ (.A1(_05485_),
    .A2(_05621_),
    .B1(_05717_),
    .B2(_05597_),
    .C1(_05718_),
    .X(_05719_));
 sky130_fd_sc_hd__nor2_1 _11041_ (.A(_03458_),
    .B(_05709_),
    .Y(_05720_));
 sky130_fd_sc_hd__nand2_1 _11042_ (.A(instr_sub),
    .B(_03582_),
    .Y(_05721_));
 sky130_fd_sc_hd__o32a_1 _11043_ (.A1(instr_sub),
    .A2(_03457_),
    .A3(_05720_),
    .B1(_05721_),
    .B2(_03585_),
    .X(_05722_));
 sky130_fd_sc_hd__nand2_1 _11044_ (.A(_03456_),
    .B(_05722_),
    .Y(_05723_));
 sky130_fd_sc_hd__or2_1 _11045_ (.A(_03456_),
    .B(_05722_),
    .X(_05724_));
 sky130_fd_sc_hd__a21oi_1 _11046_ (.A1(_05723_),
    .A2(_05724_),
    .B1(_05218_),
    .Y(_05725_));
 sky130_fd_sc_hd__or3_1 _11047_ (.A(_05716_),
    .B(_05719_),
    .C(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__clkbuf_1 _11048_ (.A(_05726_),
    .X(\alu_out[25] ));
 sky130_fd_sc_hd__and2_1 _11049_ (.A(_05513_),
    .B(_05621_),
    .X(_05727_));
 sky130_fd_sc_hd__nor2_1 _11050_ (.A(_05514_),
    .B(_05700_),
    .Y(_05728_));
 sky130_fd_sc_hd__mux2_1 _11051_ (.A0(_05044_),
    .A1(_05013_),
    .S(_05230_),
    .X(_05729_));
 sky130_fd_sc_hd__mux2_1 _11052_ (.A0(_05729_),
    .A1(_05702_),
    .S(_05266_),
    .X(_05730_));
 sky130_fd_sc_hd__or2b_1 _11053_ (.A(_05683_),
    .B_N(_05243_),
    .X(_05731_));
 sky130_fd_sc_hd__o211a_1 _11054_ (.A1(_05277_),
    .A2(_05730_),
    .B1(_05731_),
    .C1(_05251_),
    .X(_05732_));
 sky130_fd_sc_hd__o221a_1 _11055_ (.A1(_03451_),
    .A2(_05397_),
    .B1(_05221_),
    .B2(_03450_),
    .C1(_05646_),
    .X(_05733_));
 sky130_fd_sc_hd__o21ai_1 _11056_ (.A1(_03452_),
    .A2(_05357_),
    .B1(_05733_),
    .Y(_05734_));
 sky130_fd_sc_hd__a2111o_1 _11057_ (.A1(_05600_),
    .A2(_05635_),
    .B1(_05728_),
    .C1(_05732_),
    .D1(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__o21ai_1 _11058_ (.A1(_03456_),
    .A2(_03582_),
    .B1(_03587_),
    .Y(_05736_));
 sky130_fd_sc_hd__or2_1 _11059_ (.A(_03455_),
    .B(_03457_),
    .X(_05737_));
 sky130_fd_sc_hd__o21ba_1 _11060_ (.A1(_05720_),
    .A2(_05737_),
    .B1_N(_03454_),
    .X(_05738_));
 sky130_fd_sc_hd__mux2_1 _11061_ (.A0(_05736_),
    .A1(_05738_),
    .S(_05322_),
    .X(_05739_));
 sky130_fd_sc_hd__nand2_1 _11062_ (.A(_03452_),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__or2_1 _11063_ (.A(_03452_),
    .B(_05739_),
    .X(_05741_));
 sky130_fd_sc_hd__and3_1 _11064_ (.A(_05225_),
    .B(_05740_),
    .C(_05741_),
    .X(_05742_));
 sky130_fd_sc_hd__or3_1 _11065_ (.A(_05727_),
    .B(_05735_),
    .C(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__clkbuf_1 _11066_ (.A(_05743_),
    .X(\alu_out[26] ));
 sky130_fd_sc_hd__and2_1 _11067_ (.A(_05529_),
    .B(_05621_),
    .X(_05744_));
 sky130_fd_sc_hd__nor2_1 _11068_ (.A(_05530_),
    .B(_05700_),
    .Y(_05745_));
 sky130_fd_sc_hd__mux4_1 _11069_ (.A0(_05076_),
    .A1(_05044_),
    .A2(_05013_),
    .A3(_04959_),
    .S0(_05237_),
    .S1(_05266_),
    .X(_05746_));
 sky130_fd_sc_hd__or2b_1 _11070_ (.A(_05689_),
    .B_N(_05243_),
    .X(_05747_));
 sky130_fd_sc_hd__o211a_1 _11071_ (.A1(_05277_),
    .A2(_05746_),
    .B1(_05747_),
    .C1(_05251_),
    .X(_05748_));
 sky130_fd_sc_hd__o221a_1 _11072_ (.A1(_03448_),
    .A2(_05397_),
    .B1(_05221_),
    .B2(_03447_),
    .C1(_05646_),
    .X(_05749_));
 sky130_fd_sc_hd__o21ai_1 _11073_ (.A1(_03449_),
    .A2(_05357_),
    .B1(_05749_),
    .Y(_05750_));
 sky130_fd_sc_hd__a2111o_1 _11074_ (.A1(_05600_),
    .A2(_05645_),
    .B1(_05745_),
    .C1(_05748_),
    .D1(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__or2_1 _11075_ (.A(_03450_),
    .B(_05738_),
    .X(_05752_));
 sky130_fd_sc_hd__a21oi_1 _11076_ (.A1(_03452_),
    .A2(_05736_),
    .B1(_03588_),
    .Y(_05753_));
 sky130_fd_sc_hd__nor2_1 _11077_ (.A(_05323_),
    .B(_05753_),
    .Y(_05754_));
 sky130_fd_sc_hd__a31o_1 _11078_ (.A1(_05323_),
    .A2(_03451_),
    .A3(_05752_),
    .B1(_05754_),
    .X(_05755_));
 sky130_fd_sc_hd__xnor2_1 _11079_ (.A(_03449_),
    .B(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__nor2_1 _11080_ (.A(_05218_),
    .B(_05756_),
    .Y(_05757_));
 sky130_fd_sc_hd__or3_1 _11081_ (.A(_05744_),
    .B(_05751_),
    .C(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__clkbuf_1 _11082_ (.A(_05758_),
    .X(\alu_out[27] ));
 sky130_fd_sc_hd__a31o_1 _11083_ (.A1(_03448_),
    .A2(_03451_),
    .A3(_05752_),
    .B1(_03447_),
    .X(_05759_));
 sky130_fd_sc_hd__inv_2 _11084_ (.A(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__mux2_1 _11085_ (.A0(_03591_),
    .A1(_05760_),
    .S(_05363_),
    .X(_05761_));
 sky130_fd_sc_hd__xnor2_1 _11086_ (.A(_03442_),
    .B(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__a211o_1 _11087_ (.A1(_05414_),
    .A2(_05404_),
    .B1(_05545_),
    .C1(_05602_),
    .X(_05763_));
 sky130_fd_sc_hd__mux2_1 _11088_ (.A0(_05086_),
    .A1(_05076_),
    .S(_05237_),
    .X(_05764_));
 sky130_fd_sc_hd__mux4_1 _11089_ (.A0(_05764_),
    .A1(_05729_),
    .A2(_05702_),
    .A3(_05682_),
    .S0(_05266_),
    .S1(_05331_),
    .X(_05765_));
 sky130_fd_sc_hd__o221ai_2 _11090_ (.A1(_03441_),
    .A2(_05398_),
    .B1(_05367_),
    .B2(_03440_),
    .C1(_05646_),
    .Y(_05766_));
 sky130_fd_sc_hd__a221o_1 _11091_ (.A1(_03442_),
    .A2(_05220_),
    .B1(_05251_),
    .B2(_05765_),
    .C1(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__a21oi_1 _11092_ (.A1(_05601_),
    .A2(_05659_),
    .B1(_05767_),
    .Y(_05768_));
 sky130_fd_sc_hd__o211a_1 _11093_ (.A1(_05540_),
    .A2(_05700_),
    .B1(_05763_),
    .C1(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__o21ai_2 _11094_ (.A1(_05219_),
    .A2(_05762_),
    .B1(_05769_),
    .Y(\alu_out[28] ));
 sky130_fd_sc_hd__nor2_1 _11095_ (.A(_03442_),
    .B(_03591_),
    .Y(_05770_));
 sky130_fd_sc_hd__a21o_1 _11096_ (.A1(_03592_),
    .A2(_05086_),
    .B1(_05390_),
    .X(_05771_));
 sky130_fd_sc_hd__a211o_1 _11097_ (.A1(_03441_),
    .A2(_05759_),
    .B1(_05517_),
    .C1(_03440_),
    .X(_05772_));
 sky130_fd_sc_hd__o21a_1 _11098_ (.A1(_05770_),
    .A2(_05771_),
    .B1(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__xnor2_1 _11099_ (.A(_03445_),
    .B(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__or2_1 _11100_ (.A(_05564_),
    .B(_05602_),
    .X(_05775_));
 sky130_fd_sc_hd__mux4_1 _11101_ (.A0(_05143_),
    .A1(_05086_),
    .A2(_05076_),
    .A3(_05044_),
    .S0(_05324_),
    .S1(_05286_),
    .X(_05776_));
 sky130_fd_sc_hd__mux2_1 _11102_ (.A0(_05776_),
    .A1(_05713_),
    .S(_05413_),
    .X(_05777_));
 sky130_fd_sc_hd__a21o_1 _11103_ (.A1(_03444_),
    .A2(_05215_),
    .B1(_05213_),
    .X(_05778_));
 sky130_fd_sc_hd__o21ai_1 _11104_ (.A1(_03444_),
    .A2(_05398_),
    .B1(_05646_),
    .Y(_05779_));
 sky130_fd_sc_hd__a221o_1 _11105_ (.A1(_05600_),
    .A2(_05668_),
    .B1(_05778_),
    .B2(_03443_),
    .C1(_05779_),
    .X(_05780_));
 sky130_fd_sc_hd__a21oi_1 _11106_ (.A1(_05281_),
    .A2(_05777_),
    .B1(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__o211a_1 _11107_ (.A1(_05554_),
    .A2(_05700_),
    .B1(_05775_),
    .C1(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__o21ai_1 _11108_ (.A1(_05219_),
    .A2(_05774_),
    .B1(_05782_),
    .Y(\alu_out[29] ));
 sky130_fd_sc_hd__a21o_1 _11109_ (.A1(_03445_),
    .A2(_05770_),
    .B1(_03594_),
    .X(_05783_));
 sky130_fd_sc_hd__nor2_1 _11110_ (.A(net120),
    .B(_05143_),
    .Y(_05784_));
 sky130_fd_sc_hd__a211o_1 _11111_ (.A1(_03441_),
    .A2(_05759_),
    .B1(_05784_),
    .C1(_03440_),
    .X(_05785_));
 sky130_fd_sc_hd__a21o_1 _11112_ (.A1(_03444_),
    .A2(_05785_),
    .B1(_05517_),
    .X(_05786_));
 sky130_fd_sc_hd__o21ai_1 _11113_ (.A1(_05363_),
    .A2(_05783_),
    .B1(_05786_),
    .Y(_05787_));
 sky130_fd_sc_hd__xnor2_1 _11114_ (.A(_03438_),
    .B(_05787_),
    .Y(_05788_));
 sky130_fd_sc_hd__nor2_1 _11115_ (.A(_05575_),
    .B(_05700_),
    .Y(_05789_));
 sky130_fd_sc_hd__mux2_1 _11116_ (.A0(_05174_),
    .A1(_05143_),
    .S(_05324_),
    .X(_05790_));
 sky130_fd_sc_hd__mux4_1 _11117_ (.A0(_05790_),
    .A1(_05764_),
    .A2(_05729_),
    .A3(_05702_),
    .S0(_05286_),
    .S1(_05277_),
    .X(_05791_));
 sky130_fd_sc_hd__o22ai_1 _11118_ (.A1(_03435_),
    .A2(_05221_),
    .B1(_05356_),
    .B2(_03438_),
    .Y(_05792_));
 sky130_fd_sc_hd__a221o_1 _11119_ (.A1(_03436_),
    .A2(_05222_),
    .B1(_05596_),
    .B2(_05254_),
    .C1(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__a221o_1 _11120_ (.A1(_05601_),
    .A2(_05684_),
    .B1(_05791_),
    .B2(_05281_),
    .C1(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__a211o_1 _11121_ (.A1(_05574_),
    .A2(_05621_),
    .B1(_05789_),
    .C1(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__a21o_1 _11122_ (.A1(_05361_),
    .A2(_05788_),
    .B1(_05795_),
    .X(\alu_out[30] ));
 sky130_fd_sc_hd__a21oi_1 _11123_ (.A1(_03444_),
    .A2(_05785_),
    .B1(_03435_),
    .Y(_05796_));
 sky130_fd_sc_hd__a21o_1 _11124_ (.A1(_03438_),
    .A2(_05783_),
    .B1(_03595_),
    .X(_05797_));
 sky130_fd_sc_hd__nand2_1 _11125_ (.A(_05517_),
    .B(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__o31a_1 _11126_ (.A1(_05517_),
    .A2(_03436_),
    .A3(_05796_),
    .B1(_05798_),
    .X(_05799_));
 sky130_fd_sc_hd__xor2_1 _11127_ (.A(_03434_),
    .B(_05799_),
    .X(_05800_));
 sky130_fd_sc_hd__nand2_1 _11128_ (.A(_03432_),
    .B(_05301_),
    .Y(_05801_));
 sky130_fd_sc_hd__o221a_1 _11129_ (.A1(_03433_),
    .A2(_05440_),
    .B1(_05357_),
    .B2(_03434_),
    .C1(_05801_),
    .X(_05802_));
 sky130_fd_sc_hd__mux4_1 _11130_ (.A0(_05205_),
    .A1(_05174_),
    .A2(_05143_),
    .A3(_05086_),
    .S0(_05324_),
    .S1(_05286_),
    .X(_05803_));
 sky130_fd_sc_hd__or2b_1 _11131_ (.A(_05746_),
    .B_N(_05395_),
    .X(_05804_));
 sky130_fd_sc_hd__o211a_1 _11132_ (.A1(_05413_),
    .A2(_05803_),
    .B1(_05804_),
    .C1(_05251_),
    .X(_05805_));
 sky130_fd_sc_hd__a221oi_2 _11133_ (.A1(_05591_),
    .A2(_05621_),
    .B1(_05690_),
    .B2(_05601_),
    .C1(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__o211a_1 _11134_ (.A1(_05456_),
    .A2(_05700_),
    .B1(_05802_),
    .C1(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__o21ai_2 _11135_ (.A1(_05219_),
    .A2(_05800_),
    .B1(_05807_),
    .Y(\alu_out[31] ));
 sky130_fd_sc_hd__a2bb2o_2 _11136_ (.A1_N(_04040_),
    .A2_N(_04033_),
    .B1(_04030_),
    .B2(_04422_),
    .X(net259));
 sky130_fd_sc_hd__inv_2 _11137_ (.A(_04030_),
    .Y(_05808_));
 sky130_fd_sc_hd__a211o_2 _11138_ (.A1(_04040_),
    .A2(_04033_),
    .B1(_05808_),
    .C1(_04811_),
    .X(net260));
 sky130_fd_sc_hd__a211o_2 _11139_ (.A1(_04040_),
    .A2(_04037_),
    .B1(_05808_),
    .C1(_04811_),
    .X(net261));
 sky130_fd_sc_hd__a22o_2 _11140_ (.A1(_03407_),
    .A2(_05324_),
    .B1(net129),
    .B2(_04422_),
    .X(net255));
 sky130_fd_sc_hd__a22o_2 _11141_ (.A1(_03407_),
    .A2(_05286_),
    .B1(net130),
    .B2(_04422_),
    .X(net256));
 sky130_fd_sc_hd__a22o_2 _11142_ (.A1(_03407_),
    .A2(_05413_),
    .B1(net100),
    .B2(_04422_),
    .X(net226));
 sky130_fd_sc_hd__a22o_2 _11143_ (.A1(_03407_),
    .A2(_05414_),
    .B1(net101),
    .B2(_04422_),
    .X(net227));
 sky130_fd_sc_hd__a22o_2 _11144_ (.A1(_03407_),
    .A2(_05254_),
    .B1(net102),
    .B2(_04422_),
    .X(net228));
 sky130_fd_sc_hd__a22o_2 _11145_ (.A1(_03407_),
    .A2(net126),
    .B1(net103),
    .B2(_04422_),
    .X(net229));
 sky130_fd_sc_hd__a22o_2 _11146_ (.A1(_03407_),
    .A2(net127),
    .B1(net104),
    .B2(_04422_),
    .X(net230));
 sky130_fd_sc_hd__a22o_2 _11147_ (.A1(_03407_),
    .A2(net128),
    .B1(net105),
    .B2(_04422_),
    .X(net231));
 sky130_fd_sc_hd__mux2_1 _11148_ (.A0(_05324_),
    .A1(net106),
    .S(_04745_),
    .X(_05809_));
 sky130_fd_sc_hd__buf_2 _11149_ (.A(_05809_),
    .X(net232));
 sky130_fd_sc_hd__mux2_1 _11150_ (.A0(_05286_),
    .A1(net107),
    .S(_04745_),
    .X(_05810_));
 sky130_fd_sc_hd__buf_2 _11151_ (.A(_05810_),
    .X(net233));
 sky130_fd_sc_hd__mux2_1 _11152_ (.A0(_05277_),
    .A1(net108),
    .S(_04745_),
    .X(_05811_));
 sky130_fd_sc_hd__buf_2 _11153_ (.A(_05811_),
    .X(net234));
 sky130_fd_sc_hd__mux2_1 _11154_ (.A0(_05292_),
    .A1(net109),
    .S(_04745_),
    .X(_05812_));
 sky130_fd_sc_hd__buf_2 _11155_ (.A(_05812_),
    .X(net235));
 sky130_fd_sc_hd__mux2_1 _11156_ (.A0(_05254_),
    .A1(net111),
    .S(_04668_),
    .X(_05813_));
 sky130_fd_sc_hd__clkbuf_2 _11157_ (.A(_05813_),
    .X(net237));
 sky130_fd_sc_hd__mux2_1 _11158_ (.A0(net126),
    .A1(net112),
    .S(_04668_),
    .X(_05814_));
 sky130_fd_sc_hd__clkbuf_2 _11159_ (.A(_05814_),
    .X(net238));
 sky130_fd_sc_hd__mux2_1 _11160_ (.A0(net127),
    .A1(net113),
    .S(_04668_),
    .X(_05815_));
 sky130_fd_sc_hd__buf_2 _11161_ (.A(_05815_),
    .X(net239));
 sky130_fd_sc_hd__mux2_1 _11162_ (.A0(net128),
    .A1(net114),
    .S(_04668_),
    .X(_05816_));
 sky130_fd_sc_hd__clkbuf_2 _11163_ (.A(_05816_),
    .X(net240));
 sky130_fd_sc_hd__a22o_1 _11164_ (.A1(_03407_),
    .A2(_05324_),
    .B1(net129),
    .B2(_03297_),
    .X(_05817_));
 sky130_fd_sc_hd__a21o_2 _11165_ (.A1(net115),
    .A2(_04710_),
    .B1(_05817_),
    .X(net241));
 sky130_fd_sc_hd__a22o_1 _11166_ (.A1(_04038_),
    .A2(_05286_),
    .B1(net130),
    .B2(_03297_),
    .X(_05818_));
 sky130_fd_sc_hd__a21o_2 _11167_ (.A1(net116),
    .A2(_04710_),
    .B1(_05818_),
    .X(net242));
 sky130_fd_sc_hd__a22o_1 _11168_ (.A1(_04038_),
    .A2(_05277_),
    .B1(net100),
    .B2(_03297_),
    .X(_05819_));
 sky130_fd_sc_hd__a21o_2 _11169_ (.A1(net117),
    .A2(_04710_),
    .B1(_05819_),
    .X(net243));
 sky130_fd_sc_hd__a22o_1 _11170_ (.A1(_04038_),
    .A2(_05292_),
    .B1(net101),
    .B2(_03297_),
    .X(_05820_));
 sky130_fd_sc_hd__a21o_2 _11171_ (.A1(net118),
    .A2(_04710_),
    .B1(_05820_),
    .X(net244));
 sky130_fd_sc_hd__a22o_1 _11172_ (.A1(_04038_),
    .A2(_05254_),
    .B1(net102),
    .B2(_03297_),
    .X(_05821_));
 sky130_fd_sc_hd__a21o_2 _11173_ (.A1(net119),
    .A2(_04710_),
    .B1(_05821_),
    .X(net245));
 sky130_fd_sc_hd__a22o_1 _11174_ (.A1(_04038_),
    .A2(net126),
    .B1(net103),
    .B2(_03297_),
    .X(_05822_));
 sky130_fd_sc_hd__a21o_2 _11175_ (.A1(net120),
    .A2(_04710_),
    .B1(_05822_),
    .X(net246));
 sky130_fd_sc_hd__a22o_1 _11176_ (.A1(_04038_),
    .A2(net127),
    .B1(net104),
    .B2(_03297_),
    .X(_05823_));
 sky130_fd_sc_hd__a21o_2 _11177_ (.A1(net122),
    .A2(_04710_),
    .B1(_05823_),
    .X(net248));
 sky130_fd_sc_hd__a22o_1 _11178_ (.A1(_04038_),
    .A2(net128),
    .B1(net105),
    .B2(_03297_),
    .X(_05824_));
 sky130_fd_sc_hd__a21o_2 _11179_ (.A1(net123),
    .A2(_04710_),
    .B1(_05824_),
    .X(net249));
 sky130_fd_sc_hd__mux2_2 _11180_ (.A0(\reg_next_pc[2] ),
    .A1(\reg_out[2] ),
    .S(_03189_),
    .X(_05825_));
 sky130_fd_sc_hd__xor2_1 _11181_ (.A(_03217_),
    .B(_05825_),
    .X(_05826_));
 sky130_fd_sc_hd__clkbuf_4 _11182_ (.A(_03219_),
    .X(_05827_));
 sky130_fd_sc_hd__mux2_1 _11183_ (.A0(_04160_),
    .A1(_05826_),
    .S(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__buf_4 _11184_ (.A(_05828_),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_8 _11185_ (.A(_03219_),
    .X(_05829_));
 sky130_fd_sc_hd__mux2_1 _11186_ (.A0(\reg_next_pc[3] ),
    .A1(\reg_out[3] ),
    .S(_03189_),
    .X(_05830_));
 sky130_fd_sc_hd__and3_1 _11187_ (.A(_03217_),
    .B(_05825_),
    .C(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__a21oi_1 _11188_ (.A1(_03217_),
    .A2(_05825_),
    .B1(_05830_),
    .Y(_05832_));
 sky130_fd_sc_hd__o21ai_1 _11189_ (.A1(_05831_),
    .A2(_05832_),
    .B1(_05829_),
    .Y(_05833_));
 sky130_fd_sc_hd__o21a_4 _11190_ (.A1(_04198_),
    .A2(_05829_),
    .B1(_05833_),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 _11191_ (.A(_03189_),
    .X(_05834_));
 sky130_fd_sc_hd__mux2_2 _11192_ (.A0(\reg_next_pc[4] ),
    .A1(\reg_out[4] ),
    .S(_05834_),
    .X(_05835_));
 sky130_fd_sc_hd__nand2_1 _11193_ (.A(_05831_),
    .B(_05835_),
    .Y(_05836_));
 sky130_fd_sc_hd__or2_1 _11194_ (.A(_05831_),
    .B(_05835_),
    .X(_05837_));
 sky130_fd_sc_hd__buf_4 _11195_ (.A(_03841_),
    .X(_05838_));
 sky130_fd_sc_hd__and2_1 _11196_ (.A(_04251_),
    .B(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__a31o_4 _11197_ (.A1(_05829_),
    .A2(_05836_),
    .A3(_05837_),
    .B1(_05839_),
    .X(net218));
 sky130_fd_sc_hd__mux2_2 _11198_ (.A0(\reg_next_pc[5] ),
    .A1(\reg_out[5] ),
    .S(_05834_),
    .X(_05840_));
 sky130_fd_sc_hd__xnor2_1 _11199_ (.A(_05836_),
    .B(_05840_),
    .Y(_05841_));
 sky130_fd_sc_hd__mux2_1 _11200_ (.A0(_04262_),
    .A1(_05841_),
    .S(_05827_),
    .X(_05842_));
 sky130_fd_sc_hd__buf_4 _11201_ (.A(_05842_),
    .X(net219));
 sky130_fd_sc_hd__mux2_1 _11202_ (.A0(\reg_next_pc[6] ),
    .A1(\reg_out[6] ),
    .S(_05834_),
    .X(_05843_));
 sky130_fd_sc_hd__and4_1 _11203_ (.A(_05831_),
    .B(_05835_),
    .C(_05840_),
    .D(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__a31o_1 _11204_ (.A1(_05831_),
    .A2(_05835_),
    .A3(_05840_),
    .B1(_05843_),
    .X(_05845_));
 sky130_fd_sc_hd__and2b_1 _11205_ (.A_N(_05844_),
    .B(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__mux2_1 _11206_ (.A0(_04342_),
    .A1(_05846_),
    .S(_05827_),
    .X(_05847_));
 sky130_fd_sc_hd__buf_4 _11207_ (.A(_05847_),
    .X(net220));
 sky130_fd_sc_hd__mux2_2 _11208_ (.A0(\reg_next_pc[7] ),
    .A1(\reg_out[7] ),
    .S(_05834_),
    .X(_05848_));
 sky130_fd_sc_hd__xor2_1 _11209_ (.A(_05844_),
    .B(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__mux2_1 _11210_ (.A0(_04360_),
    .A1(_05849_),
    .S(_05827_),
    .X(_05850_));
 sky130_fd_sc_hd__clkbuf_4 _11211_ (.A(_05850_),
    .X(net221));
 sky130_fd_sc_hd__mux2_1 _11212_ (.A0(\reg_next_pc[8] ),
    .A1(\reg_out[8] ),
    .S(_05834_),
    .X(_05851_));
 sky130_fd_sc_hd__and3_1 _11213_ (.A(_05844_),
    .B(_05848_),
    .C(_05851_),
    .X(_05852_));
 sky130_fd_sc_hd__a21oi_1 _11214_ (.A1(_05844_),
    .A2(_05848_),
    .B1(_05851_),
    .Y(_05853_));
 sky130_fd_sc_hd__nor2_1 _11215_ (.A(_05852_),
    .B(_05853_),
    .Y(_05854_));
 sky130_fd_sc_hd__mux2_1 _11216_ (.A0(_04419_),
    .A1(_05854_),
    .S(_05827_),
    .X(_05855_));
 sky130_fd_sc_hd__clkbuf_4 _11217_ (.A(_05855_),
    .X(net222));
 sky130_fd_sc_hd__buf_2 _11218_ (.A(_03188_),
    .X(_05856_));
 sky130_fd_sc_hd__buf_2 _11219_ (.A(_05856_),
    .X(_05857_));
 sky130_fd_sc_hd__buf_2 _11220_ (.A(_05834_),
    .X(_05858_));
 sky130_fd_sc_hd__or2_1 _11221_ (.A(\reg_next_pc[9] ),
    .B(_05858_),
    .X(_05859_));
 sky130_fd_sc_hd__o21a_1 _11222_ (.A1(\reg_out[9] ),
    .A2(_05857_),
    .B1(_05859_),
    .X(_05860_));
 sky130_fd_sc_hd__nor2_1 _11223_ (.A(_05852_),
    .B(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__and2_2 _11224_ (.A(_05852_),
    .B(_05860_),
    .X(_05862_));
 sky130_fd_sc_hd__nand2_1 _11225_ (.A(_04456_),
    .B(_05838_),
    .Y(_05863_));
 sky130_fd_sc_hd__o31ai_4 _11226_ (.A1(_05838_),
    .A2(_05861_),
    .A3(_05862_),
    .B1(_05863_),
    .Y(net223));
 sky130_fd_sc_hd__mux2_2 _11227_ (.A0(\reg_next_pc[10] ),
    .A1(\reg_out[10] ),
    .S(_05858_),
    .X(_05864_));
 sky130_fd_sc_hd__nand2_1 _11228_ (.A(_05862_),
    .B(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__or2_1 _11229_ (.A(_05862_),
    .B(_05864_),
    .X(_05866_));
 sky130_fd_sc_hd__and2_1 _11230_ (.A(_04466_),
    .B(_03841_),
    .X(_05867_));
 sky130_fd_sc_hd__a31o_4 _11231_ (.A1(_05829_),
    .A2(_05865_),
    .A3(_05866_),
    .B1(_05867_),
    .X(net194));
 sky130_fd_sc_hd__mux2_2 _11232_ (.A0(\reg_next_pc[11] ),
    .A1(\reg_out[11] ),
    .S(_05858_),
    .X(_05868_));
 sky130_fd_sc_hd__xnor2_1 _11233_ (.A(_05865_),
    .B(_05868_),
    .Y(_05869_));
 sky130_fd_sc_hd__mux2_1 _11234_ (.A0(_04532_),
    .A1(_05869_),
    .S(_05827_),
    .X(_05870_));
 sky130_fd_sc_hd__buf_4 _11235_ (.A(_05870_),
    .X(net195));
 sky130_fd_sc_hd__mux2_1 _11236_ (.A0(\reg_next_pc[12] ),
    .A1(\reg_out[12] ),
    .S(_05858_),
    .X(_05871_));
 sky130_fd_sc_hd__and4_1 _11237_ (.A(_05862_),
    .B(_05864_),
    .C(_05868_),
    .D(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__a31o_1 _11238_ (.A1(_05862_),
    .A2(_05864_),
    .A3(_05868_),
    .B1(_05871_),
    .X(_05873_));
 sky130_fd_sc_hd__and2b_1 _11239_ (.A_N(_05872_),
    .B(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__mux2_1 _11240_ (.A0(_04566_),
    .A1(_05874_),
    .S(_05827_),
    .X(_05875_));
 sky130_fd_sc_hd__buf_4 _11241_ (.A(_05875_),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 _11242_ (.A(_05858_),
    .X(_05876_));
 sky130_fd_sc_hd__mux2_2 _11243_ (.A0(\reg_next_pc[13] ),
    .A1(\reg_out[13] ),
    .S(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__nand2_1 _11244_ (.A(_05872_),
    .B(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__or2_1 _11245_ (.A(_05872_),
    .B(_05877_),
    .X(_05879_));
 sky130_fd_sc_hd__and2_1 _11246_ (.A(_04602_),
    .B(_03841_),
    .X(_05880_));
 sky130_fd_sc_hd__a31o_4 _11247_ (.A1(_05829_),
    .A2(_05878_),
    .A3(_05879_),
    .B1(_05880_),
    .X(net197));
 sky130_fd_sc_hd__mux2_2 _11248_ (.A0(\reg_next_pc[14] ),
    .A1(\reg_out[14] ),
    .S(_05876_),
    .X(_05881_));
 sky130_fd_sc_hd__nand2b_1 _11249_ (.A_N(_05878_),
    .B(_05881_),
    .Y(_05882_));
 sky130_fd_sc_hd__a21o_1 _11250_ (.A1(_05872_),
    .A2(_05877_),
    .B1(_05881_),
    .X(_05883_));
 sky130_fd_sc_hd__and2_1 _11251_ (.A(_04611_),
    .B(_03841_),
    .X(_05884_));
 sky130_fd_sc_hd__a31o_4 _11252_ (.A1(_05829_),
    .A2(_05882_),
    .A3(_05883_),
    .B1(_05884_),
    .X(net198));
 sky130_fd_sc_hd__mux2_2 _11253_ (.A0(\reg_next_pc[15] ),
    .A1(\reg_out[15] ),
    .S(_05876_),
    .X(_05885_));
 sky130_fd_sc_hd__xnor2_1 _11254_ (.A(_05882_),
    .B(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__mux2_1 _11255_ (.A0(_04642_),
    .A1(_05886_),
    .S(_05827_),
    .X(_05887_));
 sky130_fd_sc_hd__clkbuf_4 _11256_ (.A(_05887_),
    .X(net199));
 sky130_fd_sc_hd__and2b_1 _11257_ (.A_N(_05882_),
    .B(_05885_),
    .X(_05888_));
 sky130_fd_sc_hd__mux2_1 _11258_ (.A0(\reg_next_pc[16] ),
    .A1(\reg_out[16] ),
    .S(_05876_),
    .X(_05889_));
 sky130_fd_sc_hd__nor2_1 _11259_ (.A(_05888_),
    .B(_05889_),
    .Y(_05890_));
 sky130_fd_sc_hd__and4b_1 _11260_ (.A_N(_05878_),
    .B(_05881_),
    .C(_05885_),
    .D(_05889_),
    .X(_05891_));
 sky130_fd_sc_hd__nand2_1 _11261_ (.A(_04708_),
    .B(_05838_),
    .Y(_05892_));
 sky130_fd_sc_hd__o31ai_4 _11262_ (.A1(_05838_),
    .A2(_05890_),
    .A3(_05891_),
    .B1(_05892_),
    .Y(net200));
 sky130_fd_sc_hd__or2_1 _11263_ (.A(\reg_next_pc[17] ),
    .B(_05876_),
    .X(_05893_));
 sky130_fd_sc_hd__o21a_1 _11264_ (.A1(\reg_out[17] ),
    .A2(_05857_),
    .B1(_05893_),
    .X(_05894_));
 sky130_fd_sc_hd__nor2_1 _11265_ (.A(_05891_),
    .B(_05894_),
    .Y(_05895_));
 sky130_fd_sc_hd__and2_2 _11266_ (.A(_05891_),
    .B(_05894_),
    .X(_05896_));
 sky130_fd_sc_hd__nand2_1 _11267_ (.A(_04744_),
    .B(_05838_),
    .Y(_05897_));
 sky130_fd_sc_hd__o31ai_4 _11268_ (.A1(_05838_),
    .A2(_05895_),
    .A3(_05896_),
    .B1(_05897_),
    .Y(net201));
 sky130_fd_sc_hd__buf_2 _11269_ (.A(_05876_),
    .X(_05898_));
 sky130_fd_sc_hd__mux2_2 _11270_ (.A0(\reg_next_pc[18] ),
    .A1(\reg_out[18] ),
    .S(_05898_),
    .X(_05899_));
 sky130_fd_sc_hd__xor2_1 _11271_ (.A(_05896_),
    .B(_05899_),
    .X(_05900_));
 sky130_fd_sc_hd__mux2_1 _11272_ (.A0(_04754_),
    .A1(_05900_),
    .S(_05827_),
    .X(_05901_));
 sky130_fd_sc_hd__clkbuf_4 _11273_ (.A(_05901_),
    .X(net202));
 sky130_fd_sc_hd__mux2_2 _11274_ (.A0(\reg_next_pc[19] ),
    .A1(\reg_out[19] ),
    .S(_05898_),
    .X(_05902_));
 sky130_fd_sc_hd__a21oi_1 _11275_ (.A1(_05896_),
    .A2(_05899_),
    .B1(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__and3_1 _11276_ (.A(_05896_),
    .B(_05899_),
    .C(_05902_),
    .X(_05904_));
 sky130_fd_sc_hd__or3_1 _11277_ (.A(_03841_),
    .B(_05903_),
    .C(_05904_),
    .X(_05905_));
 sky130_fd_sc_hd__o21ai_4 _11278_ (.A1(_03475_),
    .A2(_05829_),
    .B1(_05905_),
    .Y(net203));
 sky130_fd_sc_hd__mux2_2 _11279_ (.A0(\reg_next_pc[20] ),
    .A1(\reg_out[20] ),
    .S(_05898_),
    .X(_05906_));
 sky130_fd_sc_hd__xor2_1 _11280_ (.A(_05904_),
    .B(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__mux2_1 _11281_ (.A0(_04848_),
    .A1(_05907_),
    .S(_05827_),
    .X(_05908_));
 sky130_fd_sc_hd__clkbuf_4 _11282_ (.A(_05908_),
    .X(net204));
 sky130_fd_sc_hd__buf_2 _11283_ (.A(_05857_),
    .X(_05909_));
 sky130_fd_sc_hd__or2_1 _11284_ (.A(\reg_next_pc[21] ),
    .B(_05898_),
    .X(_05910_));
 sky130_fd_sc_hd__o21a_1 _11285_ (.A1(\reg_out[21] ),
    .A2(_05909_),
    .B1(_05910_),
    .X(_05911_));
 sky130_fd_sc_hd__a21oi_1 _11286_ (.A1(_05904_),
    .A2(_05906_),
    .B1(_05911_),
    .Y(_05912_));
 sky130_fd_sc_hd__and3_1 _11287_ (.A(_05904_),
    .B(_05906_),
    .C(_05911_),
    .X(_05913_));
 sky130_fd_sc_hd__or3_1 _11288_ (.A(_03841_),
    .B(_05912_),
    .C(_05913_),
    .X(_05914_));
 sky130_fd_sc_hd__o21ai_4 _11289_ (.A1(_03575_),
    .A2(_05829_),
    .B1(_05914_),
    .Y(net205));
 sky130_fd_sc_hd__mux2_2 _11290_ (.A0(\reg_next_pc[22] ),
    .A1(\reg_out[22] ),
    .S(_05898_),
    .X(_05915_));
 sky130_fd_sc_hd__xor2_1 _11291_ (.A(_05913_),
    .B(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__mux2_1 _11292_ (.A0(_04913_),
    .A1(_05916_),
    .S(_03219_),
    .X(_05917_));
 sky130_fd_sc_hd__buf_2 _11293_ (.A(_05917_),
    .X(net206));
 sky130_fd_sc_hd__mux2_2 _11294_ (.A0(\reg_next_pc[23] ),
    .A1(\reg_out[23] ),
    .S(_05898_),
    .X(_05918_));
 sky130_fd_sc_hd__a21oi_1 _11295_ (.A1(_05913_),
    .A2(_05915_),
    .B1(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__and3_1 _11296_ (.A(_05913_),
    .B(_05915_),
    .C(_05918_),
    .X(_05920_));
 sky130_fd_sc_hd__or3_1 _11297_ (.A(_03841_),
    .B(_05919_),
    .C(_05920_),
    .X(_05921_));
 sky130_fd_sc_hd__o21ai_4 _11298_ (.A1(_03460_),
    .A2(_05829_),
    .B1(_05921_),
    .Y(net207));
 sky130_fd_sc_hd__or2_2 _11299_ (.A(\reg_next_pc[24] ),
    .B(_05898_),
    .X(_05922_));
 sky130_fd_sc_hd__o21a_1 _11300_ (.A1(\reg_out[24] ),
    .A2(_05909_),
    .B1(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__nor2_1 _11301_ (.A(_05920_),
    .B(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__and2_1 _11302_ (.A(_05920_),
    .B(_05923_),
    .X(_05925_));
 sky130_fd_sc_hd__or3_1 _11303_ (.A(_03841_),
    .B(_05924_),
    .C(_05925_),
    .X(_05926_));
 sky130_fd_sc_hd__a21bo_1 _11304_ (.A1(_04959_),
    .A2(_05838_),
    .B1_N(_05926_),
    .X(_05927_));
 sky130_fd_sc_hd__clkbuf_2 _11305_ (.A(_05927_),
    .X(net208));
 sky130_fd_sc_hd__buf_2 _11306_ (.A(_05898_),
    .X(_05928_));
 sky130_fd_sc_hd__mux2_2 _11307_ (.A0(\reg_next_pc[25] ),
    .A1(\reg_out[25] ),
    .S(_05928_),
    .X(_05929_));
 sky130_fd_sc_hd__xor2_1 _11308_ (.A(_05925_),
    .B(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__mux2_1 _11309_ (.A0(_05013_),
    .A1(_05930_),
    .S(_03219_),
    .X(_05931_));
 sky130_fd_sc_hd__clkbuf_2 _11310_ (.A(_05931_),
    .X(net209));
 sky130_fd_sc_hd__mux2_2 _11311_ (.A0(\reg_next_pc[26] ),
    .A1(\reg_out[26] ),
    .S(_05928_),
    .X(_05932_));
 sky130_fd_sc_hd__a21oi_1 _11312_ (.A1(_05925_),
    .A2(_05929_),
    .B1(_05932_),
    .Y(_05933_));
 sky130_fd_sc_hd__and3_1 _11313_ (.A(_05925_),
    .B(_05929_),
    .C(_05932_),
    .X(_05934_));
 sky130_fd_sc_hd__or3_1 _11314_ (.A(_03841_),
    .B(_05933_),
    .C(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__a21bo_1 _11315_ (.A1(_05044_),
    .A2(_05838_),
    .B1_N(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__clkbuf_2 _11316_ (.A(_05936_),
    .X(net210));
 sky130_fd_sc_hd__mux2_2 _11317_ (.A0(\reg_next_pc[27] ),
    .A1(\reg_out[27] ),
    .S(_05928_),
    .X(_05937_));
 sky130_fd_sc_hd__and4_1 _11318_ (.A(_05925_),
    .B(_05929_),
    .C(_05932_),
    .D(_05937_),
    .X(_05938_));
 sky130_fd_sc_hd__o21ba_1 _11319_ (.A1(_05934_),
    .A2(_05937_),
    .B1_N(_05938_),
    .X(_05939_));
 sky130_fd_sc_hd__mux2_1 _11320_ (.A0(_05076_),
    .A1(_05939_),
    .S(_03219_),
    .X(_05940_));
 sky130_fd_sc_hd__clkbuf_2 _11321_ (.A(_05940_),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_4 _11322_ (.A(_05909_),
    .X(_05941_));
 sky130_fd_sc_hd__or2_1 _11323_ (.A(\reg_next_pc[28] ),
    .B(_05928_),
    .X(_05942_));
 sky130_fd_sc_hd__o21a_1 _11324_ (.A1(\reg_out[28] ),
    .A2(_05941_),
    .B1(_05942_),
    .X(_05943_));
 sky130_fd_sc_hd__xor2_1 _11325_ (.A(_05938_),
    .B(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__mux2_1 _11326_ (.A0(_05086_),
    .A1(_05944_),
    .S(_03219_),
    .X(_05945_));
 sky130_fd_sc_hd__clkbuf_2 _11327_ (.A(_05945_),
    .X(net212));
 sky130_fd_sc_hd__and2_1 _11328_ (.A(_05938_),
    .B(_05943_),
    .X(_05946_));
 sky130_fd_sc_hd__or2_1 _11329_ (.A(\reg_next_pc[29] ),
    .B(_05928_),
    .X(_05947_));
 sky130_fd_sc_hd__o21a_2 _11330_ (.A1(\reg_out[29] ),
    .A2(_05941_),
    .B1(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__xor2_1 _11331_ (.A(_05946_),
    .B(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__mux2_1 _11332_ (.A0(_05143_),
    .A1(_05949_),
    .S(_03219_),
    .X(_05950_));
 sky130_fd_sc_hd__buf_2 _11333_ (.A(_05950_),
    .X(net213));
 sky130_fd_sc_hd__or2_1 _11334_ (.A(\reg_next_pc[30] ),
    .B(_05928_),
    .X(_05951_));
 sky130_fd_sc_hd__o21a_1 _11335_ (.A1(\reg_out[30] ),
    .A2(_05941_),
    .B1(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__a21oi_1 _11336_ (.A1(_05946_),
    .A2(_05948_),
    .B1(_05952_),
    .Y(_05953_));
 sky130_fd_sc_hd__and3_1 _11337_ (.A(_05946_),
    .B(_05948_),
    .C(_05952_),
    .X(_05954_));
 sky130_fd_sc_hd__or3_1 _11338_ (.A(_03229_),
    .B(_05953_),
    .C(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__a21bo_1 _11339_ (.A1(_05174_),
    .A2(_05838_),
    .B1_N(_05955_),
    .X(_05956_));
 sky130_fd_sc_hd__buf_2 _11340_ (.A(_05956_),
    .X(net215));
 sky130_fd_sc_hd__mux2_2 _11341_ (.A0(\reg_next_pc[31] ),
    .A1(\reg_out[31] ),
    .S(_05928_),
    .X(_05957_));
 sky130_fd_sc_hd__xor2_1 _11342_ (.A(_05954_),
    .B(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__mux2_1 _11343_ (.A0(_05205_),
    .A1(_05958_),
    .S(_03219_),
    .X(_05959_));
 sky130_fd_sc_hd__clkbuf_2 _11344_ (.A(_05959_),
    .X(net216));
 sky130_fd_sc_hd__buf_2 _11345_ (.A(_03228_),
    .X(_05960_));
 sky130_fd_sc_hd__and3_1 _11346_ (.A(_03739_),
    .B(_03853_),
    .C(_03926_),
    .X(_05961_));
 sky130_fd_sc_hd__a31o_1 _11347_ (.A1(_03748_),
    .A2(_03879_),
    .A3(_03844_),
    .B1(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__nand2_1 _11348_ (.A(_03748_),
    .B(_03790_),
    .Y(_05963_));
 sky130_fd_sc_hd__a221o_1 _11349_ (.A1(_03891_),
    .A2(_03767_),
    .B1(_03770_),
    .B2(_03736_),
    .C1(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__or4_1 _11350_ (.A(_03787_),
    .B(_03762_),
    .C(_03770_),
    .D(_03736_),
    .X(_05965_));
 sky130_fd_sc_hd__nand3b_1 _11351_ (.A_N(_03948_),
    .B(_05964_),
    .C(_05965_),
    .Y(_05966_));
 sky130_fd_sc_hd__or2_1 _11352_ (.A(_05962_),
    .B(_05966_),
    .X(_05967_));
 sky130_fd_sc_hd__and3_1 _11353_ (.A(_05960_),
    .B(_03864_),
    .C(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__buf_2 _11354_ (.A(_03215_),
    .X(_05969_));
 sky130_fd_sc_hd__nand2_4 _11355_ (.A(_03199_),
    .B(_03310_),
    .Y(_05970_));
 sky130_fd_sc_hd__a21oi_1 _11356_ (.A1(_05969_),
    .A2(_03851_),
    .B1(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__inv_2 _11357_ (.A(_05971_),
    .Y(_05972_));
 sky130_fd_sc_hd__o22a_1 _11358_ (.A1(\cpuregs.raddr2[0] ),
    .A2(_03636_),
    .B1(_05968_),
    .B2(_05972_),
    .X(_00084_));
 sky130_fd_sc_hd__buf_2 _11359_ (.A(_05970_),
    .X(_05973_));
 sky130_fd_sc_hd__buf_2 _11360_ (.A(_05973_),
    .X(_05974_));
 sky130_fd_sc_hd__a21o_1 _11361_ (.A1(_05969_),
    .A2(_03874_),
    .B1(_05967_),
    .X(_05975_));
 sky130_fd_sc_hd__nand2_2 _11362_ (.A(_03228_),
    .B(_03633_),
    .Y(_05976_));
 sky130_fd_sc_hd__nor2_1 _11363_ (.A(_03979_),
    .B(_05976_),
    .Y(_05977_));
 sky130_fd_sc_hd__a31o_1 _11364_ (.A1(_05969_),
    .A2(_03634_),
    .A3(_03874_),
    .B1(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__a22o_1 _11365_ (.A1(\cpuregs.raddr2[1] ),
    .A2(_05974_),
    .B1(_05975_),
    .B2(_05978_),
    .X(_00085_));
 sky130_fd_sc_hd__and3_1 _11366_ (.A(_03783_),
    .B(_03213_),
    .C(_03876_),
    .X(_05979_));
 sky130_fd_sc_hd__or2_1 _11367_ (.A(_05967_),
    .B(_05979_),
    .X(_05980_));
 sky130_fd_sc_hd__nor2_1 _11368_ (.A(_03215_),
    .B(_05970_),
    .Y(_05981_));
 sky130_fd_sc_hd__a22o_1 _11369_ (.A1(_03885_),
    .A2(_05981_),
    .B1(_05979_),
    .B2(_03634_),
    .X(_05982_));
 sky130_fd_sc_hd__a22o_1 _11370_ (.A1(\cpuregs.raddr2[2] ),
    .A2(_05974_),
    .B1(_05980_),
    .B2(_05982_),
    .X(_00086_));
 sky130_fd_sc_hd__clkbuf_4 _11371_ (.A(_05970_),
    .X(_05983_));
 sky130_fd_sc_hd__o211a_1 _11372_ (.A1(_03895_),
    .A2(_05962_),
    .B1(_05967_),
    .C1(_05981_),
    .X(_05984_));
 sky130_fd_sc_hd__and3_1 _11373_ (.A(_05969_),
    .B(_03634_),
    .C(_03889_),
    .X(_05985_));
 sky130_fd_sc_hd__a211o_1 _11374_ (.A1(\cpuregs.raddr2[3] ),
    .A2(_05983_),
    .B1(_05984_),
    .C1(_05985_),
    .X(_00087_));
 sky130_fd_sc_hd__and3_1 _11375_ (.A(_05960_),
    .B(_03878_),
    .C(_05966_),
    .X(_05986_));
 sky130_fd_sc_hd__clkbuf_4 _11376_ (.A(_05970_),
    .X(_05987_));
 sky130_fd_sc_hd__a21o_1 _11377_ (.A1(_05969_),
    .A2(_03900_),
    .B1(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__o22a_1 _11378_ (.A1(\cpuregs.raddr2[4] ),
    .A2(_03636_),
    .B1(_05986_),
    .B2(_05988_),
    .X(_00088_));
 sky130_fd_sc_hd__nor2_1 _11379_ (.A(_03916_),
    .B(_03777_),
    .Y(_05989_));
 sky130_fd_sc_hd__or3_2 _11380_ (.A(_03787_),
    .B(_03770_),
    .C(_05989_),
    .X(_05990_));
 sky130_fd_sc_hd__inv_2 _11381_ (.A(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__o21ai_1 _11382_ (.A1(_03816_),
    .A2(_03736_),
    .B1(_03853_),
    .Y(_05992_));
 sky130_fd_sc_hd__or4_1 _11383_ (.A(_03781_),
    .B(_03789_),
    .C(_03768_),
    .D(_03736_),
    .X(_05993_));
 sky130_fd_sc_hd__o21ai_2 _11384_ (.A1(_03789_),
    .A2(_05992_),
    .B1(_05993_),
    .Y(_05994_));
 sky130_fd_sc_hd__a21o_1 _11385_ (.A1(_03739_),
    .A2(_03923_),
    .B1(_05994_),
    .X(_05995_));
 sky130_fd_sc_hd__or4_1 _11386_ (.A(_03845_),
    .B(_03971_),
    .C(_05991_),
    .D(_05995_),
    .X(_05996_));
 sky130_fd_sc_hd__or3_1 _11387_ (.A(_03228_),
    .B(_03979_),
    .C(_03814_),
    .X(_05997_));
 sky130_fd_sc_hd__or3_1 _11388_ (.A(_03800_),
    .B(_03804_),
    .C(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__or3_1 _11389_ (.A(_03756_),
    .B(_03994_),
    .C(_04000_),
    .X(_05999_));
 sky130_fd_sc_hd__or2_1 _11390_ (.A(_03954_),
    .B(_03987_),
    .X(_06000_));
 sky130_fd_sc_hd__or3b_1 _11391_ (.A(_03977_),
    .B(_06000_),
    .C_N(_03965_),
    .X(_06001_));
 sky130_fd_sc_hd__or3_1 _11392_ (.A(_05998_),
    .B(_05999_),
    .C(_06001_),
    .X(_06002_));
 sky130_fd_sc_hd__nand2_2 _11393_ (.A(_03633_),
    .B(_06002_),
    .Y(_06003_));
 sky130_fd_sc_hd__or2_1 _11394_ (.A(_03781_),
    .B(_06003_),
    .X(_06004_));
 sky130_fd_sc_hd__a22o_1 _11395_ (.A1(_03822_),
    .A2(_05996_),
    .B1(_06004_),
    .B2(_05976_),
    .X(_06005_));
 sky130_fd_sc_hd__o21a_1 _11396_ (.A1(\cpuregs.raddr1[0] ),
    .A2(_03636_),
    .B1(_06005_),
    .X(_00089_));
 sky130_fd_sc_hd__clkbuf_4 _11397_ (.A(_03635_),
    .X(_06006_));
 sky130_fd_sc_hd__o22a_1 _11398_ (.A1(_03867_),
    .A2(_03923_),
    .B1(_03971_),
    .B2(_03880_),
    .X(_06007_));
 sky130_fd_sc_hd__a21oi_1 _11399_ (.A1(_03767_),
    .A2(_03833_),
    .B1(_03947_),
    .Y(_06008_));
 sky130_fd_sc_hd__a21o_1 _11400_ (.A1(_03816_),
    .A2(_03916_),
    .B1(_03902_),
    .X(_06009_));
 sky130_fd_sc_hd__or3b_1 _11401_ (.A(_03770_),
    .B(_05989_),
    .C_N(_03867_),
    .X(_06010_));
 sky130_fd_sc_hd__o21ai_1 _11402_ (.A1(_03844_),
    .A2(_03923_),
    .B1(_03867_),
    .Y(_06011_));
 sky130_fd_sc_hd__a31o_1 _11403_ (.A1(_06009_),
    .A2(_06010_),
    .A3(_06011_),
    .B1(_03750_),
    .X(_06012_));
 sky130_fd_sc_hd__or4b_1 _11404_ (.A(_05976_),
    .B(_06007_),
    .C(_06008_),
    .D_N(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__a21o_1 _11405_ (.A1(_03867_),
    .A2(_05994_),
    .B1(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__or3_1 _11406_ (.A(_05960_),
    .B(_03910_),
    .C(_06003_),
    .X(_06015_));
 sky130_fd_sc_hd__o211a_1 _11407_ (.A1(\cpuregs.raddr1[1] ),
    .A2(_06006_),
    .B1(_06014_),
    .C1(_06015_),
    .X(_00090_));
 sky130_fd_sc_hd__clkbuf_4 _11408_ (.A(_05981_),
    .X(_06016_));
 sky130_fd_sc_hd__nand2_1 _11409_ (.A(_05969_),
    .B(_03913_),
    .Y(_06017_));
 sky130_fd_sc_hd__a2bb2o_1 _11410_ (.A1_N(_06003_),
    .A2_N(_06017_),
    .B1(\cpuregs.raddr1[2] ),
    .B2(_05973_),
    .X(_06018_));
 sky130_fd_sc_hd__a31o_1 _11411_ (.A1(_03826_),
    .A2(_06016_),
    .A3(_05996_),
    .B1(_06018_),
    .X(_00091_));
 sky130_fd_sc_hd__and3_1 _11412_ (.A(_03783_),
    .B(_03892_),
    .C(_03923_),
    .X(_06019_));
 sky130_fd_sc_hd__o41a_1 _11413_ (.A1(_03845_),
    .A2(_03971_),
    .A3(_05991_),
    .A4(_06019_),
    .B1(_05960_),
    .X(_06020_));
 sky130_fd_sc_hd__and3_1 _11414_ (.A(_03215_),
    .B(_03918_),
    .C(_06002_),
    .X(_06021_));
 sky130_fd_sc_hd__a211o_1 _11415_ (.A1(_03892_),
    .A2(_05994_),
    .B1(_06021_),
    .C1(_05973_),
    .X(_06022_));
 sky130_fd_sc_hd__o22a_1 _11416_ (.A1(\cpuregs.raddr1[3] ),
    .A2(_06006_),
    .B1(_06020_),
    .B2(_06022_),
    .X(_00092_));
 sky130_fd_sc_hd__nor2_1 _11417_ (.A(_03215_),
    .B(_03879_),
    .Y(_06023_));
 sky130_fd_sc_hd__inv_2 _11418_ (.A(_06003_),
    .Y(_06024_));
 sky130_fd_sc_hd__a32o_1 _11419_ (.A1(_05969_),
    .A2(_03920_),
    .A3(_06024_),
    .B1(_05973_),
    .B2(\cpuregs.raddr1[4] ),
    .X(_06025_));
 sky130_fd_sc_hd__a41o_1 _11420_ (.A1(_06006_),
    .A2(_03763_),
    .A3(_05995_),
    .A4(_06023_),
    .B1(_06025_),
    .X(_00093_));
 sky130_fd_sc_hd__clkbuf_8 _11421_ (.A(_03305_),
    .X(_06026_));
 sky130_fd_sc_hd__or2_1 _11422_ (.A(\irq_pending[1] ),
    .B(_03308_),
    .X(_06027_));
 sky130_fd_sc_hd__or3b_1 _11423_ (.A(_03412_),
    .B(\irq_mask[1] ),
    .C_N(\irq_pending[1] ),
    .X(_06028_));
 sky130_fd_sc_hd__a31o_1 _11424_ (.A1(_06026_),
    .A2(_06027_),
    .A3(_06028_),
    .B1(net12),
    .X(_00012_));
 sky130_fd_sc_hd__buf_2 _11425_ (.A(_03305_),
    .X(_06029_));
 sky130_fd_sc_hd__clkbuf_2 _11426_ (.A(_03412_),
    .X(_06030_));
 sky130_fd_sc_hd__or2_1 _11427_ (.A(\irq_mask[3] ),
    .B(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__a31o_1 _11428_ (.A1(_06029_),
    .A2(\irq_pending[3] ),
    .A3(_06031_),
    .B1(net26),
    .X(_00026_));
 sky130_fd_sc_hd__or2_1 _11429_ (.A(\irq_mask[4] ),
    .B(_06030_),
    .X(_06032_));
 sky130_fd_sc_hd__a31o_1 _11430_ (.A1(_06029_),
    .A2(\irq_pending[4] ),
    .A3(_06032_),
    .B1(net27),
    .X(_00027_));
 sky130_fd_sc_hd__or2_1 _11431_ (.A(\irq_mask[5] ),
    .B(_06030_),
    .X(_06033_));
 sky130_fd_sc_hd__a31o_1 _11432_ (.A1(_06029_),
    .A2(\irq_pending[5] ),
    .A3(_06033_),
    .B1(net28),
    .X(_00028_));
 sky130_fd_sc_hd__or2_1 _11433_ (.A(\irq_mask[6] ),
    .B(_06030_),
    .X(_06034_));
 sky130_fd_sc_hd__a31o_1 _11434_ (.A1(_06029_),
    .A2(\irq_pending[6] ),
    .A3(_06034_),
    .B1(net29),
    .X(_00029_));
 sky130_fd_sc_hd__or2_1 _11435_ (.A(\irq_mask[7] ),
    .B(_06030_),
    .X(_06035_));
 sky130_fd_sc_hd__a31o_1 _11436_ (.A1(_06029_),
    .A2(\irq_pending[7] ),
    .A3(_06035_),
    .B1(net30),
    .X(_00030_));
 sky130_fd_sc_hd__or2_1 _11437_ (.A(\irq_mask[8] ),
    .B(_06030_),
    .X(_06036_));
 sky130_fd_sc_hd__a31o_1 _11438_ (.A1(_06029_),
    .A2(\irq_pending[8] ),
    .A3(_06036_),
    .B1(net31),
    .X(_00031_));
 sky130_fd_sc_hd__or2_1 _11439_ (.A(\irq_mask[9] ),
    .B(_06030_),
    .X(_06037_));
 sky130_fd_sc_hd__a31o_1 _11440_ (.A1(_06029_),
    .A2(\irq_pending[9] ),
    .A3(_06037_),
    .B1(net32),
    .X(_00032_));
 sky130_fd_sc_hd__or2_1 _11441_ (.A(\irq_mask[10] ),
    .B(_06030_),
    .X(_06038_));
 sky130_fd_sc_hd__a31o_1 _11442_ (.A1(_06029_),
    .A2(\irq_pending[10] ),
    .A3(_06038_),
    .B1(net2),
    .X(_00002_));
 sky130_fd_sc_hd__or2_1 _11443_ (.A(\irq_mask[11] ),
    .B(_06030_),
    .X(_06039_));
 sky130_fd_sc_hd__a31o_1 _11444_ (.A1(_06029_),
    .A2(\irq_pending[11] ),
    .A3(_06039_),
    .B1(net3),
    .X(_00003_));
 sky130_fd_sc_hd__or2_1 _11445_ (.A(\irq_mask[12] ),
    .B(_06030_),
    .X(_06040_));
 sky130_fd_sc_hd__a31o_1 _11446_ (.A1(_06029_),
    .A2(\irq_pending[12] ),
    .A3(_06040_),
    .B1(net4),
    .X(_00004_));
 sky130_fd_sc_hd__clkbuf_4 _11447_ (.A(_03305_),
    .X(_06041_));
 sky130_fd_sc_hd__buf_2 _11448_ (.A(_03412_),
    .X(_06042_));
 sky130_fd_sc_hd__or2_1 _11449_ (.A(\irq_mask[13] ),
    .B(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__a31o_1 _11450_ (.A1(_06041_),
    .A2(\irq_pending[13] ),
    .A3(_06043_),
    .B1(net5),
    .X(_00005_));
 sky130_fd_sc_hd__or2_1 _11451_ (.A(\irq_mask[14] ),
    .B(_06042_),
    .X(_06044_));
 sky130_fd_sc_hd__a31o_1 _11452_ (.A1(_06041_),
    .A2(\irq_pending[14] ),
    .A3(_06044_),
    .B1(net6),
    .X(_00006_));
 sky130_fd_sc_hd__or2_1 _11453_ (.A(\irq_mask[15] ),
    .B(_06042_),
    .X(_06045_));
 sky130_fd_sc_hd__a31o_1 _11454_ (.A1(_06041_),
    .A2(\irq_pending[15] ),
    .A3(_06045_),
    .B1(net7),
    .X(_00007_));
 sky130_fd_sc_hd__or2_1 _11455_ (.A(\irq_mask[16] ),
    .B(_06042_),
    .X(_06046_));
 sky130_fd_sc_hd__a31o_1 _11456_ (.A1(_06041_),
    .A2(\irq_pending[16] ),
    .A3(_06046_),
    .B1(net8),
    .X(_00008_));
 sky130_fd_sc_hd__or2_1 _11457_ (.A(\irq_mask[17] ),
    .B(_06042_),
    .X(_06047_));
 sky130_fd_sc_hd__a31o_1 _11458_ (.A1(_06041_),
    .A2(\irq_pending[17] ),
    .A3(_06047_),
    .B1(net9),
    .X(_00009_));
 sky130_fd_sc_hd__or2_1 _11459_ (.A(\irq_mask[18] ),
    .B(_06042_),
    .X(_06048_));
 sky130_fd_sc_hd__a31o_1 _11460_ (.A1(_06041_),
    .A2(\irq_pending[18] ),
    .A3(_06048_),
    .B1(net10),
    .X(_00010_));
 sky130_fd_sc_hd__or2_1 _11461_ (.A(\irq_mask[19] ),
    .B(_06042_),
    .X(_06049_));
 sky130_fd_sc_hd__a31o_1 _11462_ (.A1(_06041_),
    .A2(\irq_pending[19] ),
    .A3(_06049_),
    .B1(net11),
    .X(_00011_));
 sky130_fd_sc_hd__or2_1 _11463_ (.A(\irq_mask[20] ),
    .B(_06042_),
    .X(_06050_));
 sky130_fd_sc_hd__a31o_1 _11464_ (.A1(_06041_),
    .A2(\irq_pending[20] ),
    .A3(_06050_),
    .B1(net13),
    .X(_00013_));
 sky130_fd_sc_hd__or2_1 _11465_ (.A(\irq_mask[21] ),
    .B(_06042_),
    .X(_06051_));
 sky130_fd_sc_hd__a31o_1 _11466_ (.A1(_06041_),
    .A2(\irq_pending[21] ),
    .A3(_06051_),
    .B1(net14),
    .X(_00014_));
 sky130_fd_sc_hd__or2_1 _11467_ (.A(\irq_mask[22] ),
    .B(_06042_),
    .X(_06052_));
 sky130_fd_sc_hd__a31o_1 _11468_ (.A1(_06041_),
    .A2(\irq_pending[22] ),
    .A3(_06052_),
    .B1(net15),
    .X(_00015_));
 sky130_fd_sc_hd__clkbuf_8 _11469_ (.A(_03277_),
    .X(_06053_));
 sky130_fd_sc_hd__clkbuf_4 _11470_ (.A(_06053_),
    .X(_06054_));
 sky130_fd_sc_hd__or2_1 _11471_ (.A(\irq_mask[23] ),
    .B(_03428_),
    .X(_06055_));
 sky130_fd_sc_hd__a31o_1 _11472_ (.A1(_06054_),
    .A2(\irq_pending[23] ),
    .A3(_06055_),
    .B1(net16),
    .X(_00016_));
 sky130_fd_sc_hd__or2_1 _11473_ (.A(\irq_mask[24] ),
    .B(_03428_),
    .X(_06056_));
 sky130_fd_sc_hd__a31o_1 _11474_ (.A1(_06054_),
    .A2(\irq_pending[24] ),
    .A3(_06056_),
    .B1(net17),
    .X(_00017_));
 sky130_fd_sc_hd__or2_1 _11475_ (.A(\irq_mask[25] ),
    .B(_03428_),
    .X(_06057_));
 sky130_fd_sc_hd__a31o_1 _11476_ (.A1(_06054_),
    .A2(\irq_pending[25] ),
    .A3(_06057_),
    .B1(net18),
    .X(_00018_));
 sky130_fd_sc_hd__or2_1 _11477_ (.A(\irq_mask[26] ),
    .B(_03428_),
    .X(_06058_));
 sky130_fd_sc_hd__a31o_1 _11478_ (.A1(_06054_),
    .A2(\irq_pending[26] ),
    .A3(_06058_),
    .B1(net19),
    .X(_00019_));
 sky130_fd_sc_hd__or2_1 _11479_ (.A(\irq_mask[27] ),
    .B(_03428_),
    .X(_06059_));
 sky130_fd_sc_hd__a31o_1 _11480_ (.A1(_06054_),
    .A2(\irq_pending[27] ),
    .A3(_06059_),
    .B1(net20),
    .X(_00020_));
 sky130_fd_sc_hd__or2_1 _11481_ (.A(\irq_mask[28] ),
    .B(_03428_),
    .X(_06060_));
 sky130_fd_sc_hd__a31o_1 _11482_ (.A1(_06054_),
    .A2(\irq_pending[28] ),
    .A3(_06060_),
    .B1(net21),
    .X(_00021_));
 sky130_fd_sc_hd__or2_1 _11483_ (.A(\irq_mask[29] ),
    .B(_03428_),
    .X(_06061_));
 sky130_fd_sc_hd__a31o_1 _11484_ (.A1(_06054_),
    .A2(\irq_pending[29] ),
    .A3(_06061_),
    .B1(net22),
    .X(_00022_));
 sky130_fd_sc_hd__or2_1 _11485_ (.A(\irq_mask[30] ),
    .B(_03428_),
    .X(_06062_));
 sky130_fd_sc_hd__a31o_1 _11486_ (.A1(_06054_),
    .A2(\irq_pending[30] ),
    .A3(_06062_),
    .B1(net24),
    .X(_00024_));
 sky130_fd_sc_hd__or2_1 _11487_ (.A(\irq_mask[31] ),
    .B(_03428_),
    .X(_06063_));
 sky130_fd_sc_hd__a31o_1 _11488_ (.A1(_06054_),
    .A2(\irq_pending[31] ),
    .A3(_06063_),
    .B1(net25),
    .X(_00025_));
 sky130_fd_sc_hd__and3b_1 _11489_ (.A_N(net65),
    .B(net262),
    .C(_03305_),
    .X(_06064_));
 sky130_fd_sc_hd__clkbuf_1 _11490_ (.A(_06064_),
    .X(_00094_));
 sky130_fd_sc_hd__nor2b_2 _11491_ (.A(latched_branch),
    .B_N(latched_store),
    .Y(_06065_));
 sky130_fd_sc_hd__clkbuf_4 _11492_ (.A(_06065_),
    .X(_06066_));
 sky130_fd_sc_hd__clkbuf_4 _11493_ (.A(latched_stalu),
    .X(_06067_));
 sky130_fd_sc_hd__clkbuf_4 _11494_ (.A(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__buf_4 _11495_ (.A(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__mux2_1 _11496_ (.A0(\reg_out[0] ),
    .A1(\alu_out_q[0] ),
    .S(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__clkbuf_4 _11497_ (.A(\irq_state[0] ),
    .X(_06071_));
 sky130_fd_sc_hd__clkbuf_4 _11498_ (.A(\irq_state[1] ),
    .X(_06072_));
 sky130_fd_sc_hd__a22o_1 _11499_ (.A1(_06071_),
    .A2(latched_compr),
    .B1(_03338_),
    .B2(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__nor2_1 _11500_ (.A(_03195_),
    .B(_06065_),
    .Y(_06074_));
 sky130_fd_sc_hd__clkbuf_4 _11501_ (.A(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__o21a_1 _11502_ (.A1(_06071_),
    .A2(_06075_),
    .B1(\reg_next_pc[0] ),
    .X(_06076_));
 sky130_fd_sc_hd__a211o_2 _11503_ (.A1(_06066_),
    .A2(_06070_),
    .B1(_06073_),
    .C1(_06076_),
    .X(_06077_));
 sky130_fd_sc_hd__buf_2 _11504_ (.A(_06077_),
    .X(_06078_));
 sky130_fd_sc_hd__and2b_1 _11505_ (.A_N(\cpuregs.waddr[0] ),
    .B(\cpuregs.waddr[1] ),
    .X(_06079_));
 sky130_fd_sc_hd__buf_4 _11506_ (.A(_06079_),
    .X(_06080_));
 sky130_fd_sc_hd__clkbuf_4 _11507_ (.A(\cpuregs.waddr[4] ),
    .X(_06081_));
 sky130_fd_sc_hd__clkbuf_4 _11508_ (.A(\cpuregs.waddr[3] ),
    .X(_06082_));
 sky130_fd_sc_hd__o31a_4 _11509_ (.A1(latched_branch),
    .A2(latched_store),
    .A3(_03195_),
    .B1(_03293_),
    .X(_06083_));
 sky130_fd_sc_hd__and4bb_2 _11510_ (.A_N(\cpuregs.waddr[2] ),
    .B_N(_06081_),
    .C(_06082_),
    .D(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__nand2_2 _11511_ (.A(_06080_),
    .B(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__buf_6 _11512_ (.A(_06085_),
    .X(_06086_));
 sky130_fd_sc_hd__mux2_1 _11513_ (.A0(_06078_),
    .A1(\cpuregs.regs[10][0] ),
    .S(_06086_),
    .X(_06087_));
 sky130_fd_sc_hd__clkbuf_1 _11514_ (.A(_06087_),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _11515_ (.A0(\reg_out[1] ),
    .A1(\alu_out_q[1] ),
    .S(latched_stalu),
    .X(_06088_));
 sky130_fd_sc_hd__a22o_1 _11516_ (.A1(_06071_),
    .A2(\reg_next_pc[1] ),
    .B1(_03351_),
    .B2(_06072_),
    .X(_06089_));
 sky130_fd_sc_hd__nand2b_1 _11517_ (.A_N(\reg_pc[1] ),
    .B(latched_compr),
    .Y(_06090_));
 sky130_fd_sc_hd__or2b_1 _11518_ (.A(latched_compr),
    .B_N(\reg_pc[1] ),
    .X(_06091_));
 sky130_fd_sc_hd__or2_1 _11519_ (.A(_03195_),
    .B(_06065_),
    .X(_06092_));
 sky130_fd_sc_hd__clkbuf_4 _11520_ (.A(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__a21oi_1 _11521_ (.A1(_06090_),
    .A2(_06091_),
    .B1(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__a211o_4 _11522_ (.A1(_06066_),
    .A2(_06088_),
    .B1(_06089_),
    .C1(_06094_),
    .X(_06095_));
 sky130_fd_sc_hd__buf_2 _11523_ (.A(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__mux2_1 _11524_ (.A0(_06096_),
    .A1(\cpuregs.regs[10][1] ),
    .S(_06086_),
    .X(_06097_));
 sky130_fd_sc_hd__clkbuf_1 _11525_ (.A(_06097_),
    .X(_00096_));
 sky130_fd_sc_hd__clkbuf_4 _11526_ (.A(_06065_),
    .X(_06098_));
 sky130_fd_sc_hd__mux2_1 _11527_ (.A0(\reg_out[2] ),
    .A1(\alu_out_q[2] ),
    .S(latched_stalu),
    .X(_06099_));
 sky130_fd_sc_hd__and2_1 _11528_ (.A(_06098_),
    .B(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__buf_2 _11529_ (.A(_06074_),
    .X(_06101_));
 sky130_fd_sc_hd__a221o_1 _11530_ (.A1(_06071_),
    .A2(\reg_next_pc[2] ),
    .B1(_03326_),
    .B2(_06072_),
    .C1(_06101_),
    .X(_06102_));
 sky130_fd_sc_hd__xor2_1 _11531_ (.A(\reg_pc[2] ),
    .B(_06090_),
    .X(_06103_));
 sky130_fd_sc_hd__o22a_2 _11532_ (.A1(_06100_),
    .A2(_06102_),
    .B1(_06103_),
    .B2(_06093_),
    .X(_06104_));
 sky130_fd_sc_hd__buf_2 _11533_ (.A(_06104_),
    .X(_06105_));
 sky130_fd_sc_hd__mux2_1 _11534_ (.A0(_06105_),
    .A1(\cpuregs.regs[10][2] ),
    .S(_06086_),
    .X(_06106_));
 sky130_fd_sc_hd__clkbuf_1 _11535_ (.A(_06106_),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _11536_ (.A0(\reg_out[3] ),
    .A1(\alu_out_q[3] ),
    .S(latched_stalu),
    .X(_06107_));
 sky130_fd_sc_hd__and2_1 _11537_ (.A(_06098_),
    .B(_06107_),
    .X(_06108_));
 sky130_fd_sc_hd__a221o_1 _11538_ (.A1(\irq_state[0] ),
    .A2(\reg_next_pc[3] ),
    .B1(_03344_),
    .B2(_06072_),
    .C1(_06101_),
    .X(_06109_));
 sky130_fd_sc_hd__and3_1 _11539_ (.A(\reg_pc[3] ),
    .B(\reg_pc[2] ),
    .C(_06090_),
    .X(_06110_));
 sky130_fd_sc_hd__a21oi_1 _11540_ (.A1(\reg_pc[2] ),
    .A2(_06090_),
    .B1(\reg_pc[3] ),
    .Y(_06111_));
 sky130_fd_sc_hd__nor2_1 _11541_ (.A(_06110_),
    .B(_06111_),
    .Y(_06112_));
 sky130_fd_sc_hd__o22a_2 _11542_ (.A1(_06108_),
    .A2(_06109_),
    .B1(_06112_),
    .B2(_06093_),
    .X(_06113_));
 sky130_fd_sc_hd__buf_2 _11543_ (.A(_06113_),
    .X(_06114_));
 sky130_fd_sc_hd__mux2_1 _11544_ (.A0(_06114_),
    .A1(\cpuregs.regs[10][3] ),
    .S(_06086_),
    .X(_06115_));
 sky130_fd_sc_hd__clkbuf_1 _11545_ (.A(_06115_),
    .X(_00098_));
 sky130_fd_sc_hd__clkbuf_4 _11546_ (.A(_06071_),
    .X(_06116_));
 sky130_fd_sc_hd__mux2_1 _11547_ (.A0(\reg_out[4] ),
    .A1(\alu_out_q[4] ),
    .S(latched_stalu),
    .X(_06117_));
 sky130_fd_sc_hd__buf_2 _11548_ (.A(_06074_),
    .X(_06118_));
 sky130_fd_sc_hd__a221o_1 _11549_ (.A1(_06072_),
    .A2(_03327_),
    .B1(_06098_),
    .B2(_06117_),
    .C1(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__a21oi_2 _11550_ (.A1(_06116_),
    .A2(\reg_next_pc[4] ),
    .B1(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__and2_1 _11551_ (.A(\reg_pc[4] ),
    .B(_06110_),
    .X(_06121_));
 sky130_fd_sc_hd__nor2_1 _11552_ (.A(\reg_pc[4] ),
    .B(_06110_),
    .Y(_06122_));
 sky130_fd_sc_hd__o21a_1 _11553_ (.A1(_06121_),
    .A2(_06122_),
    .B1(_06075_),
    .X(_06123_));
 sky130_fd_sc_hd__nor2_4 _11554_ (.A(_06120_),
    .B(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__buf_2 _11555_ (.A(_06124_),
    .X(_06125_));
 sky130_fd_sc_hd__mux2_1 _11556_ (.A0(_06125_),
    .A1(\cpuregs.regs[10][4] ),
    .S(_06086_),
    .X(_06126_));
 sky130_fd_sc_hd__clkbuf_1 _11557_ (.A(_06126_),
    .X(_00099_));
 sky130_fd_sc_hd__xnor2_1 _11558_ (.A(\reg_pc[5] ),
    .B(_06121_),
    .Y(_06127_));
 sky130_fd_sc_hd__mux2_1 _11559_ (.A0(\reg_out[5] ),
    .A1(\alu_out_q[5] ),
    .S(_06067_),
    .X(_06128_));
 sky130_fd_sc_hd__a221o_1 _11560_ (.A1(\irq_state[1] ),
    .A2(_03322_),
    .B1(_06098_),
    .B2(_06128_),
    .C1(_06074_),
    .X(_06129_));
 sky130_fd_sc_hd__a21oi_1 _11561_ (.A1(_06071_),
    .A2(\reg_next_pc[5] ),
    .B1(_06129_),
    .Y(_06130_));
 sky130_fd_sc_hd__a21oi_2 _11562_ (.A1(_06075_),
    .A2(_06127_),
    .B1(_06130_),
    .Y(_06131_));
 sky130_fd_sc_hd__buf_2 _11563_ (.A(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__mux2_1 _11564_ (.A0(_06132_),
    .A1(\cpuregs.regs[10][5] ),
    .S(_06086_),
    .X(_06133_));
 sky130_fd_sc_hd__clkbuf_1 _11565_ (.A(_06133_),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _11566_ (.A0(\reg_out[6] ),
    .A1(\alu_out_q[6] ),
    .S(latched_stalu),
    .X(_06134_));
 sky130_fd_sc_hd__a221o_1 _11567_ (.A1(_06072_),
    .A2(_03321_),
    .B1(_06098_),
    .B2(_06134_),
    .C1(_06118_),
    .X(_06135_));
 sky130_fd_sc_hd__a21oi_1 _11568_ (.A1(_06116_),
    .A2(\reg_next_pc[6] ),
    .B1(_06135_),
    .Y(_06136_));
 sky130_fd_sc_hd__and3_1 _11569_ (.A(\reg_pc[6] ),
    .B(\reg_pc[5] ),
    .C(_06121_),
    .X(_06137_));
 sky130_fd_sc_hd__a21oi_1 _11570_ (.A1(\reg_pc[5] ),
    .A2(_06121_),
    .B1(\reg_pc[6] ),
    .Y(_06138_));
 sky130_fd_sc_hd__o21a_1 _11571_ (.A1(_06137_),
    .A2(_06138_),
    .B1(_06075_),
    .X(_06139_));
 sky130_fd_sc_hd__nor2_2 _11572_ (.A(_06136_),
    .B(_06139_),
    .Y(_06140_));
 sky130_fd_sc_hd__buf_2 _11573_ (.A(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__mux2_1 _11574_ (.A0(_06141_),
    .A1(\cpuregs.regs[10][6] ),
    .S(_06086_),
    .X(_06142_));
 sky130_fd_sc_hd__clkbuf_1 _11575_ (.A(_06142_),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _11576_ (.A0(\reg_out[7] ),
    .A1(\alu_out_q[7] ),
    .S(_06067_),
    .X(_06143_));
 sky130_fd_sc_hd__a221o_1 _11577_ (.A1(_06072_),
    .A2(_03349_),
    .B1(_06098_),
    .B2(_06143_),
    .C1(_06118_),
    .X(_06144_));
 sky130_fd_sc_hd__a21oi_1 _11578_ (.A1(_06116_),
    .A2(\reg_next_pc[7] ),
    .B1(_06144_),
    .Y(_06145_));
 sky130_fd_sc_hd__and2_1 _11579_ (.A(\reg_pc[7] ),
    .B(_06137_),
    .X(_06146_));
 sky130_fd_sc_hd__nor2_1 _11580_ (.A(\reg_pc[7] ),
    .B(_06137_),
    .Y(_06147_));
 sky130_fd_sc_hd__o21a_1 _11581_ (.A1(_06146_),
    .A2(_06147_),
    .B1(_06075_),
    .X(_06148_));
 sky130_fd_sc_hd__nor2_2 _11582_ (.A(_06145_),
    .B(_06148_),
    .Y(_06149_));
 sky130_fd_sc_hd__buf_2 _11583_ (.A(_06149_),
    .X(_06150_));
 sky130_fd_sc_hd__mux2_1 _11584_ (.A0(_06150_),
    .A1(\cpuregs.regs[10][7] ),
    .S(_06086_),
    .X(_06151_));
 sky130_fd_sc_hd__clkbuf_1 _11585_ (.A(_06151_),
    .X(_00102_));
 sky130_fd_sc_hd__xnor2_1 _11586_ (.A(\reg_pc[8] ),
    .B(_06146_),
    .Y(_06152_));
 sky130_fd_sc_hd__mux2_1 _11587_ (.A0(\reg_out[8] ),
    .A1(\alu_out_q[8] ),
    .S(_06067_),
    .X(_06153_));
 sky130_fd_sc_hd__a221o_1 _11588_ (.A1(\irq_state[1] ),
    .A2(_03359_),
    .B1(_06065_),
    .B2(_06153_),
    .C1(_06074_),
    .X(_06154_));
 sky130_fd_sc_hd__a21oi_2 _11589_ (.A1(_06071_),
    .A2(\reg_next_pc[8] ),
    .B1(_06154_),
    .Y(_06155_));
 sky130_fd_sc_hd__a21oi_4 _11590_ (.A1(_06075_),
    .A2(_06152_),
    .B1(_06155_),
    .Y(_06156_));
 sky130_fd_sc_hd__buf_2 _11591_ (.A(_06156_),
    .X(_06157_));
 sky130_fd_sc_hd__mux2_1 _11592_ (.A0(_06157_),
    .A1(\cpuregs.regs[10][8] ),
    .S(_06086_),
    .X(_06158_));
 sky130_fd_sc_hd__clkbuf_1 _11593_ (.A(_06158_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _11594_ (.A0(\reg_out[9] ),
    .A1(\alu_out_q[9] ),
    .S(_06067_),
    .X(_06159_));
 sky130_fd_sc_hd__a221o_1 _11595_ (.A1(\irq_state[1] ),
    .A2(_03323_),
    .B1(_06098_),
    .B2(_06159_),
    .C1(_06118_),
    .X(_06160_));
 sky130_fd_sc_hd__a21oi_1 _11596_ (.A1(_06116_),
    .A2(\reg_next_pc[9] ),
    .B1(_06160_),
    .Y(_06161_));
 sky130_fd_sc_hd__and3_1 _11597_ (.A(\reg_pc[9] ),
    .B(\reg_pc[8] ),
    .C(_06146_),
    .X(_06162_));
 sky130_fd_sc_hd__a21oi_1 _11598_ (.A1(\reg_pc[8] ),
    .A2(_06146_),
    .B1(\reg_pc[9] ),
    .Y(_06163_));
 sky130_fd_sc_hd__o21a_1 _11599_ (.A1(_06162_),
    .A2(_06163_),
    .B1(_06075_),
    .X(_06164_));
 sky130_fd_sc_hd__nor2_2 _11600_ (.A(_06161_),
    .B(_06164_),
    .Y(_06165_));
 sky130_fd_sc_hd__buf_2 _11601_ (.A(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__mux2_1 _11602_ (.A0(_06166_),
    .A1(\cpuregs.regs[10][9] ),
    .S(_06086_),
    .X(_06167_));
 sky130_fd_sc_hd__clkbuf_1 _11603_ (.A(_06167_),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _11604_ (.A0(\reg_out[10] ),
    .A1(\alu_out_q[10] ),
    .S(_06067_),
    .X(_06168_));
 sky130_fd_sc_hd__a221o_1 _11605_ (.A1(\irq_state[1] ),
    .A2(_03333_),
    .B1(_06098_),
    .B2(_06168_),
    .C1(_06074_),
    .X(_06169_));
 sky130_fd_sc_hd__a21oi_1 _11606_ (.A1(_06116_),
    .A2(\reg_next_pc[10] ),
    .B1(_06169_),
    .Y(_06170_));
 sky130_fd_sc_hd__and2_1 _11607_ (.A(\reg_pc[10] ),
    .B(_06162_),
    .X(_06171_));
 sky130_fd_sc_hd__nor2_1 _11608_ (.A(\reg_pc[10] ),
    .B(_06162_),
    .Y(_06172_));
 sky130_fd_sc_hd__o21a_1 _11609_ (.A1(_06171_),
    .A2(_06172_),
    .B1(_06075_),
    .X(_06173_));
 sky130_fd_sc_hd__nor2_4 _11610_ (.A(_06170_),
    .B(_06173_),
    .Y(_06174_));
 sky130_fd_sc_hd__buf_2 _11611_ (.A(_06174_),
    .X(_06175_));
 sky130_fd_sc_hd__clkbuf_8 _11612_ (.A(_06085_),
    .X(_06176_));
 sky130_fd_sc_hd__mux2_1 _11613_ (.A0(_06175_),
    .A1(\cpuregs.regs[10][10] ),
    .S(_06176_),
    .X(_06177_));
 sky130_fd_sc_hd__clkbuf_1 _11614_ (.A(_06177_),
    .X(_00105_));
 sky130_fd_sc_hd__nand2_1 _11615_ (.A(\reg_pc[11] ),
    .B(_06171_),
    .Y(_06178_));
 sky130_fd_sc_hd__or2_1 _11616_ (.A(\reg_pc[11] ),
    .B(_06171_),
    .X(_06179_));
 sky130_fd_sc_hd__mux2_1 _11617_ (.A0(\reg_out[11] ),
    .A1(\alu_out_q[11] ),
    .S(_06067_),
    .X(_06180_));
 sky130_fd_sc_hd__a22o_1 _11618_ (.A1(\irq_state[1] ),
    .A2(_03335_),
    .B1(_06065_),
    .B2(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__a21o_1 _11619_ (.A1(_06071_),
    .A2(\reg_next_pc[11] ),
    .B1(_06181_),
    .X(_06182_));
 sky130_fd_sc_hd__a31o_2 _11620_ (.A1(_06075_),
    .A2(_06178_),
    .A3(_06179_),
    .B1(_06182_),
    .X(_06183_));
 sky130_fd_sc_hd__buf_2 _11621_ (.A(_06183_),
    .X(_06184_));
 sky130_fd_sc_hd__mux2_1 _11622_ (.A0(_06184_),
    .A1(\cpuregs.regs[10][11] ),
    .S(_06176_),
    .X(_06185_));
 sky130_fd_sc_hd__clkbuf_1 _11623_ (.A(_06185_),
    .X(_00106_));
 sky130_fd_sc_hd__buf_4 _11624_ (.A(_06071_),
    .X(_06186_));
 sky130_fd_sc_hd__and3_1 _11625_ (.A(\reg_pc[12] ),
    .B(\reg_pc[11] ),
    .C(_06171_),
    .X(_06187_));
 sky130_fd_sc_hd__a31o_1 _11626_ (.A1(\reg_pc[11] ),
    .A2(\reg_pc[10] ),
    .A3(_06162_),
    .B1(\reg_pc[12] ),
    .X(_06188_));
 sky130_fd_sc_hd__and3b_1 _11627_ (.A_N(_06187_),
    .B(_06118_),
    .C(_06188_),
    .X(_06189_));
 sky130_fd_sc_hd__mux2_1 _11628_ (.A0(\reg_out[12] ),
    .A1(\alu_out_q[12] ),
    .S(_06067_),
    .X(_06190_));
 sky130_fd_sc_hd__a22o_1 _11629_ (.A1(_03409_),
    .A2(_03357_),
    .B1(_06066_),
    .B2(_06190_),
    .X(_06191_));
 sky130_fd_sc_hd__a211o_2 _11630_ (.A1(_06186_),
    .A2(\reg_next_pc[12] ),
    .B1(_06189_),
    .C1(_06191_),
    .X(_06192_));
 sky130_fd_sc_hd__buf_2 _11631_ (.A(_06192_),
    .X(_06193_));
 sky130_fd_sc_hd__mux2_1 _11632_ (.A0(_06193_),
    .A1(\cpuregs.regs[10][12] ),
    .S(_06176_),
    .X(_06194_));
 sky130_fd_sc_hd__clkbuf_1 _11633_ (.A(_06194_),
    .X(_00107_));
 sky130_fd_sc_hd__and2_1 _11634_ (.A(\reg_pc[13] ),
    .B(_06187_),
    .X(_06195_));
 sky130_fd_sc_hd__o21ai_1 _11635_ (.A1(\reg_pc[13] ),
    .A2(_06187_),
    .B1(_06075_),
    .Y(_06196_));
 sky130_fd_sc_hd__nor2_1 _11636_ (.A(_06195_),
    .B(_06196_),
    .Y(_06197_));
 sky130_fd_sc_hd__mux2_1 _11637_ (.A0(\reg_out[13] ),
    .A1(\alu_out_q[13] ),
    .S(_06068_),
    .X(_06198_));
 sky130_fd_sc_hd__a22o_1 _11638_ (.A1(_03409_),
    .A2(_03352_),
    .B1(_06066_),
    .B2(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__a211o_4 _11639_ (.A1(_06186_),
    .A2(\reg_next_pc[13] ),
    .B1(_06197_),
    .C1(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__buf_2 _11640_ (.A(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__mux2_1 _11641_ (.A0(_06201_),
    .A1(\cpuregs.regs[10][13] ),
    .S(_06176_),
    .X(_06202_));
 sky130_fd_sc_hd__clkbuf_1 _11642_ (.A(_06202_),
    .X(_00108_));
 sky130_fd_sc_hd__a21oi_1 _11643_ (.A1(\reg_pc[14] ),
    .A2(_06195_),
    .B1(_06093_),
    .Y(_06203_));
 sky130_fd_sc_hd__o21a_1 _11644_ (.A1(\reg_pc[14] ),
    .A2(_06195_),
    .B1(_06203_),
    .X(_06204_));
 sky130_fd_sc_hd__mux2_1 _11645_ (.A0(\reg_out[14] ),
    .A1(\alu_out_q[14] ),
    .S(_06068_),
    .X(_06205_));
 sky130_fd_sc_hd__a22o_1 _11646_ (.A1(_03409_),
    .A2(_03353_),
    .B1(_06066_),
    .B2(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__a211o_2 _11647_ (.A1(_06186_),
    .A2(\reg_next_pc[14] ),
    .B1(_06204_),
    .C1(_06206_),
    .X(_06207_));
 sky130_fd_sc_hd__buf_2 _11648_ (.A(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__mux2_1 _11649_ (.A0(_06208_),
    .A1(\cpuregs.regs[10][14] ),
    .S(_06176_),
    .X(_06209_));
 sky130_fd_sc_hd__clkbuf_1 _11650_ (.A(_06209_),
    .X(_00109_));
 sky130_fd_sc_hd__and3_1 _11651_ (.A(\reg_pc[15] ),
    .B(\reg_pc[14] ),
    .C(_06195_),
    .X(_06210_));
 sky130_fd_sc_hd__a31o_1 _11652_ (.A1(\reg_pc[14] ),
    .A2(\reg_pc[13] ),
    .A3(_06187_),
    .B1(\reg_pc[15] ),
    .X(_06211_));
 sky130_fd_sc_hd__and3b_1 _11653_ (.A_N(_06210_),
    .B(_06118_),
    .C(_06211_),
    .X(_06212_));
 sky130_fd_sc_hd__mux2_1 _11654_ (.A0(\reg_out[15] ),
    .A1(\alu_out_q[15] ),
    .S(_06067_),
    .X(_06213_));
 sky130_fd_sc_hd__a22o_1 _11655_ (.A1(_03409_),
    .A2(_03356_),
    .B1(_06066_),
    .B2(_06213_),
    .X(_06214_));
 sky130_fd_sc_hd__a211o_2 _11656_ (.A1(_06186_),
    .A2(\reg_next_pc[15] ),
    .B1(_06212_),
    .C1(_06214_),
    .X(_06215_));
 sky130_fd_sc_hd__buf_2 _11657_ (.A(_06215_),
    .X(_06216_));
 sky130_fd_sc_hd__mux2_1 _11658_ (.A0(_06216_),
    .A1(\cpuregs.regs[10][15] ),
    .S(_06176_),
    .X(_06217_));
 sky130_fd_sc_hd__clkbuf_1 _11659_ (.A(_06217_),
    .X(_00110_));
 sky130_fd_sc_hd__and2_1 _11660_ (.A(\reg_pc[16] ),
    .B(_06210_),
    .X(_06218_));
 sky130_fd_sc_hd__o21ai_1 _11661_ (.A1(\reg_pc[16] ),
    .A2(_06210_),
    .B1(_06101_),
    .Y(_06219_));
 sky130_fd_sc_hd__nor2_1 _11662_ (.A(_06218_),
    .B(_06219_),
    .Y(_06220_));
 sky130_fd_sc_hd__mux2_1 _11663_ (.A0(\reg_out[16] ),
    .A1(\alu_out_q[16] ),
    .S(_06067_),
    .X(_06221_));
 sky130_fd_sc_hd__a22o_1 _11664_ (.A1(_03409_),
    .A2(_03330_),
    .B1(_06066_),
    .B2(_06221_),
    .X(_06222_));
 sky130_fd_sc_hd__a211o_4 _11665_ (.A1(_06186_),
    .A2(\reg_next_pc[16] ),
    .B1(_06220_),
    .C1(_06222_),
    .X(_06223_));
 sky130_fd_sc_hd__buf_2 _11666_ (.A(_06223_),
    .X(_06224_));
 sky130_fd_sc_hd__mux2_1 _11667_ (.A0(_06224_),
    .A1(\cpuregs.regs[10][16] ),
    .S(_06176_),
    .X(_06225_));
 sky130_fd_sc_hd__clkbuf_1 _11668_ (.A(_06225_),
    .X(_00111_));
 sky130_fd_sc_hd__clkbuf_4 _11669_ (.A(_06071_),
    .X(_06226_));
 sky130_fd_sc_hd__a21oi_1 _11670_ (.A1(\reg_pc[17] ),
    .A2(_06218_),
    .B1(_06093_),
    .Y(_06227_));
 sky130_fd_sc_hd__o21a_1 _11671_ (.A1(\reg_pc[17] ),
    .A2(_06218_),
    .B1(_06227_),
    .X(_06228_));
 sky130_fd_sc_hd__mux2_1 _11672_ (.A0(\reg_out[17] ),
    .A1(\alu_out_q[17] ),
    .S(_06068_),
    .X(_06229_));
 sky130_fd_sc_hd__a22o_1 _11673_ (.A1(_03409_),
    .A2(_03348_),
    .B1(_06066_),
    .B2(_06229_),
    .X(_06230_));
 sky130_fd_sc_hd__a211o_4 _11674_ (.A1(_06226_),
    .A2(\reg_next_pc[17] ),
    .B1(_06228_),
    .C1(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__buf_2 _11675_ (.A(_06231_),
    .X(_06232_));
 sky130_fd_sc_hd__mux2_1 _11676_ (.A0(_06232_),
    .A1(\cpuregs.regs[10][17] ),
    .S(_06176_),
    .X(_06233_));
 sky130_fd_sc_hd__clkbuf_1 _11677_ (.A(_06233_),
    .X(_00112_));
 sky130_fd_sc_hd__and3_1 _11678_ (.A(\reg_pc[18] ),
    .B(\reg_pc[17] ),
    .C(_06218_),
    .X(_06234_));
 sky130_fd_sc_hd__a31o_1 _11679_ (.A1(\reg_pc[17] ),
    .A2(\reg_pc[16] ),
    .A3(_06210_),
    .B1(\reg_pc[18] ),
    .X(_06235_));
 sky130_fd_sc_hd__and3b_1 _11680_ (.A_N(_06234_),
    .B(_06118_),
    .C(_06235_),
    .X(_06236_));
 sky130_fd_sc_hd__mux2_1 _11681_ (.A0(\reg_out[18] ),
    .A1(\alu_out_q[18] ),
    .S(_06068_),
    .X(_06237_));
 sky130_fd_sc_hd__a22o_1 _11682_ (.A1(_03409_),
    .A2(_03336_),
    .B1(_06066_),
    .B2(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__a211o_2 _11683_ (.A1(_06226_),
    .A2(\reg_next_pc[18] ),
    .B1(_06236_),
    .C1(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__buf_2 _11684_ (.A(_06239_),
    .X(_06240_));
 sky130_fd_sc_hd__mux2_1 _11685_ (.A0(_06240_),
    .A1(\cpuregs.regs[10][18] ),
    .S(_06176_),
    .X(_06241_));
 sky130_fd_sc_hd__clkbuf_1 _11686_ (.A(_06241_),
    .X(_00113_));
 sky130_fd_sc_hd__and2_1 _11687_ (.A(\reg_pc[19] ),
    .B(_06234_),
    .X(_06242_));
 sky130_fd_sc_hd__o21ai_1 _11688_ (.A1(\reg_pc[19] ),
    .A2(_06234_),
    .B1(_06101_),
    .Y(_06243_));
 sky130_fd_sc_hd__nor2_1 _11689_ (.A(_06242_),
    .B(_06243_),
    .Y(_06244_));
 sky130_fd_sc_hd__mux2_1 _11690_ (.A0(\reg_out[19] ),
    .A1(\alu_out_q[19] ),
    .S(_06068_),
    .X(_06245_));
 sky130_fd_sc_hd__a22o_1 _11691_ (.A1(_03409_),
    .A2(_03358_),
    .B1(_06066_),
    .B2(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__a211o_2 _11692_ (.A1(_06226_),
    .A2(\reg_next_pc[19] ),
    .B1(_06244_),
    .C1(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__buf_2 _11693_ (.A(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__mux2_1 _11694_ (.A0(_06248_),
    .A1(\cpuregs.regs[10][19] ),
    .S(_06176_),
    .X(_06249_));
 sky130_fd_sc_hd__clkbuf_1 _11695_ (.A(_06249_),
    .X(_00114_));
 sky130_fd_sc_hd__a21oi_1 _11696_ (.A1(\reg_pc[20] ),
    .A2(_06242_),
    .B1(_06093_),
    .Y(_06250_));
 sky130_fd_sc_hd__o21a_1 _11697_ (.A1(\reg_pc[20] ),
    .A2(_06242_),
    .B1(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__clkbuf_4 _11698_ (.A(\irq_state[1] ),
    .X(_06252_));
 sky130_fd_sc_hd__buf_2 _11699_ (.A(_06065_),
    .X(_06253_));
 sky130_fd_sc_hd__mux2_1 _11700_ (.A0(\reg_out[20] ),
    .A1(\alu_out_q[20] ),
    .S(_06068_),
    .X(_06254_));
 sky130_fd_sc_hd__a22o_1 _11701_ (.A1(_06252_),
    .A2(_03332_),
    .B1(_06253_),
    .B2(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__a211o_2 _11702_ (.A1(_06226_),
    .A2(\reg_next_pc[20] ),
    .B1(_06251_),
    .C1(_06255_),
    .X(_06256_));
 sky130_fd_sc_hd__buf_2 _11703_ (.A(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__clkbuf_8 _11704_ (.A(_06085_),
    .X(_06258_));
 sky130_fd_sc_hd__mux2_1 _11705_ (.A0(_06257_),
    .A1(\cpuregs.regs[10][20] ),
    .S(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__clkbuf_1 _11706_ (.A(_06259_),
    .X(_00115_));
 sky130_fd_sc_hd__and3_1 _11707_ (.A(\reg_pc[21] ),
    .B(\reg_pc[20] ),
    .C(_06242_),
    .X(_06260_));
 sky130_fd_sc_hd__a31o_1 _11708_ (.A1(\reg_pc[20] ),
    .A2(\reg_pc[19] ),
    .A3(_06234_),
    .B1(\reg_pc[21] ),
    .X(_06261_));
 sky130_fd_sc_hd__and3b_1 _11709_ (.A_N(_06260_),
    .B(_06118_),
    .C(_06261_),
    .X(_06262_));
 sky130_fd_sc_hd__mux2_1 _11710_ (.A0(\reg_out[21] ),
    .A1(\alu_out_q[21] ),
    .S(_06069_),
    .X(_06263_));
 sky130_fd_sc_hd__a22o_1 _11711_ (.A1(_06252_),
    .A2(_03346_),
    .B1(_06253_),
    .B2(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__a211o_2 _11712_ (.A1(_06226_),
    .A2(\reg_next_pc[21] ),
    .B1(_06262_),
    .C1(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__buf_2 _11713_ (.A(_06265_),
    .X(_06266_));
 sky130_fd_sc_hd__mux2_1 _11714_ (.A0(_06266_),
    .A1(\cpuregs.regs[10][21] ),
    .S(_06258_),
    .X(_06267_));
 sky130_fd_sc_hd__clkbuf_1 _11715_ (.A(_06267_),
    .X(_00116_));
 sky130_fd_sc_hd__and2_1 _11716_ (.A(\reg_pc[22] ),
    .B(_06260_),
    .X(_06268_));
 sky130_fd_sc_hd__o21ai_1 _11717_ (.A1(\reg_pc[22] ),
    .A2(_06260_),
    .B1(_06101_),
    .Y(_06269_));
 sky130_fd_sc_hd__nor2_1 _11718_ (.A(_06268_),
    .B(_06269_),
    .Y(_06270_));
 sky130_fd_sc_hd__mux2_1 _11719_ (.A0(\reg_out[22] ),
    .A1(\alu_out_q[22] ),
    .S(_06068_),
    .X(_06271_));
 sky130_fd_sc_hd__a22o_1 _11720_ (.A1(_06252_),
    .A2(_03320_),
    .B1(_06253_),
    .B2(_06271_),
    .X(_06272_));
 sky130_fd_sc_hd__a211o_2 _11721_ (.A1(_06226_),
    .A2(\reg_next_pc[22] ),
    .B1(_06270_),
    .C1(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__buf_2 _11722_ (.A(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__mux2_1 _11723_ (.A0(_06274_),
    .A1(\cpuregs.regs[10][22] ),
    .S(_06258_),
    .X(_06275_));
 sky130_fd_sc_hd__clkbuf_1 _11724_ (.A(_06275_),
    .X(_00117_));
 sky130_fd_sc_hd__a21oi_1 _11725_ (.A1(\reg_pc[23] ),
    .A2(_06268_),
    .B1(_06093_),
    .Y(_06276_));
 sky130_fd_sc_hd__o21a_1 _11726_ (.A1(\reg_pc[23] ),
    .A2(_06268_),
    .B1(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__mux2_1 _11727_ (.A0(\reg_out[23] ),
    .A1(\alu_out_q[23] ),
    .S(_06068_),
    .X(_06278_));
 sky130_fd_sc_hd__a22o_1 _11728_ (.A1(_06252_),
    .A2(_03343_),
    .B1(_06253_),
    .B2(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__a211o_2 _11729_ (.A1(_06226_),
    .A2(\reg_next_pc[23] ),
    .B1(_06277_),
    .C1(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__clkbuf_2 _11730_ (.A(_06280_),
    .X(_06281_));
 sky130_fd_sc_hd__mux2_1 _11731_ (.A0(_06281_),
    .A1(\cpuregs.regs[10][23] ),
    .S(_06258_),
    .X(_06282_));
 sky130_fd_sc_hd__clkbuf_1 _11732_ (.A(_06282_),
    .X(_00118_));
 sky130_fd_sc_hd__and3_1 _11733_ (.A(\reg_pc[24] ),
    .B(\reg_pc[23] ),
    .C(_06268_),
    .X(_06283_));
 sky130_fd_sc_hd__a31o_1 _11734_ (.A1(\reg_pc[23] ),
    .A2(\reg_pc[22] ),
    .A3(_06260_),
    .B1(\reg_pc[24] ),
    .X(_06284_));
 sky130_fd_sc_hd__and3b_1 _11735_ (.A_N(_06283_),
    .B(_06118_),
    .C(_06284_),
    .X(_06285_));
 sky130_fd_sc_hd__mux2_2 _11736_ (.A0(\reg_out[24] ),
    .A1(\alu_out_q[24] ),
    .S(_06068_),
    .X(_06286_));
 sky130_fd_sc_hd__a22o_1 _11737_ (.A1(_06252_),
    .A2(_03342_),
    .B1(_06253_),
    .B2(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__a211o_2 _11738_ (.A1(_06226_),
    .A2(\reg_next_pc[24] ),
    .B1(_06285_),
    .C1(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__buf_2 _11739_ (.A(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__mux2_1 _11740_ (.A0(_06289_),
    .A1(\cpuregs.regs[10][24] ),
    .S(_06258_),
    .X(_06290_));
 sky130_fd_sc_hd__clkbuf_1 _11741_ (.A(_06290_),
    .X(_00119_));
 sky130_fd_sc_hd__and2_1 _11742_ (.A(\reg_pc[25] ),
    .B(_06283_),
    .X(_06291_));
 sky130_fd_sc_hd__o21ai_1 _11743_ (.A1(\reg_pc[25] ),
    .A2(_06283_),
    .B1(_06101_),
    .Y(_06292_));
 sky130_fd_sc_hd__nor2_1 _11744_ (.A(_06291_),
    .B(_06292_),
    .Y(_06293_));
 sky130_fd_sc_hd__mux2_1 _11745_ (.A0(\reg_out[25] ),
    .A1(\alu_out_q[25] ),
    .S(_06069_),
    .X(_06294_));
 sky130_fd_sc_hd__a22o_1 _11746_ (.A1(_06252_),
    .A2(_03347_),
    .B1(_06253_),
    .B2(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__a211o_2 _11747_ (.A1(_06226_),
    .A2(\reg_next_pc[25] ),
    .B1(_06293_),
    .C1(_06295_),
    .X(_06296_));
 sky130_fd_sc_hd__buf_2 _11748_ (.A(_06296_),
    .X(_06297_));
 sky130_fd_sc_hd__mux2_1 _11749_ (.A0(_06297_),
    .A1(\cpuregs.regs[10][25] ),
    .S(_06258_),
    .X(_06298_));
 sky130_fd_sc_hd__clkbuf_1 _11750_ (.A(_06298_),
    .X(_00120_));
 sky130_fd_sc_hd__a21oi_1 _11751_ (.A1(\reg_pc[26] ),
    .A2(_06291_),
    .B1(_06093_),
    .Y(_06299_));
 sky130_fd_sc_hd__o21a_1 _11752_ (.A1(\reg_pc[26] ),
    .A2(_06291_),
    .B1(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__mux2_1 _11753_ (.A0(\reg_out[26] ),
    .A1(\alu_out_q[26] ),
    .S(_06069_),
    .X(_06301_));
 sky130_fd_sc_hd__a22o_1 _11754_ (.A1(_06252_),
    .A2(_03325_),
    .B1(_06253_),
    .B2(_06301_),
    .X(_06302_));
 sky130_fd_sc_hd__a211o_2 _11755_ (.A1(_06226_),
    .A2(\reg_next_pc[26] ),
    .B1(_06300_),
    .C1(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__buf_2 _11756_ (.A(_06303_),
    .X(_06304_));
 sky130_fd_sc_hd__mux2_1 _11757_ (.A0(_06304_),
    .A1(\cpuregs.regs[10][26] ),
    .S(_06258_),
    .X(_06305_));
 sky130_fd_sc_hd__clkbuf_1 _11758_ (.A(_06305_),
    .X(_00121_));
 sky130_fd_sc_hd__and3_1 _11759_ (.A(\reg_pc[27] ),
    .B(\reg_pc[26] ),
    .C(_06291_),
    .X(_06306_));
 sky130_fd_sc_hd__a31o_1 _11760_ (.A1(\reg_pc[26] ),
    .A2(\reg_pc[25] ),
    .A3(_06283_),
    .B1(\reg_pc[27] ),
    .X(_06307_));
 sky130_fd_sc_hd__and3b_1 _11761_ (.A_N(_06306_),
    .B(_06118_),
    .C(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__mux2_1 _11762_ (.A0(\reg_out[27] ),
    .A1(\alu_out_q[27] ),
    .S(_06069_),
    .X(_06309_));
 sky130_fd_sc_hd__a22o_1 _11763_ (.A1(_06252_),
    .A2(_03341_),
    .B1(_06253_),
    .B2(_06309_),
    .X(_06310_));
 sky130_fd_sc_hd__a211o_1 _11764_ (.A1(_06116_),
    .A2(\reg_next_pc[27] ),
    .B1(_06308_),
    .C1(_06310_),
    .X(_06311_));
 sky130_fd_sc_hd__buf_2 _11765_ (.A(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__mux2_1 _11766_ (.A0(_06312_),
    .A1(\cpuregs.regs[10][27] ),
    .S(_06258_),
    .X(_06313_));
 sky130_fd_sc_hd__clkbuf_1 _11767_ (.A(_06313_),
    .X(_00122_));
 sky130_fd_sc_hd__and2_1 _11768_ (.A(\reg_pc[28] ),
    .B(_06306_),
    .X(_06314_));
 sky130_fd_sc_hd__o21ai_1 _11769_ (.A1(\reg_pc[28] ),
    .A2(_06306_),
    .B1(_06101_),
    .Y(_06315_));
 sky130_fd_sc_hd__nor2_1 _11770_ (.A(_06314_),
    .B(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__mux2_1 _11771_ (.A0(\reg_out[28] ),
    .A1(\alu_out_q[28] ),
    .S(_06069_),
    .X(_06317_));
 sky130_fd_sc_hd__a22o_1 _11772_ (.A1(_06252_),
    .A2(_03354_),
    .B1(_06253_),
    .B2(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__a211o_2 _11773_ (.A1(_06116_),
    .A2(\reg_next_pc[28] ),
    .B1(_06316_),
    .C1(_06318_),
    .X(_06319_));
 sky130_fd_sc_hd__buf_2 _11774_ (.A(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__mux2_1 _11775_ (.A0(_06320_),
    .A1(\cpuregs.regs[10][28] ),
    .S(_06258_),
    .X(_06321_));
 sky130_fd_sc_hd__clkbuf_1 _11776_ (.A(_06321_),
    .X(_00123_));
 sky130_fd_sc_hd__and3_1 _11777_ (.A(\reg_pc[29] ),
    .B(\reg_pc[28] ),
    .C(_06306_),
    .X(_06322_));
 sky130_fd_sc_hd__o21ai_1 _11778_ (.A1(\reg_pc[29] ),
    .A2(_06314_),
    .B1(_06101_),
    .Y(_06323_));
 sky130_fd_sc_hd__nor2_1 _11779_ (.A(_06322_),
    .B(_06323_),
    .Y(_06324_));
 sky130_fd_sc_hd__mux2_1 _11780_ (.A0(\reg_out[29] ),
    .A1(\alu_out_q[29] ),
    .S(_06069_),
    .X(_06325_));
 sky130_fd_sc_hd__a22o_1 _11781_ (.A1(_06252_),
    .A2(_03337_),
    .B1(_06253_),
    .B2(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__a211o_2 _11782_ (.A1(_06116_),
    .A2(\reg_next_pc[29] ),
    .B1(_06324_),
    .C1(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__buf_2 _11783_ (.A(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__mux2_1 _11784_ (.A0(_06328_),
    .A1(\cpuregs.regs[10][29] ),
    .S(_06258_),
    .X(_06329_));
 sky130_fd_sc_hd__clkbuf_1 _11785_ (.A(_06329_),
    .X(_00124_));
 sky130_fd_sc_hd__and2_1 _11786_ (.A(\reg_pc[30] ),
    .B(_06322_),
    .X(_06330_));
 sky130_fd_sc_hd__o21ai_1 _11787_ (.A1(\reg_pc[30] ),
    .A2(_06322_),
    .B1(_06101_),
    .Y(_06331_));
 sky130_fd_sc_hd__nor2_1 _11788_ (.A(_06330_),
    .B(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__mux2_1 _11789_ (.A0(\reg_out[30] ),
    .A1(\alu_out_q[30] ),
    .S(_06069_),
    .X(_06333_));
 sky130_fd_sc_hd__a22o_1 _11790_ (.A1(_06072_),
    .A2(_03328_),
    .B1(_06098_),
    .B2(_06333_),
    .X(_06334_));
 sky130_fd_sc_hd__a211o_4 _11791_ (.A1(_06116_),
    .A2(\reg_next_pc[30] ),
    .B1(_06332_),
    .C1(_06334_),
    .X(_06335_));
 sky130_fd_sc_hd__buf_2 _11792_ (.A(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__mux2_1 _11793_ (.A0(_06336_),
    .A1(\cpuregs.regs[10][30] ),
    .S(_06085_),
    .X(_06337_));
 sky130_fd_sc_hd__clkbuf_1 _11794_ (.A(_06337_),
    .X(_00125_));
 sky130_fd_sc_hd__o21ai_1 _11795_ (.A1(\reg_pc[31] ),
    .A2(_06330_),
    .B1(_06101_),
    .Y(_06338_));
 sky130_fd_sc_hd__a21oi_1 _11796_ (.A1(\reg_pc[31] ),
    .A2(_06330_),
    .B1(_06338_),
    .Y(_06339_));
 sky130_fd_sc_hd__mux2_1 _11797_ (.A0(\reg_out[31] ),
    .A1(\alu_out_q[31] ),
    .S(_06069_),
    .X(_06340_));
 sky130_fd_sc_hd__a22o_1 _11798_ (.A1(_06072_),
    .A2(_03331_),
    .B1(_06098_),
    .B2(_06340_),
    .X(_06341_));
 sky130_fd_sc_hd__a211o_2 _11799_ (.A1(_06116_),
    .A2(\reg_next_pc[31] ),
    .B1(_06339_),
    .C1(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__buf_2 _11800_ (.A(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__mux2_1 _11801_ (.A0(_06343_),
    .A1(\cpuregs.regs[10][31] ),
    .S(_06085_),
    .X(_06344_));
 sky130_fd_sc_hd__clkbuf_1 _11802_ (.A(_06344_),
    .X(_00126_));
 sky130_fd_sc_hd__and2_1 _11803_ (.A(\cpuregs.waddr[1] ),
    .B(\cpuregs.waddr[0] ),
    .X(_06345_));
 sky130_fd_sc_hd__buf_4 _11804_ (.A(_06345_),
    .X(_06346_));
 sky130_fd_sc_hd__nand2_2 _11805_ (.A(_06084_),
    .B(_06346_),
    .Y(_06347_));
 sky130_fd_sc_hd__buf_6 _11806_ (.A(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__mux2_1 _11807_ (.A0(_06078_),
    .A1(\cpuregs.regs[11][0] ),
    .S(_06348_),
    .X(_06349_));
 sky130_fd_sc_hd__clkbuf_1 _11808_ (.A(_06349_),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _11809_ (.A0(_06096_),
    .A1(\cpuregs.regs[11][1] ),
    .S(_06348_),
    .X(_06350_));
 sky130_fd_sc_hd__clkbuf_1 _11810_ (.A(_06350_),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _11811_ (.A0(_06105_),
    .A1(\cpuregs.regs[11][2] ),
    .S(_06348_),
    .X(_06351_));
 sky130_fd_sc_hd__clkbuf_1 _11812_ (.A(_06351_),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _11813_ (.A0(_06114_),
    .A1(\cpuregs.regs[11][3] ),
    .S(_06348_),
    .X(_06352_));
 sky130_fd_sc_hd__clkbuf_1 _11814_ (.A(_06352_),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _11815_ (.A0(_06125_),
    .A1(\cpuregs.regs[11][4] ),
    .S(_06348_),
    .X(_06353_));
 sky130_fd_sc_hd__clkbuf_1 _11816_ (.A(_06353_),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _11817_ (.A0(_06132_),
    .A1(\cpuregs.regs[11][5] ),
    .S(_06348_),
    .X(_06354_));
 sky130_fd_sc_hd__clkbuf_1 _11818_ (.A(_06354_),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _11819_ (.A0(_06141_),
    .A1(\cpuregs.regs[11][6] ),
    .S(_06348_),
    .X(_06355_));
 sky130_fd_sc_hd__clkbuf_1 _11820_ (.A(_06355_),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _11821_ (.A0(_06150_),
    .A1(\cpuregs.regs[11][7] ),
    .S(_06348_),
    .X(_06356_));
 sky130_fd_sc_hd__clkbuf_1 _11822_ (.A(_06356_),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _11823_ (.A0(_06157_),
    .A1(\cpuregs.regs[11][8] ),
    .S(_06348_),
    .X(_06357_));
 sky130_fd_sc_hd__clkbuf_1 _11824_ (.A(_06357_),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _11825_ (.A0(_06166_),
    .A1(\cpuregs.regs[11][9] ),
    .S(_06348_),
    .X(_06358_));
 sky130_fd_sc_hd__clkbuf_1 _11826_ (.A(_06358_),
    .X(_00136_));
 sky130_fd_sc_hd__clkbuf_8 _11827_ (.A(_06347_),
    .X(_06359_));
 sky130_fd_sc_hd__mux2_1 _11828_ (.A0(_06175_),
    .A1(\cpuregs.regs[11][10] ),
    .S(_06359_),
    .X(_06360_));
 sky130_fd_sc_hd__clkbuf_1 _11829_ (.A(_06360_),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _11830_ (.A0(_06184_),
    .A1(\cpuregs.regs[11][11] ),
    .S(_06359_),
    .X(_06361_));
 sky130_fd_sc_hd__clkbuf_1 _11831_ (.A(_06361_),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _11832_ (.A0(_06193_),
    .A1(\cpuregs.regs[11][12] ),
    .S(_06359_),
    .X(_06362_));
 sky130_fd_sc_hd__clkbuf_1 _11833_ (.A(_06362_),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _11834_ (.A0(_06201_),
    .A1(\cpuregs.regs[11][13] ),
    .S(_06359_),
    .X(_06363_));
 sky130_fd_sc_hd__clkbuf_1 _11835_ (.A(_06363_),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _11836_ (.A0(_06208_),
    .A1(\cpuregs.regs[11][14] ),
    .S(_06359_),
    .X(_06364_));
 sky130_fd_sc_hd__clkbuf_1 _11837_ (.A(_06364_),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _11838_ (.A0(_06216_),
    .A1(\cpuregs.regs[11][15] ),
    .S(_06359_),
    .X(_06365_));
 sky130_fd_sc_hd__clkbuf_1 _11839_ (.A(_06365_),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _11840_ (.A0(_06224_),
    .A1(\cpuregs.regs[11][16] ),
    .S(_06359_),
    .X(_06366_));
 sky130_fd_sc_hd__clkbuf_1 _11841_ (.A(_06366_),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _11842_ (.A0(_06232_),
    .A1(\cpuregs.regs[11][17] ),
    .S(_06359_),
    .X(_06367_));
 sky130_fd_sc_hd__clkbuf_1 _11843_ (.A(_06367_),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _11844_ (.A0(_06240_),
    .A1(\cpuregs.regs[11][18] ),
    .S(_06359_),
    .X(_06368_));
 sky130_fd_sc_hd__clkbuf_1 _11845_ (.A(_06368_),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _11846_ (.A0(_06248_),
    .A1(\cpuregs.regs[11][19] ),
    .S(_06359_),
    .X(_06369_));
 sky130_fd_sc_hd__clkbuf_1 _11847_ (.A(_06369_),
    .X(_00146_));
 sky130_fd_sc_hd__clkbuf_8 _11848_ (.A(_06347_),
    .X(_06370_));
 sky130_fd_sc_hd__mux2_1 _11849_ (.A0(_06257_),
    .A1(\cpuregs.regs[11][20] ),
    .S(_06370_),
    .X(_06371_));
 sky130_fd_sc_hd__clkbuf_1 _11850_ (.A(_06371_),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _11851_ (.A0(_06266_),
    .A1(\cpuregs.regs[11][21] ),
    .S(_06370_),
    .X(_06372_));
 sky130_fd_sc_hd__clkbuf_1 _11852_ (.A(_06372_),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _11853_ (.A0(_06274_),
    .A1(\cpuregs.regs[11][22] ),
    .S(_06370_),
    .X(_06373_));
 sky130_fd_sc_hd__clkbuf_1 _11854_ (.A(_06373_),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _11855_ (.A0(_06281_),
    .A1(\cpuregs.regs[11][23] ),
    .S(_06370_),
    .X(_06374_));
 sky130_fd_sc_hd__clkbuf_1 _11856_ (.A(_06374_),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _11857_ (.A0(_06289_),
    .A1(\cpuregs.regs[11][24] ),
    .S(_06370_),
    .X(_06375_));
 sky130_fd_sc_hd__clkbuf_1 _11858_ (.A(_06375_),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _11859_ (.A0(_06297_),
    .A1(\cpuregs.regs[11][25] ),
    .S(_06370_),
    .X(_06376_));
 sky130_fd_sc_hd__clkbuf_1 _11860_ (.A(_06376_),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _11861_ (.A0(_06304_),
    .A1(\cpuregs.regs[11][26] ),
    .S(_06370_),
    .X(_06377_));
 sky130_fd_sc_hd__clkbuf_1 _11862_ (.A(_06377_),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _11863_ (.A0(_06312_),
    .A1(\cpuregs.regs[11][27] ),
    .S(_06370_),
    .X(_06378_));
 sky130_fd_sc_hd__clkbuf_1 _11864_ (.A(_06378_),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _11865_ (.A0(_06320_),
    .A1(\cpuregs.regs[11][28] ),
    .S(_06370_),
    .X(_06379_));
 sky130_fd_sc_hd__clkbuf_1 _11866_ (.A(_06379_),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _11867_ (.A0(_06328_),
    .A1(\cpuregs.regs[11][29] ),
    .S(_06370_),
    .X(_06380_));
 sky130_fd_sc_hd__clkbuf_1 _11868_ (.A(_06380_),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _11869_ (.A0(_06336_),
    .A1(\cpuregs.regs[11][30] ),
    .S(_06347_),
    .X(_06381_));
 sky130_fd_sc_hd__clkbuf_1 _11870_ (.A(_06381_),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _11871_ (.A0(_06343_),
    .A1(\cpuregs.regs[11][31] ),
    .S(_06347_),
    .X(_06382_));
 sky130_fd_sc_hd__clkbuf_1 _11872_ (.A(_06382_),
    .X(_00158_));
 sky130_fd_sc_hd__nor2_4 _11873_ (.A(\cpuregs.waddr[1] ),
    .B(\cpuregs.waddr[0] ),
    .Y(_06383_));
 sky130_fd_sc_hd__and2_1 _11874_ (.A(\cpuregs.waddr[2] ),
    .B(_06083_),
    .X(_06384_));
 sky130_fd_sc_hd__and3b_4 _11875_ (.A_N(_06082_),
    .B(_06384_),
    .C(_06081_),
    .X(_06385_));
 sky130_fd_sc_hd__nand2_4 _11876_ (.A(_06383_),
    .B(_06385_),
    .Y(_06386_));
 sky130_fd_sc_hd__buf_6 _11877_ (.A(_06386_),
    .X(_06387_));
 sky130_fd_sc_hd__mux2_1 _11878_ (.A0(_06078_),
    .A1(\cpuregs.regs[20][0] ),
    .S(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__clkbuf_1 _11879_ (.A(_06388_),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _11880_ (.A0(_06096_),
    .A1(\cpuregs.regs[20][1] ),
    .S(_06387_),
    .X(_06389_));
 sky130_fd_sc_hd__clkbuf_1 _11881_ (.A(_06389_),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _11882_ (.A0(_06105_),
    .A1(\cpuregs.regs[20][2] ),
    .S(_06387_),
    .X(_06390_));
 sky130_fd_sc_hd__clkbuf_1 _11883_ (.A(_06390_),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _11884_ (.A0(_06114_),
    .A1(\cpuregs.regs[20][3] ),
    .S(_06387_),
    .X(_06391_));
 sky130_fd_sc_hd__clkbuf_1 _11885_ (.A(_06391_),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _11886_ (.A0(_06125_),
    .A1(\cpuregs.regs[20][4] ),
    .S(_06387_),
    .X(_06392_));
 sky130_fd_sc_hd__clkbuf_1 _11887_ (.A(_06392_),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _11888_ (.A0(_06132_),
    .A1(\cpuregs.regs[20][5] ),
    .S(_06387_),
    .X(_06393_));
 sky130_fd_sc_hd__clkbuf_1 _11889_ (.A(_06393_),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _11890_ (.A0(_06141_),
    .A1(\cpuregs.regs[20][6] ),
    .S(_06387_),
    .X(_06394_));
 sky130_fd_sc_hd__clkbuf_1 _11891_ (.A(_06394_),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _11892_ (.A0(_06150_),
    .A1(\cpuregs.regs[20][7] ),
    .S(_06387_),
    .X(_06395_));
 sky130_fd_sc_hd__clkbuf_1 _11893_ (.A(_06395_),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _11894_ (.A0(_06157_),
    .A1(\cpuregs.regs[20][8] ),
    .S(_06387_),
    .X(_06396_));
 sky130_fd_sc_hd__clkbuf_1 _11895_ (.A(_06396_),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _11896_ (.A0(_06166_),
    .A1(\cpuregs.regs[20][9] ),
    .S(_06387_),
    .X(_06397_));
 sky130_fd_sc_hd__clkbuf_1 _11897_ (.A(_06397_),
    .X(_00168_));
 sky130_fd_sc_hd__clkbuf_8 _11898_ (.A(_06386_),
    .X(_06398_));
 sky130_fd_sc_hd__mux2_1 _11899_ (.A0(_06175_),
    .A1(\cpuregs.regs[20][10] ),
    .S(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__clkbuf_1 _11900_ (.A(_06399_),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _11901_ (.A0(_06184_),
    .A1(\cpuregs.regs[20][11] ),
    .S(_06398_),
    .X(_06400_));
 sky130_fd_sc_hd__clkbuf_1 _11902_ (.A(_06400_),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _11903_ (.A0(_06193_),
    .A1(\cpuregs.regs[20][12] ),
    .S(_06398_),
    .X(_06401_));
 sky130_fd_sc_hd__clkbuf_1 _11904_ (.A(_06401_),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _11905_ (.A0(_06201_),
    .A1(\cpuregs.regs[20][13] ),
    .S(_06398_),
    .X(_06402_));
 sky130_fd_sc_hd__clkbuf_1 _11906_ (.A(_06402_),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _11907_ (.A0(_06208_),
    .A1(\cpuregs.regs[20][14] ),
    .S(_06398_),
    .X(_06403_));
 sky130_fd_sc_hd__clkbuf_1 _11908_ (.A(_06403_),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _11909_ (.A0(_06216_),
    .A1(\cpuregs.regs[20][15] ),
    .S(_06398_),
    .X(_06404_));
 sky130_fd_sc_hd__clkbuf_1 _11910_ (.A(_06404_),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _11911_ (.A0(_06224_),
    .A1(\cpuregs.regs[20][16] ),
    .S(_06398_),
    .X(_06405_));
 sky130_fd_sc_hd__clkbuf_1 _11912_ (.A(_06405_),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _11913_ (.A0(_06232_),
    .A1(\cpuregs.regs[20][17] ),
    .S(_06398_),
    .X(_06406_));
 sky130_fd_sc_hd__clkbuf_1 _11914_ (.A(_06406_),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _11915_ (.A0(_06240_),
    .A1(\cpuregs.regs[20][18] ),
    .S(_06398_),
    .X(_06407_));
 sky130_fd_sc_hd__clkbuf_1 _11916_ (.A(_06407_),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _11917_ (.A0(_06248_),
    .A1(\cpuregs.regs[20][19] ),
    .S(_06398_),
    .X(_06408_));
 sky130_fd_sc_hd__clkbuf_1 _11918_ (.A(_06408_),
    .X(_00178_));
 sky130_fd_sc_hd__buf_6 _11919_ (.A(_06386_),
    .X(_06409_));
 sky130_fd_sc_hd__mux2_1 _11920_ (.A0(_06257_),
    .A1(\cpuregs.regs[20][20] ),
    .S(_06409_),
    .X(_06410_));
 sky130_fd_sc_hd__clkbuf_1 _11921_ (.A(_06410_),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _11922_ (.A0(_06266_),
    .A1(\cpuregs.regs[20][21] ),
    .S(_06409_),
    .X(_06411_));
 sky130_fd_sc_hd__clkbuf_1 _11923_ (.A(_06411_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _11924_ (.A0(_06274_),
    .A1(\cpuregs.regs[20][22] ),
    .S(_06409_),
    .X(_06412_));
 sky130_fd_sc_hd__clkbuf_1 _11925_ (.A(_06412_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _11926_ (.A0(_06281_),
    .A1(\cpuregs.regs[20][23] ),
    .S(_06409_),
    .X(_06413_));
 sky130_fd_sc_hd__clkbuf_1 _11927_ (.A(_06413_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _11928_ (.A0(_06289_),
    .A1(\cpuregs.regs[20][24] ),
    .S(_06409_),
    .X(_06414_));
 sky130_fd_sc_hd__clkbuf_1 _11929_ (.A(_06414_),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _11930_ (.A0(_06297_),
    .A1(\cpuregs.regs[20][25] ),
    .S(_06409_),
    .X(_06415_));
 sky130_fd_sc_hd__clkbuf_1 _11931_ (.A(_06415_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _11932_ (.A0(_06304_),
    .A1(\cpuregs.regs[20][26] ),
    .S(_06409_),
    .X(_06416_));
 sky130_fd_sc_hd__clkbuf_1 _11933_ (.A(_06416_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _11934_ (.A0(_06312_),
    .A1(\cpuregs.regs[20][27] ),
    .S(_06409_),
    .X(_06417_));
 sky130_fd_sc_hd__clkbuf_1 _11935_ (.A(_06417_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _11936_ (.A0(_06320_),
    .A1(\cpuregs.regs[20][28] ),
    .S(_06409_),
    .X(_06418_));
 sky130_fd_sc_hd__clkbuf_1 _11937_ (.A(_06418_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _11938_ (.A0(_06328_),
    .A1(\cpuregs.regs[20][29] ),
    .S(_06409_),
    .X(_06419_));
 sky130_fd_sc_hd__clkbuf_1 _11939_ (.A(_06419_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _11940_ (.A0(_06336_),
    .A1(\cpuregs.regs[20][30] ),
    .S(_06386_),
    .X(_06420_));
 sky130_fd_sc_hd__clkbuf_1 _11941_ (.A(_06420_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _11942_ (.A0(_06343_),
    .A1(\cpuregs.regs[20][31] ),
    .S(_06386_),
    .X(_06421_));
 sky130_fd_sc_hd__clkbuf_1 _11943_ (.A(_06421_),
    .X(_00190_));
 sky130_fd_sc_hd__nor2b_4 _11944_ (.A(\cpuregs.waddr[1] ),
    .B_N(\cpuregs.waddr[0] ),
    .Y(_06422_));
 sky130_fd_sc_hd__nand2_4 _11945_ (.A(_06385_),
    .B(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__buf_6 _11946_ (.A(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__mux2_1 _11947_ (.A0(_06078_),
    .A1(\cpuregs.regs[21][0] ),
    .S(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__clkbuf_1 _11948_ (.A(_06425_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _11949_ (.A0(_06096_),
    .A1(\cpuregs.regs[21][1] ),
    .S(_06424_),
    .X(_06426_));
 sky130_fd_sc_hd__clkbuf_1 _11950_ (.A(_06426_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _11951_ (.A0(_06105_),
    .A1(\cpuregs.regs[21][2] ),
    .S(_06424_),
    .X(_06427_));
 sky130_fd_sc_hd__clkbuf_1 _11952_ (.A(_06427_),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _11953_ (.A0(_06114_),
    .A1(\cpuregs.regs[21][3] ),
    .S(_06424_),
    .X(_06428_));
 sky130_fd_sc_hd__clkbuf_1 _11954_ (.A(_06428_),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _11955_ (.A0(_06125_),
    .A1(\cpuregs.regs[21][4] ),
    .S(_06424_),
    .X(_06429_));
 sky130_fd_sc_hd__clkbuf_1 _11956_ (.A(_06429_),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _11957_ (.A0(_06132_),
    .A1(\cpuregs.regs[21][5] ),
    .S(_06424_),
    .X(_06430_));
 sky130_fd_sc_hd__clkbuf_1 _11958_ (.A(_06430_),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _11959_ (.A0(_06141_),
    .A1(\cpuregs.regs[21][6] ),
    .S(_06424_),
    .X(_06431_));
 sky130_fd_sc_hd__clkbuf_1 _11960_ (.A(_06431_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _11961_ (.A0(_06150_),
    .A1(\cpuregs.regs[21][7] ),
    .S(_06424_),
    .X(_06432_));
 sky130_fd_sc_hd__clkbuf_1 _11962_ (.A(_06432_),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _11963_ (.A0(_06157_),
    .A1(\cpuregs.regs[21][8] ),
    .S(_06424_),
    .X(_06433_));
 sky130_fd_sc_hd__clkbuf_1 _11964_ (.A(_06433_),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _11965_ (.A0(_06166_),
    .A1(\cpuregs.regs[21][9] ),
    .S(_06424_),
    .X(_06434_));
 sky130_fd_sc_hd__clkbuf_1 _11966_ (.A(_06434_),
    .X(_00200_));
 sky130_fd_sc_hd__clkbuf_8 _11967_ (.A(_06423_),
    .X(_06435_));
 sky130_fd_sc_hd__mux2_1 _11968_ (.A0(_06175_),
    .A1(\cpuregs.regs[21][10] ),
    .S(_06435_),
    .X(_06436_));
 sky130_fd_sc_hd__clkbuf_1 _11969_ (.A(_06436_),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _11970_ (.A0(_06184_),
    .A1(\cpuregs.regs[21][11] ),
    .S(_06435_),
    .X(_06437_));
 sky130_fd_sc_hd__clkbuf_1 _11971_ (.A(_06437_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _11972_ (.A0(_06193_),
    .A1(\cpuregs.regs[21][12] ),
    .S(_06435_),
    .X(_06438_));
 sky130_fd_sc_hd__clkbuf_1 _11973_ (.A(_06438_),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _11974_ (.A0(_06201_),
    .A1(\cpuregs.regs[21][13] ),
    .S(_06435_),
    .X(_06439_));
 sky130_fd_sc_hd__clkbuf_1 _11975_ (.A(_06439_),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _11976_ (.A0(_06208_),
    .A1(\cpuregs.regs[21][14] ),
    .S(_06435_),
    .X(_06440_));
 sky130_fd_sc_hd__clkbuf_1 _11977_ (.A(_06440_),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _11978_ (.A0(_06216_),
    .A1(\cpuregs.regs[21][15] ),
    .S(_06435_),
    .X(_06441_));
 sky130_fd_sc_hd__clkbuf_1 _11979_ (.A(_06441_),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _11980_ (.A0(_06224_),
    .A1(\cpuregs.regs[21][16] ),
    .S(_06435_),
    .X(_06442_));
 sky130_fd_sc_hd__clkbuf_1 _11981_ (.A(_06442_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _11982_ (.A0(_06232_),
    .A1(\cpuregs.regs[21][17] ),
    .S(_06435_),
    .X(_06443_));
 sky130_fd_sc_hd__clkbuf_1 _11983_ (.A(_06443_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _11984_ (.A0(_06240_),
    .A1(\cpuregs.regs[21][18] ),
    .S(_06435_),
    .X(_06444_));
 sky130_fd_sc_hd__clkbuf_1 _11985_ (.A(_06444_),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _11986_ (.A0(_06248_),
    .A1(\cpuregs.regs[21][19] ),
    .S(_06435_),
    .X(_06445_));
 sky130_fd_sc_hd__clkbuf_1 _11987_ (.A(_06445_),
    .X(_00210_));
 sky130_fd_sc_hd__buf_6 _11988_ (.A(_06423_),
    .X(_06446_));
 sky130_fd_sc_hd__mux2_1 _11989_ (.A0(_06257_),
    .A1(\cpuregs.regs[21][20] ),
    .S(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__clkbuf_1 _11990_ (.A(_06447_),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _11991_ (.A0(_06266_),
    .A1(\cpuregs.regs[21][21] ),
    .S(_06446_),
    .X(_06448_));
 sky130_fd_sc_hd__clkbuf_1 _11992_ (.A(_06448_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _11993_ (.A0(_06274_),
    .A1(\cpuregs.regs[21][22] ),
    .S(_06446_),
    .X(_06449_));
 sky130_fd_sc_hd__clkbuf_1 _11994_ (.A(_06449_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _11995_ (.A0(_06281_),
    .A1(\cpuregs.regs[21][23] ),
    .S(_06446_),
    .X(_06450_));
 sky130_fd_sc_hd__clkbuf_1 _11996_ (.A(_06450_),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _11997_ (.A0(_06289_),
    .A1(\cpuregs.regs[21][24] ),
    .S(_06446_),
    .X(_06451_));
 sky130_fd_sc_hd__clkbuf_1 _11998_ (.A(_06451_),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _11999_ (.A0(_06297_),
    .A1(\cpuregs.regs[21][25] ),
    .S(_06446_),
    .X(_06452_));
 sky130_fd_sc_hd__clkbuf_1 _12000_ (.A(_06452_),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_1 _12001_ (.A0(_06304_),
    .A1(\cpuregs.regs[21][26] ),
    .S(_06446_),
    .X(_06453_));
 sky130_fd_sc_hd__clkbuf_1 _12002_ (.A(_06453_),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _12003_ (.A0(_06312_),
    .A1(\cpuregs.regs[21][27] ),
    .S(_06446_),
    .X(_06454_));
 sky130_fd_sc_hd__clkbuf_1 _12004_ (.A(_06454_),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _12005_ (.A0(_06320_),
    .A1(\cpuregs.regs[21][28] ),
    .S(_06446_),
    .X(_06455_));
 sky130_fd_sc_hd__clkbuf_1 _12006_ (.A(_06455_),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _12007_ (.A0(_06328_),
    .A1(\cpuregs.regs[21][29] ),
    .S(_06446_),
    .X(_06456_));
 sky130_fd_sc_hd__clkbuf_1 _12008_ (.A(_06456_),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _12009_ (.A0(_06336_),
    .A1(\cpuregs.regs[21][30] ),
    .S(_06423_),
    .X(_06457_));
 sky130_fd_sc_hd__clkbuf_1 _12010_ (.A(_06457_),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _12011_ (.A0(_06343_),
    .A1(\cpuregs.regs[21][31] ),
    .S(_06423_),
    .X(_06458_));
 sky130_fd_sc_hd__clkbuf_1 _12012_ (.A(_06458_),
    .X(_00222_));
 sky130_fd_sc_hd__nand2_4 _12013_ (.A(_06080_),
    .B(_06385_),
    .Y(_06459_));
 sky130_fd_sc_hd__clkbuf_8 _12014_ (.A(_06459_),
    .X(_06460_));
 sky130_fd_sc_hd__mux2_1 _12015_ (.A0(_06078_),
    .A1(\cpuregs.regs[22][0] ),
    .S(_06460_),
    .X(_06461_));
 sky130_fd_sc_hd__clkbuf_1 _12016_ (.A(_06461_),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _12017_ (.A0(_06096_),
    .A1(\cpuregs.regs[22][1] ),
    .S(_06460_),
    .X(_06462_));
 sky130_fd_sc_hd__clkbuf_1 _12018_ (.A(_06462_),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _12019_ (.A0(_06105_),
    .A1(\cpuregs.regs[22][2] ),
    .S(_06460_),
    .X(_06463_));
 sky130_fd_sc_hd__clkbuf_1 _12020_ (.A(_06463_),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _12021_ (.A0(_06114_),
    .A1(\cpuregs.regs[22][3] ),
    .S(_06460_),
    .X(_06464_));
 sky130_fd_sc_hd__clkbuf_1 _12022_ (.A(_06464_),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _12023_ (.A0(_06125_),
    .A1(\cpuregs.regs[22][4] ),
    .S(_06460_),
    .X(_06465_));
 sky130_fd_sc_hd__clkbuf_1 _12024_ (.A(_06465_),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _12025_ (.A0(_06132_),
    .A1(\cpuregs.regs[22][5] ),
    .S(_06460_),
    .X(_06466_));
 sky130_fd_sc_hd__clkbuf_1 _12026_ (.A(_06466_),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _12027_ (.A0(_06141_),
    .A1(\cpuregs.regs[22][6] ),
    .S(_06460_),
    .X(_06467_));
 sky130_fd_sc_hd__clkbuf_1 _12028_ (.A(_06467_),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _12029_ (.A0(_06150_),
    .A1(\cpuregs.regs[22][7] ),
    .S(_06460_),
    .X(_06468_));
 sky130_fd_sc_hd__clkbuf_1 _12030_ (.A(_06468_),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _12031_ (.A0(_06157_),
    .A1(\cpuregs.regs[22][8] ),
    .S(_06460_),
    .X(_06469_));
 sky130_fd_sc_hd__clkbuf_1 _12032_ (.A(_06469_),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _12033_ (.A0(_06166_),
    .A1(\cpuregs.regs[22][9] ),
    .S(_06460_),
    .X(_06470_));
 sky130_fd_sc_hd__clkbuf_1 _12034_ (.A(_06470_),
    .X(_00232_));
 sky130_fd_sc_hd__clkbuf_8 _12035_ (.A(_06459_),
    .X(_06471_));
 sky130_fd_sc_hd__mux2_1 _12036_ (.A0(_06175_),
    .A1(\cpuregs.regs[22][10] ),
    .S(_06471_),
    .X(_06472_));
 sky130_fd_sc_hd__clkbuf_1 _12037_ (.A(_06472_),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _12038_ (.A0(_06184_),
    .A1(\cpuregs.regs[22][11] ),
    .S(_06471_),
    .X(_06473_));
 sky130_fd_sc_hd__clkbuf_1 _12039_ (.A(_06473_),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _12040_ (.A0(_06193_),
    .A1(\cpuregs.regs[22][12] ),
    .S(_06471_),
    .X(_06474_));
 sky130_fd_sc_hd__clkbuf_1 _12041_ (.A(_06474_),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _12042_ (.A0(_06201_),
    .A1(\cpuregs.regs[22][13] ),
    .S(_06471_),
    .X(_06475_));
 sky130_fd_sc_hd__clkbuf_1 _12043_ (.A(_06475_),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _12044_ (.A0(_06208_),
    .A1(\cpuregs.regs[22][14] ),
    .S(_06471_),
    .X(_06476_));
 sky130_fd_sc_hd__clkbuf_1 _12045_ (.A(_06476_),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _12046_ (.A0(_06216_),
    .A1(\cpuregs.regs[22][15] ),
    .S(_06471_),
    .X(_06477_));
 sky130_fd_sc_hd__clkbuf_1 _12047_ (.A(_06477_),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _12048_ (.A0(_06224_),
    .A1(\cpuregs.regs[22][16] ),
    .S(_06471_),
    .X(_06478_));
 sky130_fd_sc_hd__clkbuf_1 _12049_ (.A(_06478_),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _12050_ (.A0(_06232_),
    .A1(\cpuregs.regs[22][17] ),
    .S(_06471_),
    .X(_06479_));
 sky130_fd_sc_hd__clkbuf_1 _12051_ (.A(_06479_),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _12052_ (.A0(_06240_),
    .A1(\cpuregs.regs[22][18] ),
    .S(_06471_),
    .X(_06480_));
 sky130_fd_sc_hd__clkbuf_1 _12053_ (.A(_06480_),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _12054_ (.A0(_06248_),
    .A1(\cpuregs.regs[22][19] ),
    .S(_06471_),
    .X(_06481_));
 sky130_fd_sc_hd__clkbuf_1 _12055_ (.A(_06481_),
    .X(_00242_));
 sky130_fd_sc_hd__buf_6 _12056_ (.A(_06459_),
    .X(_06482_));
 sky130_fd_sc_hd__mux2_1 _12057_ (.A0(_06257_),
    .A1(\cpuregs.regs[22][20] ),
    .S(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__clkbuf_1 _12058_ (.A(_06483_),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _12059_ (.A0(_06266_),
    .A1(\cpuregs.regs[22][21] ),
    .S(_06482_),
    .X(_06484_));
 sky130_fd_sc_hd__clkbuf_1 _12060_ (.A(_06484_),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _12061_ (.A0(_06274_),
    .A1(\cpuregs.regs[22][22] ),
    .S(_06482_),
    .X(_06485_));
 sky130_fd_sc_hd__clkbuf_1 _12062_ (.A(_06485_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _12063_ (.A0(_06281_),
    .A1(\cpuregs.regs[22][23] ),
    .S(_06482_),
    .X(_06486_));
 sky130_fd_sc_hd__clkbuf_1 _12064_ (.A(_06486_),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _12065_ (.A0(_06289_),
    .A1(\cpuregs.regs[22][24] ),
    .S(_06482_),
    .X(_06487_));
 sky130_fd_sc_hd__clkbuf_1 _12066_ (.A(_06487_),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _12067_ (.A0(_06297_),
    .A1(\cpuregs.regs[22][25] ),
    .S(_06482_),
    .X(_06488_));
 sky130_fd_sc_hd__clkbuf_1 _12068_ (.A(_06488_),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _12069_ (.A0(_06304_),
    .A1(\cpuregs.regs[22][26] ),
    .S(_06482_),
    .X(_06489_));
 sky130_fd_sc_hd__clkbuf_1 _12070_ (.A(_06489_),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _12071_ (.A0(_06312_),
    .A1(\cpuregs.regs[22][27] ),
    .S(_06482_),
    .X(_06490_));
 sky130_fd_sc_hd__clkbuf_1 _12072_ (.A(_06490_),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _12073_ (.A0(_06320_),
    .A1(\cpuregs.regs[22][28] ),
    .S(_06482_),
    .X(_06491_));
 sky130_fd_sc_hd__clkbuf_1 _12074_ (.A(_06491_),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _12075_ (.A0(_06328_),
    .A1(\cpuregs.regs[22][29] ),
    .S(_06482_),
    .X(_06492_));
 sky130_fd_sc_hd__clkbuf_1 _12076_ (.A(_06492_),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _12077_ (.A0(_06336_),
    .A1(\cpuregs.regs[22][30] ),
    .S(_06459_),
    .X(_06493_));
 sky130_fd_sc_hd__clkbuf_1 _12078_ (.A(_06493_),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _12079_ (.A0(_06343_),
    .A1(\cpuregs.regs[22][31] ),
    .S(_06459_),
    .X(_06494_));
 sky130_fd_sc_hd__clkbuf_1 _12080_ (.A(_06494_),
    .X(_00254_));
 sky130_fd_sc_hd__nand2_4 _12081_ (.A(_06346_),
    .B(_06385_),
    .Y(_06495_));
 sky130_fd_sc_hd__buf_6 _12082_ (.A(_06495_),
    .X(_06496_));
 sky130_fd_sc_hd__mux2_1 _12083_ (.A0(_06078_),
    .A1(\cpuregs.regs[23][0] ),
    .S(_06496_),
    .X(_06497_));
 sky130_fd_sc_hd__clkbuf_1 _12084_ (.A(_06497_),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _12085_ (.A0(_06096_),
    .A1(\cpuregs.regs[23][1] ),
    .S(_06496_),
    .X(_06498_));
 sky130_fd_sc_hd__clkbuf_1 _12086_ (.A(_06498_),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _12087_ (.A0(_06105_),
    .A1(\cpuregs.regs[23][2] ),
    .S(_06496_),
    .X(_06499_));
 sky130_fd_sc_hd__clkbuf_1 _12088_ (.A(_06499_),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _12089_ (.A0(_06114_),
    .A1(\cpuregs.regs[23][3] ),
    .S(_06496_),
    .X(_06500_));
 sky130_fd_sc_hd__clkbuf_1 _12090_ (.A(_06500_),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _12091_ (.A0(_06125_),
    .A1(\cpuregs.regs[23][4] ),
    .S(_06496_),
    .X(_06501_));
 sky130_fd_sc_hd__clkbuf_1 _12092_ (.A(_06501_),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _12093_ (.A0(_06132_),
    .A1(\cpuregs.regs[23][5] ),
    .S(_06496_),
    .X(_06502_));
 sky130_fd_sc_hd__clkbuf_1 _12094_ (.A(_06502_),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _12095_ (.A0(_06141_),
    .A1(\cpuregs.regs[23][6] ),
    .S(_06496_),
    .X(_06503_));
 sky130_fd_sc_hd__clkbuf_1 _12096_ (.A(_06503_),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _12097_ (.A0(_06150_),
    .A1(\cpuregs.regs[23][7] ),
    .S(_06496_),
    .X(_06504_));
 sky130_fd_sc_hd__clkbuf_1 _12098_ (.A(_06504_),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _12099_ (.A0(_06157_),
    .A1(\cpuregs.regs[23][8] ),
    .S(_06496_),
    .X(_06505_));
 sky130_fd_sc_hd__clkbuf_1 _12100_ (.A(_06505_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _12101_ (.A0(_06166_),
    .A1(\cpuregs.regs[23][9] ),
    .S(_06496_),
    .X(_06506_));
 sky130_fd_sc_hd__clkbuf_1 _12102_ (.A(_06506_),
    .X(_00264_));
 sky130_fd_sc_hd__clkbuf_8 _12103_ (.A(_06495_),
    .X(_06507_));
 sky130_fd_sc_hd__mux2_1 _12104_ (.A0(_06175_),
    .A1(\cpuregs.regs[23][10] ),
    .S(_06507_),
    .X(_06508_));
 sky130_fd_sc_hd__clkbuf_1 _12105_ (.A(_06508_),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _12106_ (.A0(_06184_),
    .A1(\cpuregs.regs[23][11] ),
    .S(_06507_),
    .X(_06509_));
 sky130_fd_sc_hd__clkbuf_1 _12107_ (.A(_06509_),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _12108_ (.A0(_06193_),
    .A1(\cpuregs.regs[23][12] ),
    .S(_06507_),
    .X(_06510_));
 sky130_fd_sc_hd__clkbuf_1 _12109_ (.A(_06510_),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _12110_ (.A0(_06201_),
    .A1(\cpuregs.regs[23][13] ),
    .S(_06507_),
    .X(_06511_));
 sky130_fd_sc_hd__clkbuf_1 _12111_ (.A(_06511_),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _12112_ (.A0(_06208_),
    .A1(\cpuregs.regs[23][14] ),
    .S(_06507_),
    .X(_06512_));
 sky130_fd_sc_hd__clkbuf_1 _12113_ (.A(_06512_),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _12114_ (.A0(_06216_),
    .A1(\cpuregs.regs[23][15] ),
    .S(_06507_),
    .X(_06513_));
 sky130_fd_sc_hd__clkbuf_1 _12115_ (.A(_06513_),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _12116_ (.A0(_06224_),
    .A1(\cpuregs.regs[23][16] ),
    .S(_06507_),
    .X(_06514_));
 sky130_fd_sc_hd__clkbuf_1 _12117_ (.A(_06514_),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _12118_ (.A0(_06232_),
    .A1(\cpuregs.regs[23][17] ),
    .S(_06507_),
    .X(_06515_));
 sky130_fd_sc_hd__clkbuf_1 _12119_ (.A(_06515_),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _12120_ (.A0(_06240_),
    .A1(\cpuregs.regs[23][18] ),
    .S(_06507_),
    .X(_06516_));
 sky130_fd_sc_hd__clkbuf_1 _12121_ (.A(_06516_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _12122_ (.A0(_06248_),
    .A1(\cpuregs.regs[23][19] ),
    .S(_06507_),
    .X(_06517_));
 sky130_fd_sc_hd__clkbuf_1 _12123_ (.A(_06517_),
    .X(_00274_));
 sky130_fd_sc_hd__buf_6 _12124_ (.A(_06495_),
    .X(_06518_));
 sky130_fd_sc_hd__mux2_1 _12125_ (.A0(_06257_),
    .A1(\cpuregs.regs[23][20] ),
    .S(_06518_),
    .X(_06519_));
 sky130_fd_sc_hd__clkbuf_1 _12126_ (.A(_06519_),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _12127_ (.A0(_06266_),
    .A1(\cpuregs.regs[23][21] ),
    .S(_06518_),
    .X(_06520_));
 sky130_fd_sc_hd__clkbuf_1 _12128_ (.A(_06520_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _12129_ (.A0(_06274_),
    .A1(\cpuregs.regs[23][22] ),
    .S(_06518_),
    .X(_06521_));
 sky130_fd_sc_hd__clkbuf_1 _12130_ (.A(_06521_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _12131_ (.A0(_06281_),
    .A1(\cpuregs.regs[23][23] ),
    .S(_06518_),
    .X(_06522_));
 sky130_fd_sc_hd__clkbuf_1 _12132_ (.A(_06522_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _12133_ (.A0(_06289_),
    .A1(\cpuregs.regs[23][24] ),
    .S(_06518_),
    .X(_06523_));
 sky130_fd_sc_hd__clkbuf_1 _12134_ (.A(_06523_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _12135_ (.A0(_06297_),
    .A1(\cpuregs.regs[23][25] ),
    .S(_06518_),
    .X(_06524_));
 sky130_fd_sc_hd__clkbuf_1 _12136_ (.A(_06524_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _12137_ (.A0(_06304_),
    .A1(\cpuregs.regs[23][26] ),
    .S(_06518_),
    .X(_06525_));
 sky130_fd_sc_hd__clkbuf_1 _12138_ (.A(_06525_),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _12139_ (.A0(_06312_),
    .A1(\cpuregs.regs[23][27] ),
    .S(_06518_),
    .X(_06526_));
 sky130_fd_sc_hd__clkbuf_1 _12140_ (.A(_06526_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _12141_ (.A0(_06320_),
    .A1(\cpuregs.regs[23][28] ),
    .S(_06518_),
    .X(_06527_));
 sky130_fd_sc_hd__clkbuf_1 _12142_ (.A(_06527_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _12143_ (.A0(_06328_),
    .A1(\cpuregs.regs[23][29] ),
    .S(_06518_),
    .X(_06528_));
 sky130_fd_sc_hd__clkbuf_1 _12144_ (.A(_06528_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _12145_ (.A0(_06336_),
    .A1(\cpuregs.regs[23][30] ),
    .S(_06495_),
    .X(_06529_));
 sky130_fd_sc_hd__clkbuf_1 _12146_ (.A(_06529_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _12147_ (.A0(_06343_),
    .A1(\cpuregs.regs[23][31] ),
    .S(_06495_),
    .X(_06530_));
 sky130_fd_sc_hd__clkbuf_1 _12148_ (.A(_06530_),
    .X(_00286_));
 sky130_fd_sc_hd__buf_2 _12149_ (.A(_06077_),
    .X(_06531_));
 sky130_fd_sc_hd__nand4b_4 _12150_ (.A_N(\cpuregs.waddr[2] ),
    .B(_06081_),
    .C(_06082_),
    .D(_06083_),
    .Y(_06532_));
 sky130_fd_sc_hd__nor3_4 _12151_ (.A(\cpuregs.waddr[1] ),
    .B(\cpuregs.waddr[0] ),
    .C(_06532_),
    .Y(_06533_));
 sky130_fd_sc_hd__clkbuf_8 _12152_ (.A(_06533_),
    .X(_06534_));
 sky130_fd_sc_hd__mux2_1 _12153_ (.A0(\cpuregs.regs[24][0] ),
    .A1(_06531_),
    .S(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__clkbuf_1 _12154_ (.A(_06535_),
    .X(_00287_));
 sky130_fd_sc_hd__buf_2 _12155_ (.A(_06095_),
    .X(_06536_));
 sky130_fd_sc_hd__mux2_1 _12156_ (.A0(\cpuregs.regs[24][1] ),
    .A1(_06536_),
    .S(_06534_),
    .X(_06537_));
 sky130_fd_sc_hd__clkbuf_1 _12157_ (.A(_06537_),
    .X(_00288_));
 sky130_fd_sc_hd__buf_2 _12158_ (.A(_06104_),
    .X(_06538_));
 sky130_fd_sc_hd__mux2_1 _12159_ (.A0(\cpuregs.regs[24][2] ),
    .A1(_06538_),
    .S(_06534_),
    .X(_06539_));
 sky130_fd_sc_hd__clkbuf_1 _12160_ (.A(_06539_),
    .X(_00289_));
 sky130_fd_sc_hd__buf_2 _12161_ (.A(_06113_),
    .X(_06540_));
 sky130_fd_sc_hd__mux2_1 _12162_ (.A0(\cpuregs.regs[24][3] ),
    .A1(_06540_),
    .S(_06534_),
    .X(_06541_));
 sky130_fd_sc_hd__clkbuf_1 _12163_ (.A(_06541_),
    .X(_00290_));
 sky130_fd_sc_hd__buf_2 _12164_ (.A(_06124_),
    .X(_06542_));
 sky130_fd_sc_hd__mux2_1 _12165_ (.A0(\cpuregs.regs[24][4] ),
    .A1(_06542_),
    .S(_06534_),
    .X(_06543_));
 sky130_fd_sc_hd__clkbuf_1 _12166_ (.A(_06543_),
    .X(_00291_));
 sky130_fd_sc_hd__buf_2 _12167_ (.A(_06131_),
    .X(_06544_));
 sky130_fd_sc_hd__mux2_1 _12168_ (.A0(\cpuregs.regs[24][5] ),
    .A1(_06544_),
    .S(_06534_),
    .X(_06545_));
 sky130_fd_sc_hd__clkbuf_1 _12169_ (.A(_06545_),
    .X(_00292_));
 sky130_fd_sc_hd__buf_2 _12170_ (.A(_06140_),
    .X(_06546_));
 sky130_fd_sc_hd__mux2_1 _12171_ (.A0(\cpuregs.regs[24][6] ),
    .A1(_06546_),
    .S(_06534_),
    .X(_06547_));
 sky130_fd_sc_hd__clkbuf_1 _12172_ (.A(_06547_),
    .X(_00293_));
 sky130_fd_sc_hd__buf_2 _12173_ (.A(_06149_),
    .X(_06548_));
 sky130_fd_sc_hd__mux2_1 _12174_ (.A0(\cpuregs.regs[24][7] ),
    .A1(_06548_),
    .S(_06534_),
    .X(_06549_));
 sky130_fd_sc_hd__clkbuf_1 _12175_ (.A(_06549_),
    .X(_00294_));
 sky130_fd_sc_hd__buf_2 _12176_ (.A(_06156_),
    .X(_06550_));
 sky130_fd_sc_hd__mux2_1 _12177_ (.A0(\cpuregs.regs[24][8] ),
    .A1(_06550_),
    .S(_06534_),
    .X(_06551_));
 sky130_fd_sc_hd__clkbuf_1 _12178_ (.A(_06551_),
    .X(_00295_));
 sky130_fd_sc_hd__buf_2 _12179_ (.A(_06165_),
    .X(_06552_));
 sky130_fd_sc_hd__mux2_1 _12180_ (.A0(\cpuregs.regs[24][9] ),
    .A1(_06552_),
    .S(_06534_),
    .X(_06553_));
 sky130_fd_sc_hd__clkbuf_1 _12181_ (.A(_06553_),
    .X(_00296_));
 sky130_fd_sc_hd__clkbuf_4 _12182_ (.A(_06174_),
    .X(_06554_));
 sky130_fd_sc_hd__clkbuf_8 _12183_ (.A(_06533_),
    .X(_06555_));
 sky130_fd_sc_hd__mux2_1 _12184_ (.A0(\cpuregs.regs[24][10] ),
    .A1(_06554_),
    .S(_06555_),
    .X(_06556_));
 sky130_fd_sc_hd__clkbuf_1 _12185_ (.A(_06556_),
    .X(_00297_));
 sky130_fd_sc_hd__buf_2 _12186_ (.A(_06183_),
    .X(_06557_));
 sky130_fd_sc_hd__mux2_1 _12187_ (.A0(\cpuregs.regs[24][11] ),
    .A1(_06557_),
    .S(_06555_),
    .X(_06558_));
 sky130_fd_sc_hd__clkbuf_1 _12188_ (.A(_06558_),
    .X(_00298_));
 sky130_fd_sc_hd__buf_2 _12189_ (.A(_06192_),
    .X(_06559_));
 sky130_fd_sc_hd__mux2_1 _12190_ (.A0(\cpuregs.regs[24][12] ),
    .A1(_06559_),
    .S(_06555_),
    .X(_06560_));
 sky130_fd_sc_hd__clkbuf_1 _12191_ (.A(_06560_),
    .X(_00299_));
 sky130_fd_sc_hd__buf_2 _12192_ (.A(_06200_),
    .X(_06561_));
 sky130_fd_sc_hd__mux2_1 _12193_ (.A0(\cpuregs.regs[24][13] ),
    .A1(_06561_),
    .S(_06555_),
    .X(_06562_));
 sky130_fd_sc_hd__clkbuf_1 _12194_ (.A(_06562_),
    .X(_00300_));
 sky130_fd_sc_hd__buf_2 _12195_ (.A(_06207_),
    .X(_06563_));
 sky130_fd_sc_hd__mux2_1 _12196_ (.A0(\cpuregs.regs[24][14] ),
    .A1(_06563_),
    .S(_06555_),
    .X(_06564_));
 sky130_fd_sc_hd__clkbuf_1 _12197_ (.A(_06564_),
    .X(_00301_));
 sky130_fd_sc_hd__buf_2 _12198_ (.A(_06215_),
    .X(_06565_));
 sky130_fd_sc_hd__mux2_1 _12199_ (.A0(\cpuregs.regs[24][15] ),
    .A1(_06565_),
    .S(_06555_),
    .X(_06566_));
 sky130_fd_sc_hd__clkbuf_1 _12200_ (.A(_06566_),
    .X(_00302_));
 sky130_fd_sc_hd__buf_2 _12201_ (.A(_06223_),
    .X(_06567_));
 sky130_fd_sc_hd__mux2_1 _12202_ (.A0(\cpuregs.regs[24][16] ),
    .A1(_06567_),
    .S(_06555_),
    .X(_06568_));
 sky130_fd_sc_hd__clkbuf_1 _12203_ (.A(_06568_),
    .X(_00303_));
 sky130_fd_sc_hd__buf_2 _12204_ (.A(_06231_),
    .X(_06569_));
 sky130_fd_sc_hd__mux2_1 _12205_ (.A0(\cpuregs.regs[24][17] ),
    .A1(_06569_),
    .S(_06555_),
    .X(_06570_));
 sky130_fd_sc_hd__clkbuf_1 _12206_ (.A(_06570_),
    .X(_00304_));
 sky130_fd_sc_hd__clkbuf_4 _12207_ (.A(_06239_),
    .X(_06571_));
 sky130_fd_sc_hd__mux2_1 _12208_ (.A0(\cpuregs.regs[24][18] ),
    .A1(_06571_),
    .S(_06555_),
    .X(_06572_));
 sky130_fd_sc_hd__clkbuf_1 _12209_ (.A(_06572_),
    .X(_00305_));
 sky130_fd_sc_hd__buf_2 _12210_ (.A(_06247_),
    .X(_06573_));
 sky130_fd_sc_hd__mux2_1 _12211_ (.A0(\cpuregs.regs[24][19] ),
    .A1(_06573_),
    .S(_06555_),
    .X(_06574_));
 sky130_fd_sc_hd__clkbuf_1 _12212_ (.A(_06574_),
    .X(_00306_));
 sky130_fd_sc_hd__buf_2 _12213_ (.A(_06256_),
    .X(_06575_));
 sky130_fd_sc_hd__clkbuf_8 _12214_ (.A(_06533_),
    .X(_06576_));
 sky130_fd_sc_hd__mux2_1 _12215_ (.A0(\cpuregs.regs[24][20] ),
    .A1(_06575_),
    .S(_06576_),
    .X(_06577_));
 sky130_fd_sc_hd__clkbuf_1 _12216_ (.A(_06577_),
    .X(_00307_));
 sky130_fd_sc_hd__buf_2 _12217_ (.A(_06265_),
    .X(_06578_));
 sky130_fd_sc_hd__mux2_1 _12218_ (.A0(\cpuregs.regs[24][21] ),
    .A1(_06578_),
    .S(_06576_),
    .X(_06579_));
 sky130_fd_sc_hd__clkbuf_1 _12219_ (.A(_06579_),
    .X(_00308_));
 sky130_fd_sc_hd__buf_2 _12220_ (.A(_06273_),
    .X(_06580_));
 sky130_fd_sc_hd__mux2_1 _12221_ (.A0(\cpuregs.regs[24][22] ),
    .A1(_06580_),
    .S(_06576_),
    .X(_06581_));
 sky130_fd_sc_hd__clkbuf_1 _12222_ (.A(_06581_),
    .X(_00309_));
 sky130_fd_sc_hd__buf_2 _12223_ (.A(_06280_),
    .X(_06582_));
 sky130_fd_sc_hd__mux2_1 _12224_ (.A0(\cpuregs.regs[24][23] ),
    .A1(_06582_),
    .S(_06576_),
    .X(_06583_));
 sky130_fd_sc_hd__clkbuf_1 _12225_ (.A(_06583_),
    .X(_00310_));
 sky130_fd_sc_hd__buf_2 _12226_ (.A(_06288_),
    .X(_06584_));
 sky130_fd_sc_hd__mux2_1 _12227_ (.A0(\cpuregs.regs[24][24] ),
    .A1(_06584_),
    .S(_06576_),
    .X(_06585_));
 sky130_fd_sc_hd__clkbuf_1 _12228_ (.A(_06585_),
    .X(_00311_));
 sky130_fd_sc_hd__buf_2 _12229_ (.A(_06296_),
    .X(_06586_));
 sky130_fd_sc_hd__mux2_1 _12230_ (.A0(\cpuregs.regs[24][25] ),
    .A1(_06586_),
    .S(_06576_),
    .X(_06587_));
 sky130_fd_sc_hd__clkbuf_1 _12231_ (.A(_06587_),
    .X(_00312_));
 sky130_fd_sc_hd__buf_2 _12232_ (.A(_06303_),
    .X(_06588_));
 sky130_fd_sc_hd__mux2_1 _12233_ (.A0(\cpuregs.regs[24][26] ),
    .A1(_06588_),
    .S(_06576_),
    .X(_06589_));
 sky130_fd_sc_hd__clkbuf_1 _12234_ (.A(_06589_),
    .X(_00313_));
 sky130_fd_sc_hd__buf_2 _12235_ (.A(_06311_),
    .X(_06590_));
 sky130_fd_sc_hd__mux2_1 _12236_ (.A0(\cpuregs.regs[24][27] ),
    .A1(_06590_),
    .S(_06576_),
    .X(_06591_));
 sky130_fd_sc_hd__clkbuf_1 _12237_ (.A(_06591_),
    .X(_00314_));
 sky130_fd_sc_hd__buf_2 _12238_ (.A(_06319_),
    .X(_06592_));
 sky130_fd_sc_hd__mux2_1 _12239_ (.A0(\cpuregs.regs[24][28] ),
    .A1(_06592_),
    .S(_06576_),
    .X(_06593_));
 sky130_fd_sc_hd__clkbuf_1 _12240_ (.A(_06593_),
    .X(_00315_));
 sky130_fd_sc_hd__buf_2 _12241_ (.A(_06327_),
    .X(_06594_));
 sky130_fd_sc_hd__mux2_1 _12242_ (.A0(\cpuregs.regs[24][29] ),
    .A1(_06594_),
    .S(_06576_),
    .X(_06595_));
 sky130_fd_sc_hd__clkbuf_1 _12243_ (.A(_06595_),
    .X(_00316_));
 sky130_fd_sc_hd__buf_2 _12244_ (.A(_06335_),
    .X(_06596_));
 sky130_fd_sc_hd__mux2_1 _12245_ (.A0(\cpuregs.regs[24][30] ),
    .A1(_06596_),
    .S(_06533_),
    .X(_06597_));
 sky130_fd_sc_hd__clkbuf_1 _12246_ (.A(_06597_),
    .X(_00317_));
 sky130_fd_sc_hd__buf_2 _12247_ (.A(_06342_),
    .X(_06598_));
 sky130_fd_sc_hd__mux2_1 _12248_ (.A0(\cpuregs.regs[24][31] ),
    .A1(_06598_),
    .S(_06533_),
    .X(_06599_));
 sky130_fd_sc_hd__clkbuf_1 _12249_ (.A(_06599_),
    .X(_00318_));
 sky130_fd_sc_hd__nand2_1 _12250_ (.A(_06083_),
    .B(_06422_),
    .Y(_06600_));
 sky130_fd_sc_hd__inv_2 _12251_ (.A(_06600_),
    .Y(_06601_));
 sky130_fd_sc_hd__and4b_1 _12252_ (.A_N(\cpuregs.waddr[2] ),
    .B(\cpuregs.waddr[4] ),
    .C(\cpuregs.waddr[3] ),
    .D(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__clkbuf_4 _12253_ (.A(_06602_),
    .X(_06603_));
 sky130_fd_sc_hd__clkbuf_8 _12254_ (.A(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__mux2_1 _12255_ (.A0(\cpuregs.regs[25][0] ),
    .A1(_06531_),
    .S(_06604_),
    .X(_06605_));
 sky130_fd_sc_hd__clkbuf_1 _12256_ (.A(_06605_),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _12257_ (.A0(\cpuregs.regs[25][1] ),
    .A1(_06536_),
    .S(_06604_),
    .X(_06606_));
 sky130_fd_sc_hd__clkbuf_1 _12258_ (.A(_06606_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _12259_ (.A0(\cpuregs.regs[25][2] ),
    .A1(_06538_),
    .S(_06604_),
    .X(_06607_));
 sky130_fd_sc_hd__clkbuf_1 _12260_ (.A(_06607_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _12261_ (.A0(\cpuregs.regs[25][3] ),
    .A1(_06540_),
    .S(_06604_),
    .X(_06608_));
 sky130_fd_sc_hd__clkbuf_1 _12262_ (.A(_06608_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _12263_ (.A0(\cpuregs.regs[25][4] ),
    .A1(_06542_),
    .S(_06604_),
    .X(_06609_));
 sky130_fd_sc_hd__clkbuf_1 _12264_ (.A(_06609_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _12265_ (.A0(\cpuregs.regs[25][5] ),
    .A1(_06544_),
    .S(_06604_),
    .X(_06610_));
 sky130_fd_sc_hd__clkbuf_1 _12266_ (.A(_06610_),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _12267_ (.A0(\cpuregs.regs[25][6] ),
    .A1(_06546_),
    .S(_06604_),
    .X(_06611_));
 sky130_fd_sc_hd__clkbuf_1 _12268_ (.A(_06611_),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _12269_ (.A0(\cpuregs.regs[25][7] ),
    .A1(_06548_),
    .S(_06604_),
    .X(_06612_));
 sky130_fd_sc_hd__clkbuf_1 _12270_ (.A(_06612_),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _12271_ (.A0(\cpuregs.regs[25][8] ),
    .A1(_06550_),
    .S(_06604_),
    .X(_06613_));
 sky130_fd_sc_hd__clkbuf_1 _12272_ (.A(_06613_),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _12273_ (.A0(\cpuregs.regs[25][9] ),
    .A1(_06552_),
    .S(_06604_),
    .X(_06614_));
 sky130_fd_sc_hd__clkbuf_1 _12274_ (.A(_06614_),
    .X(_00328_));
 sky130_fd_sc_hd__clkbuf_8 _12275_ (.A(_06603_),
    .X(_06615_));
 sky130_fd_sc_hd__mux2_1 _12276_ (.A0(\cpuregs.regs[25][10] ),
    .A1(_06554_),
    .S(_06615_),
    .X(_06616_));
 sky130_fd_sc_hd__clkbuf_1 _12277_ (.A(_06616_),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _12278_ (.A0(\cpuregs.regs[25][11] ),
    .A1(_06557_),
    .S(_06615_),
    .X(_06617_));
 sky130_fd_sc_hd__clkbuf_1 _12279_ (.A(_06617_),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _12280_ (.A0(\cpuregs.regs[25][12] ),
    .A1(_06559_),
    .S(_06615_),
    .X(_06618_));
 sky130_fd_sc_hd__clkbuf_1 _12281_ (.A(_06618_),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _12282_ (.A0(\cpuregs.regs[25][13] ),
    .A1(_06561_),
    .S(_06615_),
    .X(_06619_));
 sky130_fd_sc_hd__clkbuf_1 _12283_ (.A(_06619_),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _12284_ (.A0(\cpuregs.regs[25][14] ),
    .A1(_06563_),
    .S(_06615_),
    .X(_06620_));
 sky130_fd_sc_hd__clkbuf_1 _12285_ (.A(_06620_),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _12286_ (.A0(\cpuregs.regs[25][15] ),
    .A1(_06565_),
    .S(_06615_),
    .X(_06621_));
 sky130_fd_sc_hd__clkbuf_1 _12287_ (.A(_06621_),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _12288_ (.A0(\cpuregs.regs[25][16] ),
    .A1(_06567_),
    .S(_06615_),
    .X(_06622_));
 sky130_fd_sc_hd__clkbuf_1 _12289_ (.A(_06622_),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _12290_ (.A0(\cpuregs.regs[25][17] ),
    .A1(_06569_),
    .S(_06615_),
    .X(_06623_));
 sky130_fd_sc_hd__clkbuf_1 _12291_ (.A(_06623_),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _12292_ (.A0(\cpuregs.regs[25][18] ),
    .A1(_06571_),
    .S(_06615_),
    .X(_06624_));
 sky130_fd_sc_hd__clkbuf_1 _12293_ (.A(_06624_),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _12294_ (.A0(\cpuregs.regs[25][19] ),
    .A1(_06573_),
    .S(_06615_),
    .X(_06625_));
 sky130_fd_sc_hd__clkbuf_1 _12295_ (.A(_06625_),
    .X(_00338_));
 sky130_fd_sc_hd__clkbuf_8 _12296_ (.A(_06603_),
    .X(_06626_));
 sky130_fd_sc_hd__mux2_1 _12297_ (.A0(\cpuregs.regs[25][20] ),
    .A1(_06575_),
    .S(_06626_),
    .X(_06627_));
 sky130_fd_sc_hd__clkbuf_1 _12298_ (.A(_06627_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _12299_ (.A0(\cpuregs.regs[25][21] ),
    .A1(_06578_),
    .S(_06626_),
    .X(_06628_));
 sky130_fd_sc_hd__clkbuf_1 _12300_ (.A(_06628_),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _12301_ (.A0(\cpuregs.regs[25][22] ),
    .A1(_06580_),
    .S(_06626_),
    .X(_06629_));
 sky130_fd_sc_hd__clkbuf_1 _12302_ (.A(_06629_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _12303_ (.A0(\cpuregs.regs[25][23] ),
    .A1(_06582_),
    .S(_06626_),
    .X(_06630_));
 sky130_fd_sc_hd__clkbuf_1 _12304_ (.A(_06630_),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_1 _12305_ (.A0(\cpuregs.regs[25][24] ),
    .A1(_06584_),
    .S(_06626_),
    .X(_06631_));
 sky130_fd_sc_hd__clkbuf_1 _12306_ (.A(_06631_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _12307_ (.A0(\cpuregs.regs[25][25] ),
    .A1(_06586_),
    .S(_06626_),
    .X(_06632_));
 sky130_fd_sc_hd__clkbuf_1 _12308_ (.A(_06632_),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _12309_ (.A0(\cpuregs.regs[25][26] ),
    .A1(_06588_),
    .S(_06626_),
    .X(_06633_));
 sky130_fd_sc_hd__clkbuf_1 _12310_ (.A(_06633_),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _12311_ (.A0(\cpuregs.regs[25][27] ),
    .A1(_06590_),
    .S(_06626_),
    .X(_06634_));
 sky130_fd_sc_hd__clkbuf_1 _12312_ (.A(_06634_),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _12313_ (.A0(\cpuregs.regs[25][28] ),
    .A1(_06592_),
    .S(_06626_),
    .X(_06635_));
 sky130_fd_sc_hd__clkbuf_1 _12314_ (.A(_06635_),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _12315_ (.A0(\cpuregs.regs[25][29] ),
    .A1(_06594_),
    .S(_06626_),
    .X(_06636_));
 sky130_fd_sc_hd__clkbuf_1 _12316_ (.A(_06636_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _12317_ (.A0(\cpuregs.regs[25][30] ),
    .A1(_06596_),
    .S(_06603_),
    .X(_06637_));
 sky130_fd_sc_hd__clkbuf_1 _12318_ (.A(_06637_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _12319_ (.A0(\cpuregs.regs[25][31] ),
    .A1(_06598_),
    .S(_06603_),
    .X(_06638_));
 sky130_fd_sc_hd__clkbuf_1 _12320_ (.A(_06638_),
    .X(_00350_));
 sky130_fd_sc_hd__or2b_2 _12321_ (.A(\cpuregs.waddr[0] ),
    .B_N(\cpuregs.waddr[1] ),
    .X(_06639_));
 sky130_fd_sc_hd__nor2_4 _12322_ (.A(_06639_),
    .B(_06532_),
    .Y(_06640_));
 sky130_fd_sc_hd__clkbuf_8 _12323_ (.A(_06640_),
    .X(_06641_));
 sky130_fd_sc_hd__mux2_1 _12324_ (.A0(\cpuregs.regs[26][0] ),
    .A1(_06531_),
    .S(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__clkbuf_1 _12325_ (.A(_06642_),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _12326_ (.A0(\cpuregs.regs[26][1] ),
    .A1(_06536_),
    .S(_06641_),
    .X(_06643_));
 sky130_fd_sc_hd__clkbuf_1 _12327_ (.A(_06643_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _12328_ (.A0(\cpuregs.regs[26][2] ),
    .A1(_06538_),
    .S(_06641_),
    .X(_06644_));
 sky130_fd_sc_hd__clkbuf_1 _12329_ (.A(_06644_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _12330_ (.A0(\cpuregs.regs[26][3] ),
    .A1(_06540_),
    .S(_06641_),
    .X(_06645_));
 sky130_fd_sc_hd__clkbuf_1 _12331_ (.A(_06645_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _12332_ (.A0(\cpuregs.regs[26][4] ),
    .A1(_06542_),
    .S(_06641_),
    .X(_06646_));
 sky130_fd_sc_hd__clkbuf_1 _12333_ (.A(_06646_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _12334_ (.A0(\cpuregs.regs[26][5] ),
    .A1(_06544_),
    .S(_06641_),
    .X(_06647_));
 sky130_fd_sc_hd__clkbuf_1 _12335_ (.A(_06647_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _12336_ (.A0(\cpuregs.regs[26][6] ),
    .A1(_06546_),
    .S(_06641_),
    .X(_06648_));
 sky130_fd_sc_hd__clkbuf_1 _12337_ (.A(_06648_),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _12338_ (.A0(\cpuregs.regs[26][7] ),
    .A1(_06548_),
    .S(_06641_),
    .X(_06649_));
 sky130_fd_sc_hd__clkbuf_1 _12339_ (.A(_06649_),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _12340_ (.A0(\cpuregs.regs[26][8] ),
    .A1(_06550_),
    .S(_06641_),
    .X(_06650_));
 sky130_fd_sc_hd__clkbuf_1 _12341_ (.A(_06650_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _12342_ (.A0(\cpuregs.regs[26][9] ),
    .A1(_06552_),
    .S(_06641_),
    .X(_06651_));
 sky130_fd_sc_hd__clkbuf_1 _12343_ (.A(_06651_),
    .X(_00360_));
 sky130_fd_sc_hd__buf_6 _12344_ (.A(_06640_),
    .X(_06652_));
 sky130_fd_sc_hd__mux2_1 _12345_ (.A0(\cpuregs.regs[26][10] ),
    .A1(_06554_),
    .S(_06652_),
    .X(_06653_));
 sky130_fd_sc_hd__clkbuf_1 _12346_ (.A(_06653_),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _12347_ (.A0(\cpuregs.regs[26][11] ),
    .A1(_06557_),
    .S(_06652_),
    .X(_06654_));
 sky130_fd_sc_hd__clkbuf_1 _12348_ (.A(_06654_),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _12349_ (.A0(\cpuregs.regs[26][12] ),
    .A1(_06559_),
    .S(_06652_),
    .X(_06655_));
 sky130_fd_sc_hd__clkbuf_1 _12350_ (.A(_06655_),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _12351_ (.A0(\cpuregs.regs[26][13] ),
    .A1(_06561_),
    .S(_06652_),
    .X(_06656_));
 sky130_fd_sc_hd__clkbuf_1 _12352_ (.A(_06656_),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _12353_ (.A0(\cpuregs.regs[26][14] ),
    .A1(_06563_),
    .S(_06652_),
    .X(_06657_));
 sky130_fd_sc_hd__clkbuf_1 _12354_ (.A(_06657_),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _12355_ (.A0(\cpuregs.regs[26][15] ),
    .A1(_06565_),
    .S(_06652_),
    .X(_06658_));
 sky130_fd_sc_hd__clkbuf_1 _12356_ (.A(_06658_),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _12357_ (.A0(\cpuregs.regs[26][16] ),
    .A1(_06567_),
    .S(_06652_),
    .X(_06659_));
 sky130_fd_sc_hd__clkbuf_1 _12358_ (.A(_06659_),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _12359_ (.A0(\cpuregs.regs[26][17] ),
    .A1(_06569_),
    .S(_06652_),
    .X(_06660_));
 sky130_fd_sc_hd__clkbuf_1 _12360_ (.A(_06660_),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _12361_ (.A0(\cpuregs.regs[26][18] ),
    .A1(_06571_),
    .S(_06652_),
    .X(_06661_));
 sky130_fd_sc_hd__clkbuf_1 _12362_ (.A(_06661_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _12363_ (.A0(\cpuregs.regs[26][19] ),
    .A1(_06573_),
    .S(_06652_),
    .X(_06662_));
 sky130_fd_sc_hd__clkbuf_1 _12364_ (.A(_06662_),
    .X(_00370_));
 sky130_fd_sc_hd__clkbuf_8 _12365_ (.A(_06640_),
    .X(_06663_));
 sky130_fd_sc_hd__mux2_1 _12366_ (.A0(\cpuregs.regs[26][20] ),
    .A1(_06575_),
    .S(_06663_),
    .X(_06664_));
 sky130_fd_sc_hd__clkbuf_1 _12367_ (.A(_06664_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _12368_ (.A0(\cpuregs.regs[26][21] ),
    .A1(_06578_),
    .S(_06663_),
    .X(_06665_));
 sky130_fd_sc_hd__clkbuf_1 _12369_ (.A(_06665_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _12370_ (.A0(\cpuregs.regs[26][22] ),
    .A1(_06580_),
    .S(_06663_),
    .X(_06666_));
 sky130_fd_sc_hd__clkbuf_1 _12371_ (.A(_06666_),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _12372_ (.A0(\cpuregs.regs[26][23] ),
    .A1(_06582_),
    .S(_06663_),
    .X(_06667_));
 sky130_fd_sc_hd__clkbuf_1 _12373_ (.A(_06667_),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _12374_ (.A0(\cpuregs.regs[26][24] ),
    .A1(_06584_),
    .S(_06663_),
    .X(_06668_));
 sky130_fd_sc_hd__clkbuf_1 _12375_ (.A(_06668_),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _12376_ (.A0(\cpuregs.regs[26][25] ),
    .A1(_06586_),
    .S(_06663_),
    .X(_06669_));
 sky130_fd_sc_hd__clkbuf_1 _12377_ (.A(_06669_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _12378_ (.A0(\cpuregs.regs[26][26] ),
    .A1(_06588_),
    .S(_06663_),
    .X(_06670_));
 sky130_fd_sc_hd__clkbuf_1 _12379_ (.A(_06670_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _12380_ (.A0(\cpuregs.regs[26][27] ),
    .A1(_06590_),
    .S(_06663_),
    .X(_06671_));
 sky130_fd_sc_hd__clkbuf_1 _12381_ (.A(_06671_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(\cpuregs.regs[26][28] ),
    .A1(_06592_),
    .S(_06663_),
    .X(_06672_));
 sky130_fd_sc_hd__clkbuf_1 _12383_ (.A(_06672_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(\cpuregs.regs[26][29] ),
    .A1(_06594_),
    .S(_06663_),
    .X(_06673_));
 sky130_fd_sc_hd__clkbuf_1 _12385_ (.A(_06673_),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _12386_ (.A0(\cpuregs.regs[26][30] ),
    .A1(_06596_),
    .S(_06640_),
    .X(_06674_));
 sky130_fd_sc_hd__clkbuf_1 _12387_ (.A(_06674_),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _12388_ (.A0(\cpuregs.regs[26][31] ),
    .A1(_06598_),
    .S(_06640_),
    .X(_06675_));
 sky130_fd_sc_hd__clkbuf_1 _12389_ (.A(_06675_),
    .X(_00382_));
 sky130_fd_sc_hd__nand2_2 _12390_ (.A(\cpuregs.waddr[1] ),
    .B(\cpuregs.waddr[0] ),
    .Y(_06676_));
 sky130_fd_sc_hd__nor2_4 _12391_ (.A(_06676_),
    .B(_06532_),
    .Y(_06677_));
 sky130_fd_sc_hd__clkbuf_8 _12392_ (.A(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__mux2_1 _12393_ (.A0(\cpuregs.regs[27][0] ),
    .A1(_06531_),
    .S(_06678_),
    .X(_06679_));
 sky130_fd_sc_hd__clkbuf_1 _12394_ (.A(_06679_),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _12395_ (.A0(\cpuregs.regs[27][1] ),
    .A1(_06536_),
    .S(_06678_),
    .X(_06680_));
 sky130_fd_sc_hd__clkbuf_1 _12396_ (.A(_06680_),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _12397_ (.A0(\cpuregs.regs[27][2] ),
    .A1(_06538_),
    .S(_06678_),
    .X(_06681_));
 sky130_fd_sc_hd__clkbuf_1 _12398_ (.A(_06681_),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _12399_ (.A0(\cpuregs.regs[27][3] ),
    .A1(_06540_),
    .S(_06678_),
    .X(_06682_));
 sky130_fd_sc_hd__clkbuf_1 _12400_ (.A(_06682_),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _12401_ (.A0(\cpuregs.regs[27][4] ),
    .A1(_06542_),
    .S(_06678_),
    .X(_06683_));
 sky130_fd_sc_hd__clkbuf_1 _12402_ (.A(_06683_),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _12403_ (.A0(\cpuregs.regs[27][5] ),
    .A1(_06544_),
    .S(_06678_),
    .X(_06684_));
 sky130_fd_sc_hd__clkbuf_1 _12404_ (.A(_06684_),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _12405_ (.A0(\cpuregs.regs[27][6] ),
    .A1(_06546_),
    .S(_06678_),
    .X(_06685_));
 sky130_fd_sc_hd__clkbuf_1 _12406_ (.A(_06685_),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _12407_ (.A0(\cpuregs.regs[27][7] ),
    .A1(_06548_),
    .S(_06678_),
    .X(_06686_));
 sky130_fd_sc_hd__clkbuf_1 _12408_ (.A(_06686_),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _12409_ (.A0(\cpuregs.regs[27][8] ),
    .A1(_06550_),
    .S(_06678_),
    .X(_06687_));
 sky130_fd_sc_hd__clkbuf_1 _12410_ (.A(_06687_),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _12411_ (.A0(\cpuregs.regs[27][9] ),
    .A1(_06552_),
    .S(_06678_),
    .X(_06688_));
 sky130_fd_sc_hd__clkbuf_1 _12412_ (.A(_06688_),
    .X(_00392_));
 sky130_fd_sc_hd__clkbuf_8 _12413_ (.A(_06677_),
    .X(_06689_));
 sky130_fd_sc_hd__mux2_1 _12414_ (.A0(\cpuregs.regs[27][10] ),
    .A1(_06554_),
    .S(_06689_),
    .X(_06690_));
 sky130_fd_sc_hd__clkbuf_1 _12415_ (.A(_06690_),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _12416_ (.A0(\cpuregs.regs[27][11] ),
    .A1(_06557_),
    .S(_06689_),
    .X(_06691_));
 sky130_fd_sc_hd__clkbuf_1 _12417_ (.A(_06691_),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _12418_ (.A0(\cpuregs.regs[27][12] ),
    .A1(_06559_),
    .S(_06689_),
    .X(_06692_));
 sky130_fd_sc_hd__clkbuf_1 _12419_ (.A(_06692_),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _12420_ (.A0(\cpuregs.regs[27][13] ),
    .A1(_06561_),
    .S(_06689_),
    .X(_06693_));
 sky130_fd_sc_hd__clkbuf_1 _12421_ (.A(_06693_),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _12422_ (.A0(\cpuregs.regs[27][14] ),
    .A1(_06563_),
    .S(_06689_),
    .X(_06694_));
 sky130_fd_sc_hd__clkbuf_1 _12423_ (.A(_06694_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _12424_ (.A0(\cpuregs.regs[27][15] ),
    .A1(_06565_),
    .S(_06689_),
    .X(_06695_));
 sky130_fd_sc_hd__clkbuf_1 _12425_ (.A(_06695_),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _12426_ (.A0(\cpuregs.regs[27][16] ),
    .A1(_06567_),
    .S(_06689_),
    .X(_06696_));
 sky130_fd_sc_hd__clkbuf_1 _12427_ (.A(_06696_),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _12428_ (.A0(\cpuregs.regs[27][17] ),
    .A1(_06569_),
    .S(_06689_),
    .X(_06697_));
 sky130_fd_sc_hd__clkbuf_1 _12429_ (.A(_06697_),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _12430_ (.A0(\cpuregs.regs[27][18] ),
    .A1(_06571_),
    .S(_06689_),
    .X(_06698_));
 sky130_fd_sc_hd__clkbuf_1 _12431_ (.A(_06698_),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _12432_ (.A0(\cpuregs.regs[27][19] ),
    .A1(_06573_),
    .S(_06689_),
    .X(_06699_));
 sky130_fd_sc_hd__clkbuf_1 _12433_ (.A(_06699_),
    .X(_00402_));
 sky130_fd_sc_hd__clkbuf_8 _12434_ (.A(_06677_),
    .X(_06700_));
 sky130_fd_sc_hd__mux2_1 _12435_ (.A0(\cpuregs.regs[27][20] ),
    .A1(_06575_),
    .S(_06700_),
    .X(_06701_));
 sky130_fd_sc_hd__clkbuf_1 _12436_ (.A(_06701_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _12437_ (.A0(\cpuregs.regs[27][21] ),
    .A1(_06578_),
    .S(_06700_),
    .X(_06702_));
 sky130_fd_sc_hd__clkbuf_1 _12438_ (.A(_06702_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _12439_ (.A0(\cpuregs.regs[27][22] ),
    .A1(_06580_),
    .S(_06700_),
    .X(_06703_));
 sky130_fd_sc_hd__clkbuf_1 _12440_ (.A(_06703_),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _12441_ (.A0(\cpuregs.regs[27][23] ),
    .A1(_06582_),
    .S(_06700_),
    .X(_06704_));
 sky130_fd_sc_hd__clkbuf_1 _12442_ (.A(_06704_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _12443_ (.A0(\cpuregs.regs[27][24] ),
    .A1(_06584_),
    .S(_06700_),
    .X(_06705_));
 sky130_fd_sc_hd__clkbuf_1 _12444_ (.A(_06705_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _12445_ (.A0(\cpuregs.regs[27][25] ),
    .A1(_06586_),
    .S(_06700_),
    .X(_06706_));
 sky130_fd_sc_hd__clkbuf_1 _12446_ (.A(_06706_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _12447_ (.A0(\cpuregs.regs[27][26] ),
    .A1(_06588_),
    .S(_06700_),
    .X(_06707_));
 sky130_fd_sc_hd__clkbuf_1 _12448_ (.A(_06707_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _12449_ (.A0(\cpuregs.regs[27][27] ),
    .A1(_06590_),
    .S(_06700_),
    .X(_06708_));
 sky130_fd_sc_hd__clkbuf_1 _12450_ (.A(_06708_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _12451_ (.A0(\cpuregs.regs[27][28] ),
    .A1(_06592_),
    .S(_06700_),
    .X(_06709_));
 sky130_fd_sc_hd__clkbuf_1 _12452_ (.A(_06709_),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _12453_ (.A0(\cpuregs.regs[27][29] ),
    .A1(_06594_),
    .S(_06700_),
    .X(_06710_));
 sky130_fd_sc_hd__clkbuf_1 _12454_ (.A(_06710_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(\cpuregs.regs[27][30] ),
    .A1(_06596_),
    .S(_06677_),
    .X(_06711_));
 sky130_fd_sc_hd__clkbuf_1 _12456_ (.A(_06711_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _12457_ (.A0(\cpuregs.regs[27][31] ),
    .A1(_06598_),
    .S(_06677_),
    .X(_06712_));
 sky130_fd_sc_hd__clkbuf_1 _12458_ (.A(_06712_),
    .X(_00414_));
 sky130_fd_sc_hd__and3_4 _12459_ (.A(_06081_),
    .B(_06082_),
    .C(_06384_),
    .X(_06713_));
 sky130_fd_sc_hd__nand2_4 _12460_ (.A(_06383_),
    .B(_06713_),
    .Y(_06714_));
 sky130_fd_sc_hd__buf_6 _12461_ (.A(_06714_),
    .X(_06715_));
 sky130_fd_sc_hd__mux2_1 _12462_ (.A0(_06078_),
    .A1(\cpuregs.regs[28][0] ),
    .S(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__clkbuf_1 _12463_ (.A(_06716_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _12464_ (.A0(_06096_),
    .A1(\cpuregs.regs[28][1] ),
    .S(_06715_),
    .X(_06717_));
 sky130_fd_sc_hd__clkbuf_1 _12465_ (.A(_06717_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _12466_ (.A0(_06105_),
    .A1(\cpuregs.regs[28][2] ),
    .S(_06715_),
    .X(_06718_));
 sky130_fd_sc_hd__clkbuf_1 _12467_ (.A(_06718_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _12468_ (.A0(_06114_),
    .A1(\cpuregs.regs[28][3] ),
    .S(_06715_),
    .X(_06719_));
 sky130_fd_sc_hd__clkbuf_1 _12469_ (.A(_06719_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _12470_ (.A0(_06125_),
    .A1(\cpuregs.regs[28][4] ),
    .S(_06715_),
    .X(_06720_));
 sky130_fd_sc_hd__clkbuf_1 _12471_ (.A(_06720_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _12472_ (.A0(_06132_),
    .A1(\cpuregs.regs[28][5] ),
    .S(_06715_),
    .X(_06721_));
 sky130_fd_sc_hd__clkbuf_1 _12473_ (.A(_06721_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _12474_ (.A0(_06141_),
    .A1(\cpuregs.regs[28][6] ),
    .S(_06715_),
    .X(_06722_));
 sky130_fd_sc_hd__clkbuf_1 _12475_ (.A(_06722_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _12476_ (.A0(_06150_),
    .A1(\cpuregs.regs[28][7] ),
    .S(_06715_),
    .X(_06723_));
 sky130_fd_sc_hd__clkbuf_1 _12477_ (.A(_06723_),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _12478_ (.A0(_06157_),
    .A1(\cpuregs.regs[28][8] ),
    .S(_06715_),
    .X(_06724_));
 sky130_fd_sc_hd__clkbuf_1 _12479_ (.A(_06724_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _12480_ (.A0(_06166_),
    .A1(\cpuregs.regs[28][9] ),
    .S(_06715_),
    .X(_06725_));
 sky130_fd_sc_hd__clkbuf_1 _12481_ (.A(_06725_),
    .X(_00424_));
 sky130_fd_sc_hd__buf_6 _12482_ (.A(_06714_),
    .X(_06726_));
 sky130_fd_sc_hd__mux2_1 _12483_ (.A0(_06175_),
    .A1(\cpuregs.regs[28][10] ),
    .S(_06726_),
    .X(_06727_));
 sky130_fd_sc_hd__clkbuf_1 _12484_ (.A(_06727_),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _12485_ (.A0(_06184_),
    .A1(\cpuregs.regs[28][11] ),
    .S(_06726_),
    .X(_06728_));
 sky130_fd_sc_hd__clkbuf_1 _12486_ (.A(_06728_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _12487_ (.A0(_06193_),
    .A1(\cpuregs.regs[28][12] ),
    .S(_06726_),
    .X(_06729_));
 sky130_fd_sc_hd__clkbuf_1 _12488_ (.A(_06729_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _12489_ (.A0(_06201_),
    .A1(\cpuregs.regs[28][13] ),
    .S(_06726_),
    .X(_06730_));
 sky130_fd_sc_hd__clkbuf_1 _12490_ (.A(_06730_),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _12491_ (.A0(_06208_),
    .A1(\cpuregs.regs[28][14] ),
    .S(_06726_),
    .X(_06731_));
 sky130_fd_sc_hd__clkbuf_1 _12492_ (.A(_06731_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _12493_ (.A0(_06216_),
    .A1(\cpuregs.regs[28][15] ),
    .S(_06726_),
    .X(_06732_));
 sky130_fd_sc_hd__clkbuf_1 _12494_ (.A(_06732_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _12495_ (.A0(_06224_),
    .A1(\cpuregs.regs[28][16] ),
    .S(_06726_),
    .X(_06733_));
 sky130_fd_sc_hd__clkbuf_1 _12496_ (.A(_06733_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _12497_ (.A0(_06232_),
    .A1(\cpuregs.regs[28][17] ),
    .S(_06726_),
    .X(_06734_));
 sky130_fd_sc_hd__clkbuf_1 _12498_ (.A(_06734_),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _12499_ (.A0(_06240_),
    .A1(\cpuregs.regs[28][18] ),
    .S(_06726_),
    .X(_06735_));
 sky130_fd_sc_hd__clkbuf_1 _12500_ (.A(_06735_),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _12501_ (.A0(_06248_),
    .A1(\cpuregs.regs[28][19] ),
    .S(_06726_),
    .X(_06736_));
 sky130_fd_sc_hd__clkbuf_1 _12502_ (.A(_06736_),
    .X(_00434_));
 sky130_fd_sc_hd__buf_6 _12503_ (.A(_06714_),
    .X(_06737_));
 sky130_fd_sc_hd__mux2_1 _12504_ (.A0(_06257_),
    .A1(\cpuregs.regs[28][20] ),
    .S(_06737_),
    .X(_06738_));
 sky130_fd_sc_hd__clkbuf_1 _12505_ (.A(_06738_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _12506_ (.A0(_06266_),
    .A1(\cpuregs.regs[28][21] ),
    .S(_06737_),
    .X(_06739_));
 sky130_fd_sc_hd__clkbuf_1 _12507_ (.A(_06739_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _12508_ (.A0(_06274_),
    .A1(\cpuregs.regs[28][22] ),
    .S(_06737_),
    .X(_06740_));
 sky130_fd_sc_hd__clkbuf_1 _12509_ (.A(_06740_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _12510_ (.A0(_06281_),
    .A1(\cpuregs.regs[28][23] ),
    .S(_06737_),
    .X(_06741_));
 sky130_fd_sc_hd__clkbuf_1 _12511_ (.A(_06741_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _12512_ (.A0(_06289_),
    .A1(\cpuregs.regs[28][24] ),
    .S(_06737_),
    .X(_06742_));
 sky130_fd_sc_hd__clkbuf_1 _12513_ (.A(_06742_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _12514_ (.A0(_06297_),
    .A1(\cpuregs.regs[28][25] ),
    .S(_06737_),
    .X(_06743_));
 sky130_fd_sc_hd__clkbuf_1 _12515_ (.A(_06743_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _12516_ (.A0(_06304_),
    .A1(\cpuregs.regs[28][26] ),
    .S(_06737_),
    .X(_06744_));
 sky130_fd_sc_hd__clkbuf_1 _12517_ (.A(_06744_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _12518_ (.A0(_06312_),
    .A1(\cpuregs.regs[28][27] ),
    .S(_06737_),
    .X(_06745_));
 sky130_fd_sc_hd__clkbuf_1 _12519_ (.A(_06745_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _12520_ (.A0(_06320_),
    .A1(\cpuregs.regs[28][28] ),
    .S(_06737_),
    .X(_06746_));
 sky130_fd_sc_hd__clkbuf_1 _12521_ (.A(_06746_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _12522_ (.A0(_06328_),
    .A1(\cpuregs.regs[28][29] ),
    .S(_06737_),
    .X(_06747_));
 sky130_fd_sc_hd__clkbuf_1 _12523_ (.A(_06747_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _12524_ (.A0(_06336_),
    .A1(\cpuregs.regs[28][30] ),
    .S(_06714_),
    .X(_06748_));
 sky130_fd_sc_hd__clkbuf_1 _12525_ (.A(_06748_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _12526_ (.A0(_06343_),
    .A1(\cpuregs.regs[28][31] ),
    .S(_06714_),
    .X(_06749_));
 sky130_fd_sc_hd__clkbuf_1 _12527_ (.A(_06749_),
    .X(_00446_));
 sky130_fd_sc_hd__or4b_4 _12528_ (.A(\cpuregs.waddr[2] ),
    .B(\cpuregs.waddr[4] ),
    .C(\cpuregs.waddr[3] ),
    .D_N(_06083_),
    .X(_06750_));
 sky130_fd_sc_hd__nor2_4 _12529_ (.A(_06639_),
    .B(_06750_),
    .Y(_06751_));
 sky130_fd_sc_hd__buf_6 _12530_ (.A(_06751_),
    .X(_06752_));
 sky130_fd_sc_hd__mux2_1 _12531_ (.A0(\cpuregs.regs[2][0] ),
    .A1(_06531_),
    .S(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__clkbuf_1 _12532_ (.A(_06753_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _12533_ (.A0(\cpuregs.regs[2][1] ),
    .A1(_06536_),
    .S(_06752_),
    .X(_06754_));
 sky130_fd_sc_hd__clkbuf_1 _12534_ (.A(_06754_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _12535_ (.A0(\cpuregs.regs[2][2] ),
    .A1(_06538_),
    .S(_06752_),
    .X(_06755_));
 sky130_fd_sc_hd__clkbuf_1 _12536_ (.A(_06755_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _12537_ (.A0(\cpuregs.regs[2][3] ),
    .A1(_06540_),
    .S(_06752_),
    .X(_06756_));
 sky130_fd_sc_hd__clkbuf_1 _12538_ (.A(_06756_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _12539_ (.A0(\cpuregs.regs[2][4] ),
    .A1(_06542_),
    .S(_06752_),
    .X(_06757_));
 sky130_fd_sc_hd__clkbuf_1 _12540_ (.A(_06757_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(\cpuregs.regs[2][5] ),
    .A1(_06544_),
    .S(_06752_),
    .X(_06758_));
 sky130_fd_sc_hd__clkbuf_1 _12542_ (.A(_06758_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _12543_ (.A0(\cpuregs.regs[2][6] ),
    .A1(_06546_),
    .S(_06752_),
    .X(_06759_));
 sky130_fd_sc_hd__clkbuf_1 _12544_ (.A(_06759_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _12545_ (.A0(\cpuregs.regs[2][7] ),
    .A1(_06548_),
    .S(_06752_),
    .X(_06760_));
 sky130_fd_sc_hd__clkbuf_1 _12546_ (.A(_06760_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _12547_ (.A0(\cpuregs.regs[2][8] ),
    .A1(_06550_),
    .S(_06752_),
    .X(_06761_));
 sky130_fd_sc_hd__clkbuf_1 _12548_ (.A(_06761_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _12549_ (.A0(\cpuregs.regs[2][9] ),
    .A1(_06552_),
    .S(_06752_),
    .X(_06762_));
 sky130_fd_sc_hd__clkbuf_1 _12550_ (.A(_06762_),
    .X(_00456_));
 sky130_fd_sc_hd__clkbuf_8 _12551_ (.A(_06751_),
    .X(_06763_));
 sky130_fd_sc_hd__mux2_1 _12552_ (.A0(\cpuregs.regs[2][10] ),
    .A1(_06554_),
    .S(_06763_),
    .X(_06764_));
 sky130_fd_sc_hd__clkbuf_1 _12553_ (.A(_06764_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _12554_ (.A0(\cpuregs.regs[2][11] ),
    .A1(_06557_),
    .S(_06763_),
    .X(_06765_));
 sky130_fd_sc_hd__clkbuf_1 _12555_ (.A(_06765_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _12556_ (.A0(\cpuregs.regs[2][12] ),
    .A1(_06559_),
    .S(_06763_),
    .X(_06766_));
 sky130_fd_sc_hd__clkbuf_1 _12557_ (.A(_06766_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _12558_ (.A0(\cpuregs.regs[2][13] ),
    .A1(_06561_),
    .S(_06763_),
    .X(_06767_));
 sky130_fd_sc_hd__clkbuf_1 _12559_ (.A(_06767_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _12560_ (.A0(\cpuregs.regs[2][14] ),
    .A1(_06563_),
    .S(_06763_),
    .X(_06768_));
 sky130_fd_sc_hd__clkbuf_1 _12561_ (.A(_06768_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _12562_ (.A0(\cpuregs.regs[2][15] ),
    .A1(_06565_),
    .S(_06763_),
    .X(_06769_));
 sky130_fd_sc_hd__clkbuf_1 _12563_ (.A(_06769_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _12564_ (.A0(\cpuregs.regs[2][16] ),
    .A1(_06567_),
    .S(_06763_),
    .X(_06770_));
 sky130_fd_sc_hd__clkbuf_1 _12565_ (.A(_06770_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _12566_ (.A0(\cpuregs.regs[2][17] ),
    .A1(_06569_),
    .S(_06763_),
    .X(_06771_));
 sky130_fd_sc_hd__clkbuf_1 _12567_ (.A(_06771_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _12568_ (.A0(\cpuregs.regs[2][18] ),
    .A1(_06571_),
    .S(_06763_),
    .X(_06772_));
 sky130_fd_sc_hd__clkbuf_1 _12569_ (.A(_06772_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _12570_ (.A0(\cpuregs.regs[2][19] ),
    .A1(_06573_),
    .S(_06763_),
    .X(_06773_));
 sky130_fd_sc_hd__clkbuf_1 _12571_ (.A(_06773_),
    .X(_00466_));
 sky130_fd_sc_hd__buf_6 _12572_ (.A(_06751_),
    .X(_06774_));
 sky130_fd_sc_hd__mux2_1 _12573_ (.A0(\cpuregs.regs[2][20] ),
    .A1(_06575_),
    .S(_06774_),
    .X(_06775_));
 sky130_fd_sc_hd__clkbuf_1 _12574_ (.A(_06775_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _12575_ (.A0(\cpuregs.regs[2][21] ),
    .A1(_06578_),
    .S(_06774_),
    .X(_06776_));
 sky130_fd_sc_hd__clkbuf_1 _12576_ (.A(_06776_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _12577_ (.A0(\cpuregs.regs[2][22] ),
    .A1(_06580_),
    .S(_06774_),
    .X(_06777_));
 sky130_fd_sc_hd__clkbuf_1 _12578_ (.A(_06777_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _12579_ (.A0(\cpuregs.regs[2][23] ),
    .A1(_06582_),
    .S(_06774_),
    .X(_06778_));
 sky130_fd_sc_hd__clkbuf_1 _12580_ (.A(_06778_),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _12581_ (.A0(\cpuregs.regs[2][24] ),
    .A1(_06584_),
    .S(_06774_),
    .X(_06779_));
 sky130_fd_sc_hd__clkbuf_1 _12582_ (.A(_06779_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _12583_ (.A0(\cpuregs.regs[2][25] ),
    .A1(_06586_),
    .S(_06774_),
    .X(_06780_));
 sky130_fd_sc_hd__clkbuf_1 _12584_ (.A(_06780_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _12585_ (.A0(\cpuregs.regs[2][26] ),
    .A1(_06588_),
    .S(_06774_),
    .X(_06781_));
 sky130_fd_sc_hd__clkbuf_1 _12586_ (.A(_06781_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _12587_ (.A0(\cpuregs.regs[2][27] ),
    .A1(_06590_),
    .S(_06774_),
    .X(_06782_));
 sky130_fd_sc_hd__clkbuf_1 _12588_ (.A(_06782_),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _12589_ (.A0(\cpuregs.regs[2][28] ),
    .A1(_06592_),
    .S(_06774_),
    .X(_06783_));
 sky130_fd_sc_hd__clkbuf_1 _12590_ (.A(_06783_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _12591_ (.A0(\cpuregs.regs[2][29] ),
    .A1(_06594_),
    .S(_06774_),
    .X(_06784_));
 sky130_fd_sc_hd__clkbuf_1 _12592_ (.A(_06784_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _12593_ (.A0(\cpuregs.regs[2][30] ),
    .A1(_06596_),
    .S(_06751_),
    .X(_06785_));
 sky130_fd_sc_hd__clkbuf_1 _12594_ (.A(_06785_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _12595_ (.A0(\cpuregs.regs[2][31] ),
    .A1(_06598_),
    .S(_06751_),
    .X(_06786_));
 sky130_fd_sc_hd__clkbuf_1 _12596_ (.A(_06786_),
    .X(_00478_));
 sky130_fd_sc_hd__nand2_4 _12597_ (.A(_06080_),
    .B(_06713_),
    .Y(_06787_));
 sky130_fd_sc_hd__clkbuf_8 _12598_ (.A(_06787_),
    .X(_06788_));
 sky130_fd_sc_hd__mux2_1 _12599_ (.A0(_06078_),
    .A1(\cpuregs.regs[30][0] ),
    .S(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__clkbuf_1 _12600_ (.A(_06789_),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _12601_ (.A0(_06096_),
    .A1(\cpuregs.regs[30][1] ),
    .S(_06788_),
    .X(_06790_));
 sky130_fd_sc_hd__clkbuf_1 _12602_ (.A(_06790_),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _12603_ (.A0(_06105_),
    .A1(\cpuregs.regs[30][2] ),
    .S(_06788_),
    .X(_06791_));
 sky130_fd_sc_hd__clkbuf_1 _12604_ (.A(_06791_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _12605_ (.A0(_06114_),
    .A1(\cpuregs.regs[30][3] ),
    .S(_06788_),
    .X(_06792_));
 sky130_fd_sc_hd__clkbuf_1 _12606_ (.A(_06792_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _12607_ (.A0(_06125_),
    .A1(\cpuregs.regs[30][4] ),
    .S(_06788_),
    .X(_06793_));
 sky130_fd_sc_hd__clkbuf_1 _12608_ (.A(_06793_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _12609_ (.A0(_06132_),
    .A1(\cpuregs.regs[30][5] ),
    .S(_06788_),
    .X(_06794_));
 sky130_fd_sc_hd__clkbuf_1 _12610_ (.A(_06794_),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _12611_ (.A0(_06141_),
    .A1(\cpuregs.regs[30][6] ),
    .S(_06788_),
    .X(_06795_));
 sky130_fd_sc_hd__clkbuf_1 _12612_ (.A(_06795_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _12613_ (.A0(_06150_),
    .A1(\cpuregs.regs[30][7] ),
    .S(_06788_),
    .X(_06796_));
 sky130_fd_sc_hd__clkbuf_1 _12614_ (.A(_06796_),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _12615_ (.A0(_06157_),
    .A1(\cpuregs.regs[30][8] ),
    .S(_06788_),
    .X(_06797_));
 sky130_fd_sc_hd__clkbuf_1 _12616_ (.A(_06797_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _12617_ (.A0(_06166_),
    .A1(\cpuregs.regs[30][9] ),
    .S(_06788_),
    .X(_06798_));
 sky130_fd_sc_hd__clkbuf_1 _12618_ (.A(_06798_),
    .X(_00488_));
 sky130_fd_sc_hd__buf_6 _12619_ (.A(_06787_),
    .X(_06799_));
 sky130_fd_sc_hd__mux2_1 _12620_ (.A0(_06175_),
    .A1(\cpuregs.regs[30][10] ),
    .S(_06799_),
    .X(_06800_));
 sky130_fd_sc_hd__clkbuf_1 _12621_ (.A(_06800_),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _12622_ (.A0(_06184_),
    .A1(\cpuregs.regs[30][11] ),
    .S(_06799_),
    .X(_06801_));
 sky130_fd_sc_hd__clkbuf_1 _12623_ (.A(_06801_),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _12624_ (.A0(_06193_),
    .A1(\cpuregs.regs[30][12] ),
    .S(_06799_),
    .X(_06802_));
 sky130_fd_sc_hd__clkbuf_1 _12625_ (.A(_06802_),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _12626_ (.A0(_06201_),
    .A1(\cpuregs.regs[30][13] ),
    .S(_06799_),
    .X(_06803_));
 sky130_fd_sc_hd__clkbuf_1 _12627_ (.A(_06803_),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _12628_ (.A0(_06208_),
    .A1(\cpuregs.regs[30][14] ),
    .S(_06799_),
    .X(_06804_));
 sky130_fd_sc_hd__clkbuf_1 _12629_ (.A(_06804_),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _12630_ (.A0(_06216_),
    .A1(\cpuregs.regs[30][15] ),
    .S(_06799_),
    .X(_06805_));
 sky130_fd_sc_hd__clkbuf_1 _12631_ (.A(_06805_),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _12632_ (.A0(_06224_),
    .A1(\cpuregs.regs[30][16] ),
    .S(_06799_),
    .X(_06806_));
 sky130_fd_sc_hd__clkbuf_1 _12633_ (.A(_06806_),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _12634_ (.A0(_06232_),
    .A1(\cpuregs.regs[30][17] ),
    .S(_06799_),
    .X(_06807_));
 sky130_fd_sc_hd__clkbuf_1 _12635_ (.A(_06807_),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _12636_ (.A0(_06240_),
    .A1(\cpuregs.regs[30][18] ),
    .S(_06799_),
    .X(_06808_));
 sky130_fd_sc_hd__clkbuf_1 _12637_ (.A(_06808_),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _12638_ (.A0(_06248_),
    .A1(\cpuregs.regs[30][19] ),
    .S(_06799_),
    .X(_06809_));
 sky130_fd_sc_hd__clkbuf_1 _12639_ (.A(_06809_),
    .X(_00498_));
 sky130_fd_sc_hd__clkbuf_8 _12640_ (.A(_06787_),
    .X(_06810_));
 sky130_fd_sc_hd__mux2_1 _12641_ (.A0(_06257_),
    .A1(\cpuregs.regs[30][20] ),
    .S(_06810_),
    .X(_06811_));
 sky130_fd_sc_hd__clkbuf_1 _12642_ (.A(_06811_),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _12643_ (.A0(_06266_),
    .A1(\cpuregs.regs[30][21] ),
    .S(_06810_),
    .X(_06812_));
 sky130_fd_sc_hd__clkbuf_1 _12644_ (.A(_06812_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _12645_ (.A0(_06274_),
    .A1(\cpuregs.regs[30][22] ),
    .S(_06810_),
    .X(_06813_));
 sky130_fd_sc_hd__clkbuf_1 _12646_ (.A(_06813_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _12647_ (.A0(_06281_),
    .A1(\cpuregs.regs[30][23] ),
    .S(_06810_),
    .X(_06814_));
 sky130_fd_sc_hd__clkbuf_1 _12648_ (.A(_06814_),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _12649_ (.A0(_06289_),
    .A1(\cpuregs.regs[30][24] ),
    .S(_06810_),
    .X(_06815_));
 sky130_fd_sc_hd__clkbuf_1 _12650_ (.A(_06815_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _12651_ (.A0(_06297_),
    .A1(\cpuregs.regs[30][25] ),
    .S(_06810_),
    .X(_06816_));
 sky130_fd_sc_hd__clkbuf_1 _12652_ (.A(_06816_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _12653_ (.A0(_06304_),
    .A1(\cpuregs.regs[30][26] ),
    .S(_06810_),
    .X(_06817_));
 sky130_fd_sc_hd__clkbuf_1 _12654_ (.A(_06817_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _12655_ (.A0(_06312_),
    .A1(\cpuregs.regs[30][27] ),
    .S(_06810_),
    .X(_06818_));
 sky130_fd_sc_hd__clkbuf_1 _12656_ (.A(_06818_),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _12657_ (.A0(_06320_),
    .A1(\cpuregs.regs[30][28] ),
    .S(_06810_),
    .X(_06819_));
 sky130_fd_sc_hd__clkbuf_1 _12658_ (.A(_06819_),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _12659_ (.A0(_06328_),
    .A1(\cpuregs.regs[30][29] ),
    .S(_06810_),
    .X(_06820_));
 sky130_fd_sc_hd__clkbuf_1 _12660_ (.A(_06820_),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _12661_ (.A0(_06336_),
    .A1(\cpuregs.regs[30][30] ),
    .S(_06787_),
    .X(_06821_));
 sky130_fd_sc_hd__clkbuf_1 _12662_ (.A(_06821_),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _12663_ (.A0(_06343_),
    .A1(\cpuregs.regs[30][31] ),
    .S(_06787_),
    .X(_06822_));
 sky130_fd_sc_hd__clkbuf_1 _12664_ (.A(_06822_),
    .X(_00510_));
 sky130_fd_sc_hd__and3b_2 _12665_ (.A_N(_06081_),
    .B(_06082_),
    .C(_06384_),
    .X(_06823_));
 sky130_fd_sc_hd__nand2_2 _12666_ (.A(_06383_),
    .B(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__clkbuf_8 _12667_ (.A(_06824_),
    .X(_06825_));
 sky130_fd_sc_hd__mux2_1 _12668_ (.A0(_06078_),
    .A1(\cpuregs.regs[12][0] ),
    .S(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__clkbuf_1 _12669_ (.A(_06826_),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _12670_ (.A0(_06096_),
    .A1(\cpuregs.regs[12][1] ),
    .S(_06825_),
    .X(_06827_));
 sky130_fd_sc_hd__clkbuf_1 _12671_ (.A(_06827_),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _12672_ (.A0(_06105_),
    .A1(\cpuregs.regs[12][2] ),
    .S(_06825_),
    .X(_06828_));
 sky130_fd_sc_hd__clkbuf_1 _12673_ (.A(_06828_),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _12674_ (.A0(_06114_),
    .A1(\cpuregs.regs[12][3] ),
    .S(_06825_),
    .X(_06829_));
 sky130_fd_sc_hd__clkbuf_1 _12675_ (.A(_06829_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _12676_ (.A0(_06125_),
    .A1(\cpuregs.regs[12][4] ),
    .S(_06825_),
    .X(_06830_));
 sky130_fd_sc_hd__clkbuf_1 _12677_ (.A(_06830_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _12678_ (.A0(_06132_),
    .A1(\cpuregs.regs[12][5] ),
    .S(_06825_),
    .X(_06831_));
 sky130_fd_sc_hd__clkbuf_1 _12679_ (.A(_06831_),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _12680_ (.A0(_06141_),
    .A1(\cpuregs.regs[12][6] ),
    .S(_06825_),
    .X(_06832_));
 sky130_fd_sc_hd__clkbuf_1 _12681_ (.A(_06832_),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _12682_ (.A0(_06150_),
    .A1(\cpuregs.regs[12][7] ),
    .S(_06825_),
    .X(_06833_));
 sky130_fd_sc_hd__clkbuf_1 _12683_ (.A(_06833_),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _12684_ (.A0(_06157_),
    .A1(\cpuregs.regs[12][8] ),
    .S(_06825_),
    .X(_06834_));
 sky130_fd_sc_hd__clkbuf_1 _12685_ (.A(_06834_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _12686_ (.A0(_06166_),
    .A1(\cpuregs.regs[12][9] ),
    .S(_06825_),
    .X(_06835_));
 sky130_fd_sc_hd__clkbuf_1 _12687_ (.A(_06835_),
    .X(_00520_));
 sky130_fd_sc_hd__buf_6 _12688_ (.A(_06824_),
    .X(_06836_));
 sky130_fd_sc_hd__mux2_1 _12689_ (.A0(_06175_),
    .A1(\cpuregs.regs[12][10] ),
    .S(_06836_),
    .X(_06837_));
 sky130_fd_sc_hd__clkbuf_1 _12690_ (.A(_06837_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _12691_ (.A0(_06184_),
    .A1(\cpuregs.regs[12][11] ),
    .S(_06836_),
    .X(_06838_));
 sky130_fd_sc_hd__clkbuf_1 _12692_ (.A(_06838_),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _12693_ (.A0(_06193_),
    .A1(\cpuregs.regs[12][12] ),
    .S(_06836_),
    .X(_06839_));
 sky130_fd_sc_hd__clkbuf_1 _12694_ (.A(_06839_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _12695_ (.A0(_06201_),
    .A1(\cpuregs.regs[12][13] ),
    .S(_06836_),
    .X(_06840_));
 sky130_fd_sc_hd__clkbuf_1 _12696_ (.A(_06840_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _12697_ (.A0(_06208_),
    .A1(\cpuregs.regs[12][14] ),
    .S(_06836_),
    .X(_06841_));
 sky130_fd_sc_hd__clkbuf_1 _12698_ (.A(_06841_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _12699_ (.A0(_06216_),
    .A1(\cpuregs.regs[12][15] ),
    .S(_06836_),
    .X(_06842_));
 sky130_fd_sc_hd__clkbuf_1 _12700_ (.A(_06842_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _12701_ (.A0(_06224_),
    .A1(\cpuregs.regs[12][16] ),
    .S(_06836_),
    .X(_06843_));
 sky130_fd_sc_hd__clkbuf_1 _12702_ (.A(_06843_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _12703_ (.A0(_06232_),
    .A1(\cpuregs.regs[12][17] ),
    .S(_06836_),
    .X(_06844_));
 sky130_fd_sc_hd__clkbuf_1 _12704_ (.A(_06844_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _12705_ (.A0(_06240_),
    .A1(\cpuregs.regs[12][18] ),
    .S(_06836_),
    .X(_06845_));
 sky130_fd_sc_hd__clkbuf_1 _12706_ (.A(_06845_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _12707_ (.A0(_06248_),
    .A1(\cpuregs.regs[12][19] ),
    .S(_06836_),
    .X(_06846_));
 sky130_fd_sc_hd__clkbuf_1 _12708_ (.A(_06846_),
    .X(_00530_));
 sky130_fd_sc_hd__clkbuf_8 _12709_ (.A(_06824_),
    .X(_06847_));
 sky130_fd_sc_hd__mux2_1 _12710_ (.A0(_06257_),
    .A1(\cpuregs.regs[12][20] ),
    .S(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__clkbuf_1 _12711_ (.A(_06848_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _12712_ (.A0(_06266_),
    .A1(\cpuregs.regs[12][21] ),
    .S(_06847_),
    .X(_06849_));
 sky130_fd_sc_hd__clkbuf_1 _12713_ (.A(_06849_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _12714_ (.A0(_06274_),
    .A1(\cpuregs.regs[12][22] ),
    .S(_06847_),
    .X(_06850_));
 sky130_fd_sc_hd__clkbuf_1 _12715_ (.A(_06850_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _12716_ (.A0(_06281_),
    .A1(\cpuregs.regs[12][23] ),
    .S(_06847_),
    .X(_06851_));
 sky130_fd_sc_hd__clkbuf_1 _12717_ (.A(_06851_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _12718_ (.A0(_06289_),
    .A1(\cpuregs.regs[12][24] ),
    .S(_06847_),
    .X(_06852_));
 sky130_fd_sc_hd__clkbuf_1 _12719_ (.A(_06852_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _12720_ (.A0(_06297_),
    .A1(\cpuregs.regs[12][25] ),
    .S(_06847_),
    .X(_06853_));
 sky130_fd_sc_hd__clkbuf_1 _12721_ (.A(_06853_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _12722_ (.A0(_06304_),
    .A1(\cpuregs.regs[12][26] ),
    .S(_06847_),
    .X(_06854_));
 sky130_fd_sc_hd__clkbuf_1 _12723_ (.A(_06854_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _12724_ (.A0(_06312_),
    .A1(\cpuregs.regs[12][27] ),
    .S(_06847_),
    .X(_06855_));
 sky130_fd_sc_hd__clkbuf_1 _12725_ (.A(_06855_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _12726_ (.A0(_06320_),
    .A1(\cpuregs.regs[12][28] ),
    .S(_06847_),
    .X(_06856_));
 sky130_fd_sc_hd__clkbuf_1 _12727_ (.A(_06856_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _12728_ (.A0(_06328_),
    .A1(\cpuregs.regs[12][29] ),
    .S(_06847_),
    .X(_06857_));
 sky130_fd_sc_hd__clkbuf_1 _12729_ (.A(_06857_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _12730_ (.A0(_06336_),
    .A1(\cpuregs.regs[12][30] ),
    .S(_06824_),
    .X(_06858_));
 sky130_fd_sc_hd__clkbuf_1 _12731_ (.A(_06858_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _12732_ (.A0(_06343_),
    .A1(\cpuregs.regs[12][31] ),
    .S(_06824_),
    .X(_06859_));
 sky130_fd_sc_hd__clkbuf_1 _12733_ (.A(_06859_),
    .X(_00542_));
 sky130_fd_sc_hd__nand2_4 _12734_ (.A(_03298_),
    .B(_03277_),
    .Y(_06860_));
 sky130_fd_sc_hd__nor2_2 _12735_ (.A(\cpu_state[3] ),
    .B(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__a31oi_4 _12736_ (.A1(_03309_),
    .A2(_03384_),
    .A3(_06053_),
    .B1(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__clkbuf_4 _12737_ (.A(_03364_),
    .X(_06863_));
 sky130_fd_sc_hd__nor2_1 _12738_ (.A(_06186_),
    .B(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__a21o_1 _12739_ (.A1(\decoded_rd[0] ),
    .A2(_06863_),
    .B1(_06864_),
    .X(_06865_));
 sky130_fd_sc_hd__a22o_1 _12740_ (.A1(\cpuregs.waddr[0] ),
    .A2(_06862_),
    .B1(_06865_),
    .B2(_06861_),
    .X(_00543_));
 sky130_fd_sc_hd__a21o_1 _12741_ (.A1(\decoded_rd[1] ),
    .A2(_06863_),
    .B1(_06864_),
    .X(_06866_));
 sky130_fd_sc_hd__a22o_1 _12742_ (.A1(\cpuregs.waddr[1] ),
    .A2(_06862_),
    .B1(_06866_),
    .B2(_06861_),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _12743_ (.A0(_06186_),
    .A1(\decoded_rd[2] ),
    .S(_06863_),
    .X(_06867_));
 sky130_fd_sc_hd__a22o_1 _12744_ (.A1(\cpuregs.waddr[2] ),
    .A2(_06862_),
    .B1(_06867_),
    .B2(_06861_),
    .X(_00545_));
 sky130_fd_sc_hd__and4bb_4 _12745_ (.A_N(\cpuregs.waddr[2] ),
    .B_N(_06081_),
    .C(_06082_),
    .D(_06601_),
    .X(_06868_));
 sky130_fd_sc_hd__buf_6 _12746_ (.A(_06868_),
    .X(_06869_));
 sky130_fd_sc_hd__mux2_1 _12747_ (.A0(\cpuregs.regs[9][0] ),
    .A1(_06531_),
    .S(_06869_),
    .X(_06870_));
 sky130_fd_sc_hd__clkbuf_1 _12748_ (.A(_06870_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _12749_ (.A0(\cpuregs.regs[9][1] ),
    .A1(_06536_),
    .S(_06869_),
    .X(_06871_));
 sky130_fd_sc_hd__clkbuf_1 _12750_ (.A(_06871_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _12751_ (.A0(\cpuregs.regs[9][2] ),
    .A1(_06538_),
    .S(_06869_),
    .X(_06872_));
 sky130_fd_sc_hd__clkbuf_1 _12752_ (.A(_06872_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _12753_ (.A0(\cpuregs.regs[9][3] ),
    .A1(_06540_),
    .S(_06869_),
    .X(_06873_));
 sky130_fd_sc_hd__clkbuf_1 _12754_ (.A(_06873_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _12755_ (.A0(\cpuregs.regs[9][4] ),
    .A1(_06542_),
    .S(_06869_),
    .X(_06874_));
 sky130_fd_sc_hd__clkbuf_1 _12756_ (.A(_06874_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _12757_ (.A0(\cpuregs.regs[9][5] ),
    .A1(_06544_),
    .S(_06869_),
    .X(_06875_));
 sky130_fd_sc_hd__clkbuf_1 _12758_ (.A(_06875_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _12759_ (.A0(\cpuregs.regs[9][6] ),
    .A1(_06546_),
    .S(_06869_),
    .X(_06876_));
 sky130_fd_sc_hd__clkbuf_1 _12760_ (.A(_06876_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _12761_ (.A0(\cpuregs.regs[9][7] ),
    .A1(_06548_),
    .S(_06869_),
    .X(_06877_));
 sky130_fd_sc_hd__clkbuf_1 _12762_ (.A(_06877_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _12763_ (.A0(\cpuregs.regs[9][8] ),
    .A1(_06550_),
    .S(_06869_),
    .X(_06878_));
 sky130_fd_sc_hd__clkbuf_1 _12764_ (.A(_06878_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _12765_ (.A0(\cpuregs.regs[9][9] ),
    .A1(_06552_),
    .S(_06869_),
    .X(_06879_));
 sky130_fd_sc_hd__clkbuf_1 _12766_ (.A(_06879_),
    .X(_00555_));
 sky130_fd_sc_hd__clkbuf_8 _12767_ (.A(_06868_),
    .X(_06880_));
 sky130_fd_sc_hd__mux2_1 _12768_ (.A0(\cpuregs.regs[9][10] ),
    .A1(_06554_),
    .S(_06880_),
    .X(_06881_));
 sky130_fd_sc_hd__clkbuf_1 _12769_ (.A(_06881_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _12770_ (.A0(\cpuregs.regs[9][11] ),
    .A1(_06557_),
    .S(_06880_),
    .X(_06882_));
 sky130_fd_sc_hd__clkbuf_1 _12771_ (.A(_06882_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _12772_ (.A0(\cpuregs.regs[9][12] ),
    .A1(_06559_),
    .S(_06880_),
    .X(_06883_));
 sky130_fd_sc_hd__clkbuf_1 _12773_ (.A(_06883_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _12774_ (.A0(\cpuregs.regs[9][13] ),
    .A1(_06561_),
    .S(_06880_),
    .X(_06884_));
 sky130_fd_sc_hd__clkbuf_1 _12775_ (.A(_06884_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _12776_ (.A0(\cpuregs.regs[9][14] ),
    .A1(_06563_),
    .S(_06880_),
    .X(_06885_));
 sky130_fd_sc_hd__clkbuf_1 _12777_ (.A(_06885_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _12778_ (.A0(\cpuregs.regs[9][15] ),
    .A1(_06565_),
    .S(_06880_),
    .X(_06886_));
 sky130_fd_sc_hd__clkbuf_1 _12779_ (.A(_06886_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _12780_ (.A0(\cpuregs.regs[9][16] ),
    .A1(_06567_),
    .S(_06880_),
    .X(_06887_));
 sky130_fd_sc_hd__clkbuf_1 _12781_ (.A(_06887_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _12782_ (.A0(\cpuregs.regs[9][17] ),
    .A1(_06569_),
    .S(_06880_),
    .X(_06888_));
 sky130_fd_sc_hd__clkbuf_1 _12783_ (.A(_06888_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _12784_ (.A0(\cpuregs.regs[9][18] ),
    .A1(_06571_),
    .S(_06880_),
    .X(_06889_));
 sky130_fd_sc_hd__clkbuf_1 _12785_ (.A(_06889_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _12786_ (.A0(\cpuregs.regs[9][19] ),
    .A1(_06573_),
    .S(_06880_),
    .X(_06890_));
 sky130_fd_sc_hd__clkbuf_1 _12787_ (.A(_06890_),
    .X(_00565_));
 sky130_fd_sc_hd__clkbuf_8 _12788_ (.A(_06868_),
    .X(_06891_));
 sky130_fd_sc_hd__mux2_1 _12789_ (.A0(\cpuregs.regs[9][20] ),
    .A1(_06575_),
    .S(_06891_),
    .X(_06892_));
 sky130_fd_sc_hd__clkbuf_1 _12790_ (.A(_06892_),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _12791_ (.A0(\cpuregs.regs[9][21] ),
    .A1(_06578_),
    .S(_06891_),
    .X(_06893_));
 sky130_fd_sc_hd__clkbuf_1 _12792_ (.A(_06893_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _12793_ (.A0(\cpuregs.regs[9][22] ),
    .A1(_06580_),
    .S(_06891_),
    .X(_06894_));
 sky130_fd_sc_hd__clkbuf_1 _12794_ (.A(_06894_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _12795_ (.A0(\cpuregs.regs[9][23] ),
    .A1(_06582_),
    .S(_06891_),
    .X(_06895_));
 sky130_fd_sc_hd__clkbuf_1 _12796_ (.A(_06895_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _12797_ (.A0(\cpuregs.regs[9][24] ),
    .A1(_06584_),
    .S(_06891_),
    .X(_06896_));
 sky130_fd_sc_hd__clkbuf_1 _12798_ (.A(_06896_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _12799_ (.A0(\cpuregs.regs[9][25] ),
    .A1(_06586_),
    .S(_06891_),
    .X(_06897_));
 sky130_fd_sc_hd__clkbuf_1 _12800_ (.A(_06897_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _12801_ (.A0(\cpuregs.regs[9][26] ),
    .A1(_06588_),
    .S(_06891_),
    .X(_06898_));
 sky130_fd_sc_hd__clkbuf_1 _12802_ (.A(_06898_),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _12803_ (.A0(\cpuregs.regs[9][27] ),
    .A1(_06590_),
    .S(_06891_),
    .X(_06899_));
 sky130_fd_sc_hd__clkbuf_1 _12804_ (.A(_06899_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _12805_ (.A0(\cpuregs.regs[9][28] ),
    .A1(_06592_),
    .S(_06891_),
    .X(_06900_));
 sky130_fd_sc_hd__clkbuf_1 _12806_ (.A(_06900_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _12807_ (.A0(\cpuregs.regs[9][29] ),
    .A1(_06594_),
    .S(_06891_),
    .X(_06901_));
 sky130_fd_sc_hd__clkbuf_1 _12808_ (.A(_06901_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _12809_ (.A0(\cpuregs.regs[9][30] ),
    .A1(_06596_),
    .S(_06868_),
    .X(_06902_));
 sky130_fd_sc_hd__clkbuf_1 _12810_ (.A(_06902_),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _12811_ (.A0(\cpuregs.regs[9][31] ),
    .A1(_06598_),
    .S(_06868_),
    .X(_06903_));
 sky130_fd_sc_hd__clkbuf_1 _12812_ (.A(_06903_),
    .X(_00577_));
 sky130_fd_sc_hd__and4bb_4 _12813_ (.A_N(_06081_),
    .B_N(_06082_),
    .C(_06083_),
    .D(\cpuregs.waddr[2] ),
    .X(_06904_));
 sky130_fd_sc_hd__nand2_4 _12814_ (.A(_06080_),
    .B(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__buf_6 _12815_ (.A(_06905_),
    .X(_06906_));
 sky130_fd_sc_hd__mux2_1 _12816_ (.A0(_06078_),
    .A1(\cpuregs.regs[6][0] ),
    .S(_06906_),
    .X(_06907_));
 sky130_fd_sc_hd__clkbuf_1 _12817_ (.A(_06907_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _12818_ (.A0(_06096_),
    .A1(\cpuregs.regs[6][1] ),
    .S(_06906_),
    .X(_06908_));
 sky130_fd_sc_hd__clkbuf_1 _12819_ (.A(_06908_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _12820_ (.A0(_06105_),
    .A1(\cpuregs.regs[6][2] ),
    .S(_06906_),
    .X(_06909_));
 sky130_fd_sc_hd__clkbuf_1 _12821_ (.A(_06909_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _12822_ (.A0(_06114_),
    .A1(\cpuregs.regs[6][3] ),
    .S(_06906_),
    .X(_06910_));
 sky130_fd_sc_hd__clkbuf_1 _12823_ (.A(_06910_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _12824_ (.A0(_06125_),
    .A1(\cpuregs.regs[6][4] ),
    .S(_06906_),
    .X(_06911_));
 sky130_fd_sc_hd__clkbuf_1 _12825_ (.A(_06911_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _12826_ (.A0(_06132_),
    .A1(\cpuregs.regs[6][5] ),
    .S(_06906_),
    .X(_06912_));
 sky130_fd_sc_hd__clkbuf_1 _12827_ (.A(_06912_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _12828_ (.A0(_06141_),
    .A1(\cpuregs.regs[6][6] ),
    .S(_06906_),
    .X(_06913_));
 sky130_fd_sc_hd__clkbuf_1 _12829_ (.A(_06913_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _12830_ (.A0(_06150_),
    .A1(\cpuregs.regs[6][7] ),
    .S(_06906_),
    .X(_06914_));
 sky130_fd_sc_hd__clkbuf_1 _12831_ (.A(_06914_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _12832_ (.A0(_06157_),
    .A1(\cpuregs.regs[6][8] ),
    .S(_06906_),
    .X(_06915_));
 sky130_fd_sc_hd__clkbuf_1 _12833_ (.A(_06915_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _12834_ (.A0(_06166_),
    .A1(\cpuregs.regs[6][9] ),
    .S(_06906_),
    .X(_06916_));
 sky130_fd_sc_hd__clkbuf_1 _12835_ (.A(_06916_),
    .X(_00587_));
 sky130_fd_sc_hd__clkbuf_8 _12836_ (.A(_06905_),
    .X(_06917_));
 sky130_fd_sc_hd__mux2_1 _12837_ (.A0(_06175_),
    .A1(\cpuregs.regs[6][10] ),
    .S(_06917_),
    .X(_06918_));
 sky130_fd_sc_hd__clkbuf_1 _12838_ (.A(_06918_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _12839_ (.A0(_06184_),
    .A1(\cpuregs.regs[6][11] ),
    .S(_06917_),
    .X(_06919_));
 sky130_fd_sc_hd__clkbuf_1 _12840_ (.A(_06919_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _12841_ (.A0(_06193_),
    .A1(\cpuregs.regs[6][12] ),
    .S(_06917_),
    .X(_06920_));
 sky130_fd_sc_hd__clkbuf_1 _12842_ (.A(_06920_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _12843_ (.A0(_06201_),
    .A1(\cpuregs.regs[6][13] ),
    .S(_06917_),
    .X(_06921_));
 sky130_fd_sc_hd__clkbuf_1 _12844_ (.A(_06921_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _12845_ (.A0(_06208_),
    .A1(\cpuregs.regs[6][14] ),
    .S(_06917_),
    .X(_06922_));
 sky130_fd_sc_hd__clkbuf_1 _12846_ (.A(_06922_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _12847_ (.A0(_06216_),
    .A1(\cpuregs.regs[6][15] ),
    .S(_06917_),
    .X(_06923_));
 sky130_fd_sc_hd__clkbuf_1 _12848_ (.A(_06923_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _12849_ (.A0(_06224_),
    .A1(\cpuregs.regs[6][16] ),
    .S(_06917_),
    .X(_06924_));
 sky130_fd_sc_hd__clkbuf_1 _12850_ (.A(_06924_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _12851_ (.A0(_06232_),
    .A1(\cpuregs.regs[6][17] ),
    .S(_06917_),
    .X(_06925_));
 sky130_fd_sc_hd__clkbuf_1 _12852_ (.A(_06925_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _12853_ (.A0(_06240_),
    .A1(\cpuregs.regs[6][18] ),
    .S(_06917_),
    .X(_06926_));
 sky130_fd_sc_hd__clkbuf_1 _12854_ (.A(_06926_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _12855_ (.A0(_06248_),
    .A1(\cpuregs.regs[6][19] ),
    .S(_06917_),
    .X(_06927_));
 sky130_fd_sc_hd__clkbuf_1 _12856_ (.A(_06927_),
    .X(_00597_));
 sky130_fd_sc_hd__clkbuf_8 _12857_ (.A(_06905_),
    .X(_06928_));
 sky130_fd_sc_hd__mux2_1 _12858_ (.A0(_06257_),
    .A1(\cpuregs.regs[6][20] ),
    .S(_06928_),
    .X(_06929_));
 sky130_fd_sc_hd__clkbuf_1 _12859_ (.A(_06929_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _12860_ (.A0(_06266_),
    .A1(\cpuregs.regs[6][21] ),
    .S(_06928_),
    .X(_06930_));
 sky130_fd_sc_hd__clkbuf_1 _12861_ (.A(_06930_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _12862_ (.A0(_06274_),
    .A1(\cpuregs.regs[6][22] ),
    .S(_06928_),
    .X(_06931_));
 sky130_fd_sc_hd__clkbuf_1 _12863_ (.A(_06931_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _12864_ (.A0(_06281_),
    .A1(\cpuregs.regs[6][23] ),
    .S(_06928_),
    .X(_06932_));
 sky130_fd_sc_hd__clkbuf_1 _12865_ (.A(_06932_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _12866_ (.A0(_06289_),
    .A1(\cpuregs.regs[6][24] ),
    .S(_06928_),
    .X(_06933_));
 sky130_fd_sc_hd__clkbuf_1 _12867_ (.A(_06933_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _12868_ (.A0(_06297_),
    .A1(\cpuregs.regs[6][25] ),
    .S(_06928_),
    .X(_06934_));
 sky130_fd_sc_hd__clkbuf_1 _12869_ (.A(_06934_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _12870_ (.A0(_06304_),
    .A1(\cpuregs.regs[6][26] ),
    .S(_06928_),
    .X(_06935_));
 sky130_fd_sc_hd__clkbuf_1 _12871_ (.A(_06935_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _12872_ (.A0(_06312_),
    .A1(\cpuregs.regs[6][27] ),
    .S(_06928_),
    .X(_06936_));
 sky130_fd_sc_hd__clkbuf_1 _12873_ (.A(_06936_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _12874_ (.A0(_06320_),
    .A1(\cpuregs.regs[6][28] ),
    .S(_06928_),
    .X(_06937_));
 sky130_fd_sc_hd__clkbuf_1 _12875_ (.A(_06937_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _12876_ (.A0(_06328_),
    .A1(\cpuregs.regs[6][29] ),
    .S(_06928_),
    .X(_06938_));
 sky130_fd_sc_hd__clkbuf_1 _12877_ (.A(_06938_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _12878_ (.A0(_06336_),
    .A1(\cpuregs.regs[6][30] ),
    .S(_06905_),
    .X(_06939_));
 sky130_fd_sc_hd__clkbuf_1 _12879_ (.A(_06939_),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _12880_ (.A0(_06343_),
    .A1(\cpuregs.regs[6][31] ),
    .S(_06905_),
    .X(_06940_));
 sky130_fd_sc_hd__clkbuf_1 _12881_ (.A(_06940_),
    .X(_00609_));
 sky130_fd_sc_hd__buf_2 _12882_ (.A(_06077_),
    .X(_06941_));
 sky130_fd_sc_hd__nand2_4 _12883_ (.A(_06346_),
    .B(_06713_),
    .Y(_06942_));
 sky130_fd_sc_hd__buf_6 _12884_ (.A(_06942_),
    .X(_06943_));
 sky130_fd_sc_hd__mux2_1 _12885_ (.A0(_06941_),
    .A1(\cpuregs.regs[31][0] ),
    .S(_06943_),
    .X(_06944_));
 sky130_fd_sc_hd__clkbuf_1 _12886_ (.A(_06944_),
    .X(_00610_));
 sky130_fd_sc_hd__buf_2 _12887_ (.A(_06095_),
    .X(_06945_));
 sky130_fd_sc_hd__mux2_1 _12888_ (.A0(_06945_),
    .A1(\cpuregs.regs[31][1] ),
    .S(_06943_),
    .X(_06946_));
 sky130_fd_sc_hd__clkbuf_1 _12889_ (.A(_06946_),
    .X(_00611_));
 sky130_fd_sc_hd__buf_2 _12890_ (.A(_06104_),
    .X(_06947_));
 sky130_fd_sc_hd__mux2_1 _12891_ (.A0(_06947_),
    .A1(\cpuregs.regs[31][2] ),
    .S(_06943_),
    .X(_06948_));
 sky130_fd_sc_hd__clkbuf_1 _12892_ (.A(_06948_),
    .X(_00612_));
 sky130_fd_sc_hd__clkbuf_4 _12893_ (.A(_06113_),
    .X(_06949_));
 sky130_fd_sc_hd__mux2_1 _12894_ (.A0(_06949_),
    .A1(\cpuregs.regs[31][3] ),
    .S(_06943_),
    .X(_06950_));
 sky130_fd_sc_hd__clkbuf_1 _12895_ (.A(_06950_),
    .X(_00613_));
 sky130_fd_sc_hd__buf_2 _12896_ (.A(_06124_),
    .X(_06951_));
 sky130_fd_sc_hd__mux2_1 _12897_ (.A0(_06951_),
    .A1(\cpuregs.regs[31][4] ),
    .S(_06943_),
    .X(_06952_));
 sky130_fd_sc_hd__clkbuf_1 _12898_ (.A(_06952_),
    .X(_00614_));
 sky130_fd_sc_hd__buf_2 _12899_ (.A(_06131_),
    .X(_06953_));
 sky130_fd_sc_hd__mux2_1 _12900_ (.A0(_06953_),
    .A1(\cpuregs.regs[31][5] ),
    .S(_06943_),
    .X(_06954_));
 sky130_fd_sc_hd__clkbuf_1 _12901_ (.A(_06954_),
    .X(_00615_));
 sky130_fd_sc_hd__buf_2 _12902_ (.A(_06140_),
    .X(_06955_));
 sky130_fd_sc_hd__mux2_1 _12903_ (.A0(_06955_),
    .A1(\cpuregs.regs[31][6] ),
    .S(_06943_),
    .X(_06956_));
 sky130_fd_sc_hd__clkbuf_1 _12904_ (.A(_06956_),
    .X(_00616_));
 sky130_fd_sc_hd__buf_2 _12905_ (.A(_06149_),
    .X(_06957_));
 sky130_fd_sc_hd__mux2_1 _12906_ (.A0(_06957_),
    .A1(\cpuregs.regs[31][7] ),
    .S(_06943_),
    .X(_06958_));
 sky130_fd_sc_hd__clkbuf_1 _12907_ (.A(_06958_),
    .X(_00617_));
 sky130_fd_sc_hd__buf_2 _12908_ (.A(_06156_),
    .X(_06959_));
 sky130_fd_sc_hd__mux2_1 _12909_ (.A0(_06959_),
    .A1(\cpuregs.regs[31][8] ),
    .S(_06943_),
    .X(_06960_));
 sky130_fd_sc_hd__clkbuf_1 _12910_ (.A(_06960_),
    .X(_00618_));
 sky130_fd_sc_hd__buf_2 _12911_ (.A(_06165_),
    .X(_06961_));
 sky130_fd_sc_hd__mux2_1 _12912_ (.A0(_06961_),
    .A1(\cpuregs.regs[31][9] ),
    .S(_06943_),
    .X(_06962_));
 sky130_fd_sc_hd__clkbuf_1 _12913_ (.A(_06962_),
    .X(_00619_));
 sky130_fd_sc_hd__buf_2 _12914_ (.A(_06174_),
    .X(_06963_));
 sky130_fd_sc_hd__buf_6 _12915_ (.A(_06942_),
    .X(_06964_));
 sky130_fd_sc_hd__mux2_1 _12916_ (.A0(_06963_),
    .A1(\cpuregs.regs[31][10] ),
    .S(_06964_),
    .X(_06965_));
 sky130_fd_sc_hd__clkbuf_1 _12917_ (.A(_06965_),
    .X(_00620_));
 sky130_fd_sc_hd__buf_2 _12918_ (.A(_06183_),
    .X(_06966_));
 sky130_fd_sc_hd__mux2_1 _12919_ (.A0(_06966_),
    .A1(\cpuregs.regs[31][11] ),
    .S(_06964_),
    .X(_06967_));
 sky130_fd_sc_hd__clkbuf_1 _12920_ (.A(_06967_),
    .X(_00621_));
 sky130_fd_sc_hd__buf_2 _12921_ (.A(_06192_),
    .X(_06968_));
 sky130_fd_sc_hd__mux2_1 _12922_ (.A0(_06968_),
    .A1(\cpuregs.regs[31][12] ),
    .S(_06964_),
    .X(_06969_));
 sky130_fd_sc_hd__clkbuf_1 _12923_ (.A(_06969_),
    .X(_00622_));
 sky130_fd_sc_hd__buf_2 _12924_ (.A(_06200_),
    .X(_06970_));
 sky130_fd_sc_hd__mux2_1 _12925_ (.A0(_06970_),
    .A1(\cpuregs.regs[31][13] ),
    .S(_06964_),
    .X(_06971_));
 sky130_fd_sc_hd__clkbuf_1 _12926_ (.A(_06971_),
    .X(_00623_));
 sky130_fd_sc_hd__buf_2 _12927_ (.A(_06207_),
    .X(_06972_));
 sky130_fd_sc_hd__mux2_1 _12928_ (.A0(_06972_),
    .A1(\cpuregs.regs[31][14] ),
    .S(_06964_),
    .X(_06973_));
 sky130_fd_sc_hd__clkbuf_1 _12929_ (.A(_06973_),
    .X(_00624_));
 sky130_fd_sc_hd__clkbuf_4 _12930_ (.A(_06215_),
    .X(_06974_));
 sky130_fd_sc_hd__mux2_1 _12931_ (.A0(_06974_),
    .A1(\cpuregs.regs[31][15] ),
    .S(_06964_),
    .X(_06975_));
 sky130_fd_sc_hd__clkbuf_1 _12932_ (.A(_06975_),
    .X(_00625_));
 sky130_fd_sc_hd__buf_2 _12933_ (.A(_06223_),
    .X(_06976_));
 sky130_fd_sc_hd__mux2_1 _12934_ (.A0(_06976_),
    .A1(\cpuregs.regs[31][16] ),
    .S(_06964_),
    .X(_06977_));
 sky130_fd_sc_hd__clkbuf_1 _12935_ (.A(_06977_),
    .X(_00626_));
 sky130_fd_sc_hd__buf_2 _12936_ (.A(_06231_),
    .X(_06978_));
 sky130_fd_sc_hd__mux2_1 _12937_ (.A0(_06978_),
    .A1(\cpuregs.regs[31][17] ),
    .S(_06964_),
    .X(_06979_));
 sky130_fd_sc_hd__clkbuf_1 _12938_ (.A(_06979_),
    .X(_00627_));
 sky130_fd_sc_hd__buf_2 _12939_ (.A(_06239_),
    .X(_06980_));
 sky130_fd_sc_hd__mux2_1 _12940_ (.A0(_06980_),
    .A1(\cpuregs.regs[31][18] ),
    .S(_06964_),
    .X(_06981_));
 sky130_fd_sc_hd__clkbuf_1 _12941_ (.A(_06981_),
    .X(_00628_));
 sky130_fd_sc_hd__buf_2 _12942_ (.A(_06247_),
    .X(_06982_));
 sky130_fd_sc_hd__mux2_1 _12943_ (.A0(_06982_),
    .A1(\cpuregs.regs[31][19] ),
    .S(_06964_),
    .X(_06983_));
 sky130_fd_sc_hd__clkbuf_1 _12944_ (.A(_06983_),
    .X(_00629_));
 sky130_fd_sc_hd__buf_2 _12945_ (.A(_06256_),
    .X(_06984_));
 sky130_fd_sc_hd__buf_6 _12946_ (.A(_06942_),
    .X(_06985_));
 sky130_fd_sc_hd__mux2_1 _12947_ (.A0(_06984_),
    .A1(\cpuregs.regs[31][20] ),
    .S(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__clkbuf_1 _12948_ (.A(_06986_),
    .X(_00630_));
 sky130_fd_sc_hd__buf_2 _12949_ (.A(_06265_),
    .X(_06987_));
 sky130_fd_sc_hd__mux2_1 _12950_ (.A0(_06987_),
    .A1(\cpuregs.regs[31][21] ),
    .S(_06985_),
    .X(_06988_));
 sky130_fd_sc_hd__clkbuf_1 _12951_ (.A(_06988_),
    .X(_00631_));
 sky130_fd_sc_hd__buf_2 _12952_ (.A(_06273_),
    .X(_06989_));
 sky130_fd_sc_hd__mux2_1 _12953_ (.A0(_06989_),
    .A1(\cpuregs.regs[31][22] ),
    .S(_06985_),
    .X(_06990_));
 sky130_fd_sc_hd__clkbuf_1 _12954_ (.A(_06990_),
    .X(_00632_));
 sky130_fd_sc_hd__buf_2 _12955_ (.A(_06280_),
    .X(_06991_));
 sky130_fd_sc_hd__mux2_1 _12956_ (.A0(_06991_),
    .A1(\cpuregs.regs[31][23] ),
    .S(_06985_),
    .X(_06992_));
 sky130_fd_sc_hd__clkbuf_1 _12957_ (.A(_06992_),
    .X(_00633_));
 sky130_fd_sc_hd__buf_2 _12958_ (.A(_06288_),
    .X(_06993_));
 sky130_fd_sc_hd__mux2_1 _12959_ (.A0(_06993_),
    .A1(\cpuregs.regs[31][24] ),
    .S(_06985_),
    .X(_06994_));
 sky130_fd_sc_hd__clkbuf_1 _12960_ (.A(_06994_),
    .X(_00634_));
 sky130_fd_sc_hd__buf_2 _12961_ (.A(_06296_),
    .X(_06995_));
 sky130_fd_sc_hd__mux2_1 _12962_ (.A0(_06995_),
    .A1(\cpuregs.regs[31][25] ),
    .S(_06985_),
    .X(_06996_));
 sky130_fd_sc_hd__clkbuf_1 _12963_ (.A(_06996_),
    .X(_00635_));
 sky130_fd_sc_hd__buf_2 _12964_ (.A(_06303_),
    .X(_06997_));
 sky130_fd_sc_hd__mux2_1 _12965_ (.A0(_06997_),
    .A1(\cpuregs.regs[31][26] ),
    .S(_06985_),
    .X(_06998_));
 sky130_fd_sc_hd__clkbuf_1 _12966_ (.A(_06998_),
    .X(_00636_));
 sky130_fd_sc_hd__buf_2 _12967_ (.A(_06311_),
    .X(_06999_));
 sky130_fd_sc_hd__mux2_1 _12968_ (.A0(_06999_),
    .A1(\cpuregs.regs[31][27] ),
    .S(_06985_),
    .X(_07000_));
 sky130_fd_sc_hd__clkbuf_1 _12969_ (.A(_07000_),
    .X(_00637_));
 sky130_fd_sc_hd__buf_2 _12970_ (.A(_06319_),
    .X(_07001_));
 sky130_fd_sc_hd__mux2_1 _12971_ (.A0(_07001_),
    .A1(\cpuregs.regs[31][28] ),
    .S(_06985_),
    .X(_07002_));
 sky130_fd_sc_hd__clkbuf_1 _12972_ (.A(_07002_),
    .X(_00638_));
 sky130_fd_sc_hd__buf_2 _12973_ (.A(_06327_),
    .X(_07003_));
 sky130_fd_sc_hd__mux2_1 _12974_ (.A0(_07003_),
    .A1(\cpuregs.regs[31][29] ),
    .S(_06985_),
    .X(_07004_));
 sky130_fd_sc_hd__clkbuf_1 _12975_ (.A(_07004_),
    .X(_00639_));
 sky130_fd_sc_hd__buf_2 _12976_ (.A(_06335_),
    .X(_07005_));
 sky130_fd_sc_hd__mux2_1 _12977_ (.A0(_07005_),
    .A1(\cpuregs.regs[31][30] ),
    .S(_06942_),
    .X(_07006_));
 sky130_fd_sc_hd__clkbuf_1 _12978_ (.A(_07006_),
    .X(_00640_));
 sky130_fd_sc_hd__buf_2 _12979_ (.A(_06342_),
    .X(_07007_));
 sky130_fd_sc_hd__mux2_1 _12980_ (.A0(_07007_),
    .A1(\cpuregs.regs[31][31] ),
    .S(_06942_),
    .X(_07008_));
 sky130_fd_sc_hd__clkbuf_1 _12981_ (.A(_07008_),
    .X(_00641_));
 sky130_fd_sc_hd__nor2_4 _12982_ (.A(_06676_),
    .B(_06750_),
    .Y(_07009_));
 sky130_fd_sc_hd__buf_6 _12983_ (.A(_07009_),
    .X(_07010_));
 sky130_fd_sc_hd__mux2_1 _12984_ (.A0(\cpuregs.regs[3][0] ),
    .A1(_06531_),
    .S(_07010_),
    .X(_07011_));
 sky130_fd_sc_hd__clkbuf_1 _12985_ (.A(_07011_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _12986_ (.A0(\cpuregs.regs[3][1] ),
    .A1(_06536_),
    .S(_07010_),
    .X(_07012_));
 sky130_fd_sc_hd__clkbuf_1 _12987_ (.A(_07012_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _12988_ (.A0(\cpuregs.regs[3][2] ),
    .A1(_06538_),
    .S(_07010_),
    .X(_07013_));
 sky130_fd_sc_hd__clkbuf_1 _12989_ (.A(_07013_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _12990_ (.A0(\cpuregs.regs[3][3] ),
    .A1(_06540_),
    .S(_07010_),
    .X(_07014_));
 sky130_fd_sc_hd__clkbuf_1 _12991_ (.A(_07014_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _12992_ (.A0(\cpuregs.regs[3][4] ),
    .A1(_06542_),
    .S(_07010_),
    .X(_07015_));
 sky130_fd_sc_hd__clkbuf_1 _12993_ (.A(_07015_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _12994_ (.A0(\cpuregs.regs[3][5] ),
    .A1(_06544_),
    .S(_07010_),
    .X(_07016_));
 sky130_fd_sc_hd__clkbuf_1 _12995_ (.A(_07016_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _12996_ (.A0(\cpuregs.regs[3][6] ),
    .A1(_06546_),
    .S(_07010_),
    .X(_07017_));
 sky130_fd_sc_hd__clkbuf_1 _12997_ (.A(_07017_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _12998_ (.A0(\cpuregs.regs[3][7] ),
    .A1(_06548_),
    .S(_07010_),
    .X(_07018_));
 sky130_fd_sc_hd__clkbuf_1 _12999_ (.A(_07018_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _13000_ (.A0(\cpuregs.regs[3][8] ),
    .A1(_06550_),
    .S(_07010_),
    .X(_07019_));
 sky130_fd_sc_hd__clkbuf_1 _13001_ (.A(_07019_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _13002_ (.A0(\cpuregs.regs[3][9] ),
    .A1(_06552_),
    .S(_07010_),
    .X(_07020_));
 sky130_fd_sc_hd__clkbuf_1 _13003_ (.A(_07020_),
    .X(_00651_));
 sky130_fd_sc_hd__clkbuf_8 _13004_ (.A(_07009_),
    .X(_07021_));
 sky130_fd_sc_hd__mux2_1 _13005_ (.A0(\cpuregs.regs[3][10] ),
    .A1(_06554_),
    .S(_07021_),
    .X(_07022_));
 sky130_fd_sc_hd__clkbuf_1 _13006_ (.A(_07022_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _13007_ (.A0(\cpuregs.regs[3][11] ),
    .A1(_06557_),
    .S(_07021_),
    .X(_07023_));
 sky130_fd_sc_hd__clkbuf_1 _13008_ (.A(_07023_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _13009_ (.A0(\cpuregs.regs[3][12] ),
    .A1(_06559_),
    .S(_07021_),
    .X(_07024_));
 sky130_fd_sc_hd__clkbuf_1 _13010_ (.A(_07024_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _13011_ (.A0(\cpuregs.regs[3][13] ),
    .A1(_06561_),
    .S(_07021_),
    .X(_07025_));
 sky130_fd_sc_hd__clkbuf_1 _13012_ (.A(_07025_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _13013_ (.A0(\cpuregs.regs[3][14] ),
    .A1(_06563_),
    .S(_07021_),
    .X(_07026_));
 sky130_fd_sc_hd__clkbuf_1 _13014_ (.A(_07026_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _13015_ (.A0(\cpuregs.regs[3][15] ),
    .A1(_06565_),
    .S(_07021_),
    .X(_07027_));
 sky130_fd_sc_hd__clkbuf_1 _13016_ (.A(_07027_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _13017_ (.A0(\cpuregs.regs[3][16] ),
    .A1(_06567_),
    .S(_07021_),
    .X(_07028_));
 sky130_fd_sc_hd__clkbuf_1 _13018_ (.A(_07028_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _13019_ (.A0(\cpuregs.regs[3][17] ),
    .A1(_06569_),
    .S(_07021_),
    .X(_07029_));
 sky130_fd_sc_hd__clkbuf_1 _13020_ (.A(_07029_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _13021_ (.A0(\cpuregs.regs[3][18] ),
    .A1(_06571_),
    .S(_07021_),
    .X(_07030_));
 sky130_fd_sc_hd__clkbuf_1 _13022_ (.A(_07030_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _13023_ (.A0(\cpuregs.regs[3][19] ),
    .A1(_06573_),
    .S(_07021_),
    .X(_07031_));
 sky130_fd_sc_hd__clkbuf_1 _13024_ (.A(_07031_),
    .X(_00661_));
 sky130_fd_sc_hd__buf_6 _13025_ (.A(_07009_),
    .X(_07032_));
 sky130_fd_sc_hd__mux2_1 _13026_ (.A0(\cpuregs.regs[3][20] ),
    .A1(_06575_),
    .S(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__clkbuf_1 _13027_ (.A(_07033_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _13028_ (.A0(\cpuregs.regs[3][21] ),
    .A1(_06578_),
    .S(_07032_),
    .X(_07034_));
 sky130_fd_sc_hd__clkbuf_1 _13029_ (.A(_07034_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _13030_ (.A0(\cpuregs.regs[3][22] ),
    .A1(_06580_),
    .S(_07032_),
    .X(_07035_));
 sky130_fd_sc_hd__clkbuf_1 _13031_ (.A(_07035_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _13032_ (.A0(\cpuregs.regs[3][23] ),
    .A1(_06582_),
    .S(_07032_),
    .X(_07036_));
 sky130_fd_sc_hd__clkbuf_1 _13033_ (.A(_07036_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _13034_ (.A0(\cpuregs.regs[3][24] ),
    .A1(_06584_),
    .S(_07032_),
    .X(_07037_));
 sky130_fd_sc_hd__clkbuf_1 _13035_ (.A(_07037_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _13036_ (.A0(\cpuregs.regs[3][25] ),
    .A1(_06586_),
    .S(_07032_),
    .X(_07038_));
 sky130_fd_sc_hd__clkbuf_1 _13037_ (.A(_07038_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _13038_ (.A0(\cpuregs.regs[3][26] ),
    .A1(_06588_),
    .S(_07032_),
    .X(_07039_));
 sky130_fd_sc_hd__clkbuf_1 _13039_ (.A(_07039_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _13040_ (.A0(\cpuregs.regs[3][27] ),
    .A1(_06590_),
    .S(_07032_),
    .X(_07040_));
 sky130_fd_sc_hd__clkbuf_1 _13041_ (.A(_07040_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _13042_ (.A0(\cpuregs.regs[3][28] ),
    .A1(_06592_),
    .S(_07032_),
    .X(_07041_));
 sky130_fd_sc_hd__clkbuf_1 _13043_ (.A(_07041_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _13044_ (.A0(\cpuregs.regs[3][29] ),
    .A1(_06594_),
    .S(_07032_),
    .X(_07042_));
 sky130_fd_sc_hd__clkbuf_1 _13045_ (.A(_07042_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _13046_ (.A0(\cpuregs.regs[3][30] ),
    .A1(_06596_),
    .S(_07009_),
    .X(_07043_));
 sky130_fd_sc_hd__clkbuf_1 _13047_ (.A(_07043_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _13048_ (.A0(\cpuregs.regs[3][31] ),
    .A1(_06598_),
    .S(_07009_),
    .X(_07044_));
 sky130_fd_sc_hd__clkbuf_1 _13049_ (.A(_07044_),
    .X(_00673_));
 sky130_fd_sc_hd__nand2_4 _13050_ (.A(_06346_),
    .B(_06904_),
    .Y(_07045_));
 sky130_fd_sc_hd__buf_6 _13051_ (.A(_07045_),
    .X(_07046_));
 sky130_fd_sc_hd__mux2_1 _13052_ (.A0(_06941_),
    .A1(\cpuregs.regs[7][0] ),
    .S(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__clkbuf_1 _13053_ (.A(_07047_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _13054_ (.A0(_06945_),
    .A1(\cpuregs.regs[7][1] ),
    .S(_07046_),
    .X(_07048_));
 sky130_fd_sc_hd__clkbuf_1 _13055_ (.A(_07048_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _13056_ (.A0(_06947_),
    .A1(\cpuregs.regs[7][2] ),
    .S(_07046_),
    .X(_07049_));
 sky130_fd_sc_hd__clkbuf_1 _13057_ (.A(_07049_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _13058_ (.A0(_06949_),
    .A1(\cpuregs.regs[7][3] ),
    .S(_07046_),
    .X(_07050_));
 sky130_fd_sc_hd__clkbuf_1 _13059_ (.A(_07050_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _13060_ (.A0(_06951_),
    .A1(\cpuregs.regs[7][4] ),
    .S(_07046_),
    .X(_07051_));
 sky130_fd_sc_hd__clkbuf_1 _13061_ (.A(_07051_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _13062_ (.A0(_06953_),
    .A1(\cpuregs.regs[7][5] ),
    .S(_07046_),
    .X(_07052_));
 sky130_fd_sc_hd__clkbuf_1 _13063_ (.A(_07052_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _13064_ (.A0(_06955_),
    .A1(\cpuregs.regs[7][6] ),
    .S(_07046_),
    .X(_07053_));
 sky130_fd_sc_hd__clkbuf_1 _13065_ (.A(_07053_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _13066_ (.A0(_06957_),
    .A1(\cpuregs.regs[7][7] ),
    .S(_07046_),
    .X(_07054_));
 sky130_fd_sc_hd__clkbuf_1 _13067_ (.A(_07054_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _13068_ (.A0(_06959_),
    .A1(\cpuregs.regs[7][8] ),
    .S(_07046_),
    .X(_07055_));
 sky130_fd_sc_hd__clkbuf_1 _13069_ (.A(_07055_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _13070_ (.A0(_06961_),
    .A1(\cpuregs.regs[7][9] ),
    .S(_07046_),
    .X(_07056_));
 sky130_fd_sc_hd__clkbuf_1 _13071_ (.A(_07056_),
    .X(_00683_));
 sky130_fd_sc_hd__clkbuf_8 _13072_ (.A(_07045_),
    .X(_07057_));
 sky130_fd_sc_hd__mux2_1 _13073_ (.A0(_06963_),
    .A1(\cpuregs.regs[7][10] ),
    .S(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__clkbuf_1 _13074_ (.A(_07058_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _13075_ (.A0(_06966_),
    .A1(\cpuregs.regs[7][11] ),
    .S(_07057_),
    .X(_07059_));
 sky130_fd_sc_hd__clkbuf_1 _13076_ (.A(_07059_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _13077_ (.A0(_06968_),
    .A1(\cpuregs.regs[7][12] ),
    .S(_07057_),
    .X(_07060_));
 sky130_fd_sc_hd__clkbuf_1 _13078_ (.A(_07060_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _13079_ (.A0(_06970_),
    .A1(\cpuregs.regs[7][13] ),
    .S(_07057_),
    .X(_07061_));
 sky130_fd_sc_hd__clkbuf_1 _13080_ (.A(_07061_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _13081_ (.A0(_06972_),
    .A1(\cpuregs.regs[7][14] ),
    .S(_07057_),
    .X(_07062_));
 sky130_fd_sc_hd__clkbuf_1 _13082_ (.A(_07062_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _13083_ (.A0(_06974_),
    .A1(\cpuregs.regs[7][15] ),
    .S(_07057_),
    .X(_07063_));
 sky130_fd_sc_hd__clkbuf_1 _13084_ (.A(_07063_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _13085_ (.A0(_06976_),
    .A1(\cpuregs.regs[7][16] ),
    .S(_07057_),
    .X(_07064_));
 sky130_fd_sc_hd__clkbuf_1 _13086_ (.A(_07064_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _13087_ (.A0(_06978_),
    .A1(\cpuregs.regs[7][17] ),
    .S(_07057_),
    .X(_07065_));
 sky130_fd_sc_hd__clkbuf_1 _13088_ (.A(_07065_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _13089_ (.A0(_06980_),
    .A1(\cpuregs.regs[7][18] ),
    .S(_07057_),
    .X(_07066_));
 sky130_fd_sc_hd__clkbuf_1 _13090_ (.A(_07066_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _13091_ (.A0(_06982_),
    .A1(\cpuregs.regs[7][19] ),
    .S(_07057_),
    .X(_07067_));
 sky130_fd_sc_hd__clkbuf_1 _13092_ (.A(_07067_),
    .X(_00693_));
 sky130_fd_sc_hd__clkbuf_8 _13093_ (.A(_07045_),
    .X(_07068_));
 sky130_fd_sc_hd__mux2_1 _13094_ (.A0(_06984_),
    .A1(\cpuregs.regs[7][20] ),
    .S(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__clkbuf_1 _13095_ (.A(_07069_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _13096_ (.A0(_06987_),
    .A1(\cpuregs.regs[7][21] ),
    .S(_07068_),
    .X(_07070_));
 sky130_fd_sc_hd__clkbuf_1 _13097_ (.A(_07070_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _13098_ (.A0(_06989_),
    .A1(\cpuregs.regs[7][22] ),
    .S(_07068_),
    .X(_07071_));
 sky130_fd_sc_hd__clkbuf_1 _13099_ (.A(_07071_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _13100_ (.A0(_06991_),
    .A1(\cpuregs.regs[7][23] ),
    .S(_07068_),
    .X(_07072_));
 sky130_fd_sc_hd__clkbuf_1 _13101_ (.A(_07072_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _13102_ (.A0(_06993_),
    .A1(\cpuregs.regs[7][24] ),
    .S(_07068_),
    .X(_07073_));
 sky130_fd_sc_hd__clkbuf_1 _13103_ (.A(_07073_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _13104_ (.A0(_06995_),
    .A1(\cpuregs.regs[7][25] ),
    .S(_07068_),
    .X(_07074_));
 sky130_fd_sc_hd__clkbuf_1 _13105_ (.A(_07074_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _13106_ (.A0(_06997_),
    .A1(\cpuregs.regs[7][26] ),
    .S(_07068_),
    .X(_07075_));
 sky130_fd_sc_hd__clkbuf_1 _13107_ (.A(_07075_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _13108_ (.A0(_06999_),
    .A1(\cpuregs.regs[7][27] ),
    .S(_07068_),
    .X(_07076_));
 sky130_fd_sc_hd__clkbuf_1 _13109_ (.A(_07076_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _13110_ (.A0(_07001_),
    .A1(\cpuregs.regs[7][28] ),
    .S(_07068_),
    .X(_07077_));
 sky130_fd_sc_hd__clkbuf_1 _13111_ (.A(_07077_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _13112_ (.A0(_07003_),
    .A1(\cpuregs.regs[7][29] ),
    .S(_07068_),
    .X(_07078_));
 sky130_fd_sc_hd__clkbuf_1 _13113_ (.A(_07078_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _13114_ (.A0(_07005_),
    .A1(\cpuregs.regs[7][30] ),
    .S(_07045_),
    .X(_07079_));
 sky130_fd_sc_hd__clkbuf_1 _13115_ (.A(_07079_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _13116_ (.A0(_07007_),
    .A1(\cpuregs.regs[7][31] ),
    .S(_07045_),
    .X(_07080_));
 sky130_fd_sc_hd__clkbuf_1 _13117_ (.A(_07080_),
    .X(_00705_));
 sky130_fd_sc_hd__nand2_4 _13118_ (.A(_06383_),
    .B(_06904_),
    .Y(_07081_));
 sky130_fd_sc_hd__buf_6 _13119_ (.A(_07081_),
    .X(_07082_));
 sky130_fd_sc_hd__mux2_1 _13120_ (.A0(_06941_),
    .A1(\cpuregs.regs[4][0] ),
    .S(_07082_),
    .X(_07083_));
 sky130_fd_sc_hd__clkbuf_1 _13121_ (.A(_07083_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _13122_ (.A0(_06945_),
    .A1(\cpuregs.regs[4][1] ),
    .S(_07082_),
    .X(_07084_));
 sky130_fd_sc_hd__clkbuf_1 _13123_ (.A(_07084_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _13124_ (.A0(_06947_),
    .A1(\cpuregs.regs[4][2] ),
    .S(_07082_),
    .X(_07085_));
 sky130_fd_sc_hd__clkbuf_1 _13125_ (.A(_07085_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _13126_ (.A0(_06949_),
    .A1(\cpuregs.regs[4][3] ),
    .S(_07082_),
    .X(_07086_));
 sky130_fd_sc_hd__clkbuf_1 _13127_ (.A(_07086_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _13128_ (.A0(_06951_),
    .A1(\cpuregs.regs[4][4] ),
    .S(_07082_),
    .X(_07087_));
 sky130_fd_sc_hd__clkbuf_1 _13129_ (.A(_07087_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _13130_ (.A0(_06953_),
    .A1(\cpuregs.regs[4][5] ),
    .S(_07082_),
    .X(_07088_));
 sky130_fd_sc_hd__clkbuf_1 _13131_ (.A(_07088_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _13132_ (.A0(_06955_),
    .A1(\cpuregs.regs[4][6] ),
    .S(_07082_),
    .X(_07089_));
 sky130_fd_sc_hd__clkbuf_1 _13133_ (.A(_07089_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _13134_ (.A0(_06957_),
    .A1(\cpuregs.regs[4][7] ),
    .S(_07082_),
    .X(_07090_));
 sky130_fd_sc_hd__clkbuf_1 _13135_ (.A(_07090_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _13136_ (.A0(_06959_),
    .A1(\cpuregs.regs[4][8] ),
    .S(_07082_),
    .X(_07091_));
 sky130_fd_sc_hd__clkbuf_1 _13137_ (.A(_07091_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _13138_ (.A0(_06961_),
    .A1(\cpuregs.regs[4][9] ),
    .S(_07082_),
    .X(_07092_));
 sky130_fd_sc_hd__clkbuf_1 _13139_ (.A(_07092_),
    .X(_00715_));
 sky130_fd_sc_hd__clkbuf_8 _13140_ (.A(_07081_),
    .X(_07093_));
 sky130_fd_sc_hd__mux2_1 _13141_ (.A0(_06963_),
    .A1(\cpuregs.regs[4][10] ),
    .S(_07093_),
    .X(_07094_));
 sky130_fd_sc_hd__clkbuf_1 _13142_ (.A(_07094_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _13143_ (.A0(_06966_),
    .A1(\cpuregs.regs[4][11] ),
    .S(_07093_),
    .X(_07095_));
 sky130_fd_sc_hd__clkbuf_1 _13144_ (.A(_07095_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _13145_ (.A0(_06968_),
    .A1(\cpuregs.regs[4][12] ),
    .S(_07093_),
    .X(_07096_));
 sky130_fd_sc_hd__clkbuf_1 _13146_ (.A(_07096_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _13147_ (.A0(_06970_),
    .A1(\cpuregs.regs[4][13] ),
    .S(_07093_),
    .X(_07097_));
 sky130_fd_sc_hd__clkbuf_1 _13148_ (.A(_07097_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _13149_ (.A0(_06972_),
    .A1(\cpuregs.regs[4][14] ),
    .S(_07093_),
    .X(_07098_));
 sky130_fd_sc_hd__clkbuf_1 _13150_ (.A(_07098_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _13151_ (.A0(_06974_),
    .A1(\cpuregs.regs[4][15] ),
    .S(_07093_),
    .X(_07099_));
 sky130_fd_sc_hd__clkbuf_1 _13152_ (.A(_07099_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _13153_ (.A0(_06976_),
    .A1(\cpuregs.regs[4][16] ),
    .S(_07093_),
    .X(_07100_));
 sky130_fd_sc_hd__clkbuf_1 _13154_ (.A(_07100_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _13155_ (.A0(_06978_),
    .A1(\cpuregs.regs[4][17] ),
    .S(_07093_),
    .X(_07101_));
 sky130_fd_sc_hd__clkbuf_1 _13156_ (.A(_07101_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _13157_ (.A0(_06980_),
    .A1(\cpuregs.regs[4][18] ),
    .S(_07093_),
    .X(_07102_));
 sky130_fd_sc_hd__clkbuf_1 _13158_ (.A(_07102_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _13159_ (.A0(_06982_),
    .A1(\cpuregs.regs[4][19] ),
    .S(_07093_),
    .X(_07103_));
 sky130_fd_sc_hd__clkbuf_1 _13160_ (.A(_07103_),
    .X(_00725_));
 sky130_fd_sc_hd__clkbuf_8 _13161_ (.A(_07081_),
    .X(_07104_));
 sky130_fd_sc_hd__mux2_1 _13162_ (.A0(_06984_),
    .A1(\cpuregs.regs[4][20] ),
    .S(_07104_),
    .X(_07105_));
 sky130_fd_sc_hd__clkbuf_1 _13163_ (.A(_07105_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _13164_ (.A0(_06987_),
    .A1(\cpuregs.regs[4][21] ),
    .S(_07104_),
    .X(_07106_));
 sky130_fd_sc_hd__clkbuf_1 _13165_ (.A(_07106_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _13166_ (.A0(_06989_),
    .A1(\cpuregs.regs[4][22] ),
    .S(_07104_),
    .X(_07107_));
 sky130_fd_sc_hd__clkbuf_1 _13167_ (.A(_07107_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _13168_ (.A0(_06991_),
    .A1(\cpuregs.regs[4][23] ),
    .S(_07104_),
    .X(_07108_));
 sky130_fd_sc_hd__clkbuf_1 _13169_ (.A(_07108_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _13170_ (.A0(_06993_),
    .A1(\cpuregs.regs[4][24] ),
    .S(_07104_),
    .X(_07109_));
 sky130_fd_sc_hd__clkbuf_1 _13171_ (.A(_07109_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _13172_ (.A0(_06995_),
    .A1(\cpuregs.regs[4][25] ),
    .S(_07104_),
    .X(_07110_));
 sky130_fd_sc_hd__clkbuf_1 _13173_ (.A(_07110_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _13174_ (.A0(_06997_),
    .A1(\cpuregs.regs[4][26] ),
    .S(_07104_),
    .X(_07111_));
 sky130_fd_sc_hd__clkbuf_1 _13175_ (.A(_07111_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _13176_ (.A0(_06999_),
    .A1(\cpuregs.regs[4][27] ),
    .S(_07104_),
    .X(_07112_));
 sky130_fd_sc_hd__clkbuf_1 _13177_ (.A(_07112_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _13178_ (.A0(_07001_),
    .A1(\cpuregs.regs[4][28] ),
    .S(_07104_),
    .X(_07113_));
 sky130_fd_sc_hd__clkbuf_1 _13179_ (.A(_07113_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _13180_ (.A0(_07003_),
    .A1(\cpuregs.regs[4][29] ),
    .S(_07104_),
    .X(_07114_));
 sky130_fd_sc_hd__clkbuf_1 _13181_ (.A(_07114_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _13182_ (.A0(_07005_),
    .A1(\cpuregs.regs[4][30] ),
    .S(_07081_),
    .X(_07115_));
 sky130_fd_sc_hd__clkbuf_1 _13183_ (.A(_07115_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _13184_ (.A0(_07007_),
    .A1(\cpuregs.regs[4][31] ),
    .S(_07081_),
    .X(_07116_));
 sky130_fd_sc_hd__clkbuf_1 _13185_ (.A(_07116_),
    .X(_00737_));
 sky130_fd_sc_hd__nand2_2 _13186_ (.A(_06383_),
    .B(_06084_),
    .Y(_07117_));
 sky130_fd_sc_hd__buf_6 _13187_ (.A(_07117_),
    .X(_07118_));
 sky130_fd_sc_hd__mux2_1 _13188_ (.A0(_06941_),
    .A1(\cpuregs.regs[8][0] ),
    .S(_07118_),
    .X(_07119_));
 sky130_fd_sc_hd__clkbuf_1 _13189_ (.A(_07119_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _13190_ (.A0(_06945_),
    .A1(\cpuregs.regs[8][1] ),
    .S(_07118_),
    .X(_07120_));
 sky130_fd_sc_hd__clkbuf_1 _13191_ (.A(_07120_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _13192_ (.A0(_06947_),
    .A1(\cpuregs.regs[8][2] ),
    .S(_07118_),
    .X(_07121_));
 sky130_fd_sc_hd__clkbuf_1 _13193_ (.A(_07121_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _13194_ (.A0(_06949_),
    .A1(\cpuregs.regs[8][3] ),
    .S(_07118_),
    .X(_07122_));
 sky130_fd_sc_hd__clkbuf_1 _13195_ (.A(_07122_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _13196_ (.A0(_06951_),
    .A1(\cpuregs.regs[8][4] ),
    .S(_07118_),
    .X(_07123_));
 sky130_fd_sc_hd__clkbuf_1 _13197_ (.A(_07123_),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _13198_ (.A0(_06953_),
    .A1(\cpuregs.regs[8][5] ),
    .S(_07118_),
    .X(_07124_));
 sky130_fd_sc_hd__clkbuf_1 _13199_ (.A(_07124_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _13200_ (.A0(_06955_),
    .A1(\cpuregs.regs[8][6] ),
    .S(_07118_),
    .X(_07125_));
 sky130_fd_sc_hd__clkbuf_1 _13201_ (.A(_07125_),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _13202_ (.A0(_06957_),
    .A1(\cpuregs.regs[8][7] ),
    .S(_07118_),
    .X(_07126_));
 sky130_fd_sc_hd__clkbuf_1 _13203_ (.A(_07126_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _13204_ (.A0(_06959_),
    .A1(\cpuregs.regs[8][8] ),
    .S(_07118_),
    .X(_07127_));
 sky130_fd_sc_hd__clkbuf_1 _13205_ (.A(_07127_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _13206_ (.A0(_06961_),
    .A1(\cpuregs.regs[8][9] ),
    .S(_07118_),
    .X(_07128_));
 sky130_fd_sc_hd__clkbuf_1 _13207_ (.A(_07128_),
    .X(_00747_));
 sky130_fd_sc_hd__clkbuf_8 _13208_ (.A(_07117_),
    .X(_07129_));
 sky130_fd_sc_hd__mux2_1 _13209_ (.A0(_06963_),
    .A1(\cpuregs.regs[8][10] ),
    .S(_07129_),
    .X(_07130_));
 sky130_fd_sc_hd__clkbuf_1 _13210_ (.A(_07130_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _13211_ (.A0(_06966_),
    .A1(\cpuregs.regs[8][11] ),
    .S(_07129_),
    .X(_07131_));
 sky130_fd_sc_hd__clkbuf_1 _13212_ (.A(_07131_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _13213_ (.A0(_06968_),
    .A1(\cpuregs.regs[8][12] ),
    .S(_07129_),
    .X(_07132_));
 sky130_fd_sc_hd__clkbuf_1 _13214_ (.A(_07132_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _13215_ (.A0(_06970_),
    .A1(\cpuregs.regs[8][13] ),
    .S(_07129_),
    .X(_07133_));
 sky130_fd_sc_hd__clkbuf_1 _13216_ (.A(_07133_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _13217_ (.A0(_06972_),
    .A1(\cpuregs.regs[8][14] ),
    .S(_07129_),
    .X(_07134_));
 sky130_fd_sc_hd__clkbuf_1 _13218_ (.A(_07134_),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _13219_ (.A0(_06974_),
    .A1(\cpuregs.regs[8][15] ),
    .S(_07129_),
    .X(_07135_));
 sky130_fd_sc_hd__clkbuf_1 _13220_ (.A(_07135_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _13221_ (.A0(_06976_),
    .A1(\cpuregs.regs[8][16] ),
    .S(_07129_),
    .X(_07136_));
 sky130_fd_sc_hd__clkbuf_1 _13222_ (.A(_07136_),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _13223_ (.A0(_06978_),
    .A1(\cpuregs.regs[8][17] ),
    .S(_07129_),
    .X(_07137_));
 sky130_fd_sc_hd__clkbuf_1 _13224_ (.A(_07137_),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_1 _13225_ (.A0(_06980_),
    .A1(\cpuregs.regs[8][18] ),
    .S(_07129_),
    .X(_07138_));
 sky130_fd_sc_hd__clkbuf_1 _13226_ (.A(_07138_),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _13227_ (.A0(_06982_),
    .A1(\cpuregs.regs[8][19] ),
    .S(_07129_),
    .X(_07139_));
 sky130_fd_sc_hd__clkbuf_1 _13228_ (.A(_07139_),
    .X(_00757_));
 sky130_fd_sc_hd__buf_6 _13229_ (.A(_07117_),
    .X(_07140_));
 sky130_fd_sc_hd__mux2_1 _13230_ (.A0(_06984_),
    .A1(\cpuregs.regs[8][20] ),
    .S(_07140_),
    .X(_07141_));
 sky130_fd_sc_hd__clkbuf_1 _13231_ (.A(_07141_),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _13232_ (.A0(_06987_),
    .A1(\cpuregs.regs[8][21] ),
    .S(_07140_),
    .X(_07142_));
 sky130_fd_sc_hd__clkbuf_1 _13233_ (.A(_07142_),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _13234_ (.A0(_06989_),
    .A1(\cpuregs.regs[8][22] ),
    .S(_07140_),
    .X(_07143_));
 sky130_fd_sc_hd__clkbuf_1 _13235_ (.A(_07143_),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _13236_ (.A0(_06991_),
    .A1(\cpuregs.regs[8][23] ),
    .S(_07140_),
    .X(_07144_));
 sky130_fd_sc_hd__clkbuf_1 _13237_ (.A(_07144_),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _13238_ (.A0(_06993_),
    .A1(\cpuregs.regs[8][24] ),
    .S(_07140_),
    .X(_07145_));
 sky130_fd_sc_hd__clkbuf_1 _13239_ (.A(_07145_),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _13240_ (.A0(_06995_),
    .A1(\cpuregs.regs[8][25] ),
    .S(_07140_),
    .X(_07146_));
 sky130_fd_sc_hd__clkbuf_1 _13241_ (.A(_07146_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _13242_ (.A0(_06997_),
    .A1(\cpuregs.regs[8][26] ),
    .S(_07140_),
    .X(_07147_));
 sky130_fd_sc_hd__clkbuf_1 _13243_ (.A(_07147_),
    .X(_00764_));
 sky130_fd_sc_hd__mux2_1 _13244_ (.A0(_06999_),
    .A1(\cpuregs.regs[8][27] ),
    .S(_07140_),
    .X(_07148_));
 sky130_fd_sc_hd__clkbuf_1 _13245_ (.A(_07148_),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _13246_ (.A0(_07001_),
    .A1(\cpuregs.regs[8][28] ),
    .S(_07140_),
    .X(_07149_));
 sky130_fd_sc_hd__clkbuf_1 _13247_ (.A(_07149_),
    .X(_00766_));
 sky130_fd_sc_hd__mux2_1 _13248_ (.A0(_07003_),
    .A1(\cpuregs.regs[8][29] ),
    .S(_07140_),
    .X(_07150_));
 sky130_fd_sc_hd__clkbuf_1 _13249_ (.A(_07150_),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _13250_ (.A0(_07005_),
    .A1(\cpuregs.regs[8][30] ),
    .S(_07117_),
    .X(_07151_));
 sky130_fd_sc_hd__clkbuf_1 _13251_ (.A(_07151_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _13252_ (.A0(_07007_),
    .A1(\cpuregs.regs[8][31] ),
    .S(_07117_),
    .X(_07152_));
 sky130_fd_sc_hd__clkbuf_1 _13253_ (.A(_07152_),
    .X(_00769_));
 sky130_fd_sc_hd__nand2_4 _13254_ (.A(_06422_),
    .B(_06904_),
    .Y(_07153_));
 sky130_fd_sc_hd__buf_6 _13255_ (.A(_07153_),
    .X(_07154_));
 sky130_fd_sc_hd__mux2_1 _13256_ (.A0(_06941_),
    .A1(\cpuregs.regs[5][0] ),
    .S(_07154_),
    .X(_07155_));
 sky130_fd_sc_hd__clkbuf_1 _13257_ (.A(_07155_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _13258_ (.A0(_06945_),
    .A1(\cpuregs.regs[5][1] ),
    .S(_07154_),
    .X(_07156_));
 sky130_fd_sc_hd__clkbuf_1 _13259_ (.A(_07156_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _13260_ (.A0(_06947_),
    .A1(\cpuregs.regs[5][2] ),
    .S(_07154_),
    .X(_07157_));
 sky130_fd_sc_hd__clkbuf_1 _13261_ (.A(_07157_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _13262_ (.A0(_06949_),
    .A1(\cpuregs.regs[5][3] ),
    .S(_07154_),
    .X(_07158_));
 sky130_fd_sc_hd__clkbuf_1 _13263_ (.A(_07158_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _13264_ (.A0(_06951_),
    .A1(\cpuregs.regs[5][4] ),
    .S(_07154_),
    .X(_07159_));
 sky130_fd_sc_hd__clkbuf_1 _13265_ (.A(_07159_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _13266_ (.A0(_06953_),
    .A1(\cpuregs.regs[5][5] ),
    .S(_07154_),
    .X(_07160_));
 sky130_fd_sc_hd__clkbuf_1 _13267_ (.A(_07160_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _13268_ (.A0(_06955_),
    .A1(\cpuregs.regs[5][6] ),
    .S(_07154_),
    .X(_07161_));
 sky130_fd_sc_hd__clkbuf_1 _13269_ (.A(_07161_),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _13270_ (.A0(_06957_),
    .A1(\cpuregs.regs[5][7] ),
    .S(_07154_),
    .X(_07162_));
 sky130_fd_sc_hd__clkbuf_1 _13271_ (.A(_07162_),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _13272_ (.A0(_06959_),
    .A1(\cpuregs.regs[5][8] ),
    .S(_07154_),
    .X(_07163_));
 sky130_fd_sc_hd__clkbuf_1 _13273_ (.A(_07163_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _13274_ (.A0(_06961_),
    .A1(\cpuregs.regs[5][9] ),
    .S(_07154_),
    .X(_07164_));
 sky130_fd_sc_hd__clkbuf_1 _13275_ (.A(_07164_),
    .X(_00779_));
 sky130_fd_sc_hd__buf_6 _13276_ (.A(_07153_),
    .X(_07165_));
 sky130_fd_sc_hd__mux2_1 _13277_ (.A0(_06963_),
    .A1(\cpuregs.regs[5][10] ),
    .S(_07165_),
    .X(_07166_));
 sky130_fd_sc_hd__clkbuf_1 _13278_ (.A(_07166_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _13279_ (.A0(_06966_),
    .A1(\cpuregs.regs[5][11] ),
    .S(_07165_),
    .X(_07167_));
 sky130_fd_sc_hd__clkbuf_1 _13280_ (.A(_07167_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _13281_ (.A0(_06968_),
    .A1(\cpuregs.regs[5][12] ),
    .S(_07165_),
    .X(_07168_));
 sky130_fd_sc_hd__clkbuf_1 _13282_ (.A(_07168_),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _13283_ (.A0(_06970_),
    .A1(\cpuregs.regs[5][13] ),
    .S(_07165_),
    .X(_07169_));
 sky130_fd_sc_hd__clkbuf_1 _13284_ (.A(_07169_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _13285_ (.A0(_06972_),
    .A1(\cpuregs.regs[5][14] ),
    .S(_07165_),
    .X(_07170_));
 sky130_fd_sc_hd__clkbuf_1 _13286_ (.A(_07170_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _13287_ (.A0(_06974_),
    .A1(\cpuregs.regs[5][15] ),
    .S(_07165_),
    .X(_07171_));
 sky130_fd_sc_hd__clkbuf_1 _13288_ (.A(_07171_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _13289_ (.A0(_06976_),
    .A1(\cpuregs.regs[5][16] ),
    .S(_07165_),
    .X(_07172_));
 sky130_fd_sc_hd__clkbuf_1 _13290_ (.A(_07172_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _13291_ (.A0(_06978_),
    .A1(\cpuregs.regs[5][17] ),
    .S(_07165_),
    .X(_07173_));
 sky130_fd_sc_hd__clkbuf_1 _13292_ (.A(_07173_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _13293_ (.A0(_06980_),
    .A1(\cpuregs.regs[5][18] ),
    .S(_07165_),
    .X(_07174_));
 sky130_fd_sc_hd__clkbuf_1 _13294_ (.A(_07174_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _13295_ (.A0(_06982_),
    .A1(\cpuregs.regs[5][19] ),
    .S(_07165_),
    .X(_07175_));
 sky130_fd_sc_hd__clkbuf_1 _13296_ (.A(_07175_),
    .X(_00789_));
 sky130_fd_sc_hd__buf_6 _13297_ (.A(_07153_),
    .X(_07176_));
 sky130_fd_sc_hd__mux2_1 _13298_ (.A0(_06984_),
    .A1(\cpuregs.regs[5][20] ),
    .S(_07176_),
    .X(_07177_));
 sky130_fd_sc_hd__clkbuf_1 _13299_ (.A(_07177_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _13300_ (.A0(_06987_),
    .A1(\cpuregs.regs[5][21] ),
    .S(_07176_),
    .X(_07178_));
 sky130_fd_sc_hd__clkbuf_1 _13301_ (.A(_07178_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _13302_ (.A0(_06989_),
    .A1(\cpuregs.regs[5][22] ),
    .S(_07176_),
    .X(_07179_));
 sky130_fd_sc_hd__clkbuf_1 _13303_ (.A(_07179_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _13304_ (.A0(_06991_),
    .A1(\cpuregs.regs[5][23] ),
    .S(_07176_),
    .X(_07180_));
 sky130_fd_sc_hd__clkbuf_1 _13305_ (.A(_07180_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _13306_ (.A0(_06993_),
    .A1(\cpuregs.regs[5][24] ),
    .S(_07176_),
    .X(_07181_));
 sky130_fd_sc_hd__clkbuf_1 _13307_ (.A(_07181_),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _13308_ (.A0(_06995_),
    .A1(\cpuregs.regs[5][25] ),
    .S(_07176_),
    .X(_07182_));
 sky130_fd_sc_hd__clkbuf_1 _13309_ (.A(_07182_),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _13310_ (.A0(_06997_),
    .A1(\cpuregs.regs[5][26] ),
    .S(_07176_),
    .X(_07183_));
 sky130_fd_sc_hd__clkbuf_1 _13311_ (.A(_07183_),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _13312_ (.A0(_06999_),
    .A1(\cpuregs.regs[5][27] ),
    .S(_07176_),
    .X(_07184_));
 sky130_fd_sc_hd__clkbuf_1 _13313_ (.A(_07184_),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _13314_ (.A0(_07001_),
    .A1(\cpuregs.regs[5][28] ),
    .S(_07176_),
    .X(_07185_));
 sky130_fd_sc_hd__clkbuf_1 _13315_ (.A(_07185_),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _13316_ (.A0(_07003_),
    .A1(\cpuregs.regs[5][29] ),
    .S(_07176_),
    .X(_07186_));
 sky130_fd_sc_hd__clkbuf_1 _13317_ (.A(_07186_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _13318_ (.A0(_07005_),
    .A1(\cpuregs.regs[5][30] ),
    .S(_07153_),
    .X(_07187_));
 sky130_fd_sc_hd__clkbuf_1 _13319_ (.A(_07187_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _13320_ (.A0(_07007_),
    .A1(\cpuregs.regs[5][31] ),
    .S(_07153_),
    .X(_07188_));
 sky130_fd_sc_hd__clkbuf_1 _13321_ (.A(_07188_),
    .X(_00801_));
 sky130_fd_sc_hd__nor2_1 _13322_ (.A(_03312_),
    .B(_03274_),
    .Y(_07189_));
 sky130_fd_sc_hd__buf_2 _13323_ (.A(_07189_),
    .X(_07190_));
 sky130_fd_sc_hd__clkbuf_4 _13324_ (.A(_07190_),
    .X(_07191_));
 sky130_fd_sc_hd__mux4_1 _13325_ (.A0(\cpuregs.regs[28][0] ),
    .A1(\cpuregs.regs[29][0] ),
    .A2(\cpuregs.regs[30][0] ),
    .A3(\cpuregs.regs[31][0] ),
    .S0(_04282_),
    .S1(_04285_),
    .X(_07192_));
 sky130_fd_sc_hd__mux4_1 _13326_ (.A0(\cpuregs.regs[24][0] ),
    .A1(\cpuregs.regs[25][0] ),
    .A2(\cpuregs.regs[26][0] ),
    .A3(\cpuregs.regs[27][0] ),
    .S0(_04758_),
    .S1(_04759_),
    .X(_07193_));
 sky130_fd_sc_hd__mux2_1 _13327_ (.A0(_07192_),
    .A1(_07193_),
    .S(_04287_),
    .X(_07194_));
 sky130_fd_sc_hd__nand2_1 _13328_ (.A(_04272_),
    .B(_07194_),
    .Y(_07195_));
 sky130_fd_sc_hd__mux4_1 _13329_ (.A0(\cpuregs.regs[20][0] ),
    .A1(\cpuregs.regs[21][0] ),
    .A2(\cpuregs.regs[22][0] ),
    .A3(\cpuregs.regs[23][0] ),
    .S0(_04207_),
    .S1(_04208_),
    .X(_07196_));
 sky130_fd_sc_hd__mux4_1 _13330_ (.A0(\cpuregs.regs[16][0] ),
    .A1(\cpuregs.regs[17][0] ),
    .A2(\cpuregs.regs[18][0] ),
    .A3(\cpuregs.regs[19][0] ),
    .S0(_04207_),
    .S1(_04208_),
    .X(_07197_));
 sky130_fd_sc_hd__mux2_1 _13331_ (.A0(_07196_),
    .A1(_07197_),
    .S(_04211_),
    .X(_07198_));
 sky130_fd_sc_hd__a21oi_1 _13332_ (.A1(_04215_),
    .A2(_07198_),
    .B1(_04225_),
    .Y(_07199_));
 sky130_fd_sc_hd__mux4_1 _13333_ (.A0(\cpuregs.regs[4][0] ),
    .A1(\cpuregs.regs[5][0] ),
    .A2(\cpuregs.regs[6][0] ),
    .A3(\cpuregs.regs[7][0] ),
    .S0(_04758_),
    .S1(_04759_),
    .X(_07200_));
 sky130_fd_sc_hd__mux4_1 _13334_ (.A0(\cpuregs.regs[0][0] ),
    .A1(\cpuregs.regs[1][0] ),
    .A2(\cpuregs.regs[2][0] ),
    .A3(\cpuregs.regs[3][0] ),
    .S0(_04758_),
    .S1(_04759_),
    .X(_07201_));
 sky130_fd_sc_hd__mux2_1 _13335_ (.A0(_07200_),
    .A1(_07201_),
    .S(_04211_),
    .X(_07202_));
 sky130_fd_sc_hd__mux4_1 _13336_ (.A0(\cpuregs.regs[12][0] ),
    .A1(\cpuregs.regs[13][0] ),
    .A2(\cpuregs.regs[14][0] ),
    .A3(\cpuregs.regs[15][0] ),
    .S0(_04579_),
    .S1(_04284_),
    .X(_07203_));
 sky130_fd_sc_hd__mux4_1 _13337_ (.A0(\cpuregs.regs[8][0] ),
    .A1(\cpuregs.regs[9][0] ),
    .A2(\cpuregs.regs[10][0] ),
    .A3(\cpuregs.regs[11][0] ),
    .S0(_04579_),
    .S1(_04284_),
    .X(_07204_));
 sky130_fd_sc_hd__mux2_1 _13338_ (.A0(_07203_),
    .A1(_07204_),
    .S(_04575_),
    .X(_07205_));
 sky130_fd_sc_hd__a21o_1 _13339_ (.A1(_04054_),
    .A2(_07205_),
    .B1(_04296_),
    .X(_07206_));
 sky130_fd_sc_hd__a21oi_1 _13340_ (.A1(_04215_),
    .A2(_07202_),
    .B1(_07206_),
    .Y(_07207_));
 sky130_fd_sc_hd__a211o_4 _13341_ (.A1(_07195_),
    .A2(_07199_),
    .B1(_04227_),
    .C1(_07207_),
    .X(_07208_));
 sky130_fd_sc_hd__clkinv_4 _13342_ (.A(is_lui_auipc_jal),
    .Y(_07209_));
 sky130_fd_sc_hd__nor2_2 _13343_ (.A(instr_lui),
    .B(_07209_),
    .Y(_07210_));
 sky130_fd_sc_hd__clkbuf_4 _13344_ (.A(_07210_),
    .X(_07211_));
 sky130_fd_sc_hd__a2bb2o_1 _13345_ (.A1_N(_03387_),
    .A2_N(_07208_),
    .B1(_07211_),
    .B2(\reg_next_pc[0] ),
    .X(_07212_));
 sky130_fd_sc_hd__a21oi_1 _13346_ (.A1(_04037_),
    .A2(\decoded_imm[0] ),
    .B1(_03311_),
    .Y(_07213_));
 sky130_fd_sc_hd__o21a_1 _13347_ (.A1(_04037_),
    .A2(\decoded_imm[0] ),
    .B1(_07213_),
    .X(_07214_));
 sky130_fd_sc_hd__and2_1 _13348_ (.A(\cpu_state[4] ),
    .B(_03399_),
    .X(_07215_));
 sky130_fd_sc_hd__clkbuf_4 _13349_ (.A(_07215_),
    .X(_07216_));
 sky130_fd_sc_hd__clkbuf_4 _13350_ (.A(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__o221a_1 _13351_ (.A1(_04251_),
    .A2(_03313_),
    .B1(_07217_),
    .B2(_04118_),
    .C1(_05260_),
    .X(_07218_));
 sky130_fd_sc_hd__a211o_1 _13352_ (.A1(_07191_),
    .A2(_07212_),
    .B1(_07214_),
    .C1(_07218_),
    .X(_07219_));
 sky130_fd_sc_hd__or2_1 _13353_ (.A(\cpu_state[4] ),
    .B(_03274_),
    .X(_07220_));
 sky130_fd_sc_hd__clkbuf_4 _13354_ (.A(_07220_),
    .X(_07221_));
 sky130_fd_sc_hd__o22a_1 _13355_ (.A1(\cpu_state[2] ),
    .A2(_07221_),
    .B1(_05211_),
    .B2(_03400_),
    .X(_07222_));
 sky130_fd_sc_hd__and3b_1 _13356_ (.A_N(_03316_),
    .B(_07222_),
    .C(_03281_),
    .X(_07223_));
 sky130_fd_sc_hd__buf_4 _13357_ (.A(_07223_),
    .X(_07224_));
 sky130_fd_sc_hd__buf_4 _13358_ (.A(_07224_),
    .X(_07225_));
 sky130_fd_sc_hd__mux2_1 _13359_ (.A0(_04037_),
    .A1(_07219_),
    .S(_07225_),
    .X(_07226_));
 sky130_fd_sc_hd__clkbuf_1 _13360_ (.A(_07226_),
    .X(_00802_));
 sky130_fd_sc_hd__nand2_1 _13361_ (.A(_04040_),
    .B(\decoded_imm[1] ),
    .Y(_07227_));
 sky130_fd_sc_hd__or2_1 _13362_ (.A(net78),
    .B(\decoded_imm[1] ),
    .X(_07228_));
 sky130_fd_sc_hd__and4_1 _13363_ (.A(_04036_),
    .B(\decoded_imm[0] ),
    .C(_07227_),
    .D(_07228_),
    .X(_07229_));
 sky130_fd_sc_hd__inv_2 _13364_ (.A(_07229_),
    .Y(_07230_));
 sky130_fd_sc_hd__a22o_1 _13365_ (.A1(_04037_),
    .A2(\decoded_imm[0] ),
    .B1(_07227_),
    .B2(_07228_),
    .X(_07231_));
 sky130_fd_sc_hd__clkbuf_4 _13366_ (.A(_07189_),
    .X(_07232_));
 sky130_fd_sc_hd__a2bb2o_1 _13367_ (.A1_N(_03387_),
    .A2_N(_04101_),
    .B1(_07210_),
    .B2(\reg_pc[1] ),
    .X(_07233_));
 sky130_fd_sc_hd__mux2_1 _13368_ (.A0(_04036_),
    .A1(_04160_),
    .S(_05257_),
    .X(_07234_));
 sky130_fd_sc_hd__or2_1 _13369_ (.A(_03399_),
    .B(_07234_),
    .X(_07235_));
 sky130_fd_sc_hd__clkbuf_4 _13370_ (.A(_05258_),
    .X(_07236_));
 sky130_fd_sc_hd__and2_1 _13371_ (.A(\cpu_state[4] ),
    .B(_03313_),
    .X(_07237_));
 sky130_fd_sc_hd__clkbuf_4 _13372_ (.A(_07237_),
    .X(_07238_));
 sky130_fd_sc_hd__a31o_1 _13373_ (.A1(_03312_),
    .A2(_04262_),
    .A3(_07236_),
    .B1(_07238_),
    .X(_07239_));
 sky130_fd_sc_hd__a22o_1 _13374_ (.A1(_07232_),
    .A2(_07233_),
    .B1(_07235_),
    .B2(_07239_),
    .X(_07240_));
 sky130_fd_sc_hd__a31o_1 _13375_ (.A1(_03276_),
    .A2(_07230_),
    .A3(_07231_),
    .B1(_07240_),
    .X(_07241_));
 sky130_fd_sc_hd__mux2_1 _13376_ (.A0(_04040_),
    .A1(_07241_),
    .S(_07225_),
    .X(_07242_));
 sky130_fd_sc_hd__clkbuf_1 _13377_ (.A(_07242_),
    .X(_00803_));
 sky130_fd_sc_hd__nand2_1 _13378_ (.A(net89),
    .B(\decoded_imm[2] ),
    .Y(_07243_));
 sky130_fd_sc_hd__or2_1 _13379_ (.A(net89),
    .B(\decoded_imm[2] ),
    .X(_07244_));
 sky130_fd_sc_hd__and2_1 _13380_ (.A(net78),
    .B(\decoded_imm[1] ),
    .X(_07245_));
 sky130_fd_sc_hd__a31o_1 _13381_ (.A1(net67),
    .A2(\decoded_imm[0] ),
    .A3(_07228_),
    .B1(_07245_),
    .X(_07246_));
 sky130_fd_sc_hd__and3_1 _13382_ (.A(_07243_),
    .B(_07244_),
    .C(_07246_),
    .X(_07247_));
 sky130_fd_sc_hd__inv_2 _13383_ (.A(_07247_),
    .Y(_07248_));
 sky130_fd_sc_hd__a21o_1 _13384_ (.A1(_07243_),
    .A2(_07244_),
    .B1(_07246_),
    .X(_07249_));
 sky130_fd_sc_hd__inv_2 _13385_ (.A(_04142_),
    .Y(_07250_));
 sky130_fd_sc_hd__a22o_1 _13386_ (.A1(_07209_),
    .A2(_07250_),
    .B1(_07211_),
    .B2(\reg_pc[2] ),
    .X(_07251_));
 sky130_fd_sc_hd__mux2_1 _13387_ (.A0(_04039_),
    .A1(_04198_),
    .S(_05257_),
    .X(_07252_));
 sky130_fd_sc_hd__or2_1 _13388_ (.A(_03399_),
    .B(_07252_),
    .X(_07253_));
 sky130_fd_sc_hd__clkbuf_4 _13389_ (.A(_07237_),
    .X(_07254_));
 sky130_fd_sc_hd__a31o_1 _13390_ (.A1(_03312_),
    .A2(_04342_),
    .A3(_05259_),
    .B1(_07254_),
    .X(_07255_));
 sky130_fd_sc_hd__a22o_1 _13391_ (.A1(_07232_),
    .A2(_07251_),
    .B1(_07253_),
    .B2(_07255_),
    .X(_07256_));
 sky130_fd_sc_hd__a31o_1 _13392_ (.A1(_03276_),
    .A2(_07248_),
    .A3(_07249_),
    .B1(_07256_),
    .X(_07257_));
 sky130_fd_sc_hd__mux2_1 _13393_ (.A0(_04160_),
    .A1(_07257_),
    .S(_07225_),
    .X(_07258_));
 sky130_fd_sc_hd__clkbuf_1 _13394_ (.A(_07258_),
    .X(_00804_));
 sky130_fd_sc_hd__nand2_1 _13395_ (.A(net92),
    .B(\decoded_imm[3] ),
    .Y(_07259_));
 sky130_fd_sc_hd__or2_1 _13396_ (.A(net92),
    .B(\decoded_imm[3] ),
    .X(_07260_));
 sky130_fd_sc_hd__a21bo_1 _13397_ (.A1(_07244_),
    .A2(_07246_),
    .B1_N(_07243_),
    .X(_07261_));
 sky130_fd_sc_hd__nand3_1 _13398_ (.A(_07259_),
    .B(_07260_),
    .C(_07261_),
    .Y(_07262_));
 sky130_fd_sc_hd__a21o_1 _13399_ (.A1(_07259_),
    .A2(_07260_),
    .B1(_07261_),
    .X(_07263_));
 sky130_fd_sc_hd__a22o_1 _13400_ (.A1(_07209_),
    .A2(_04186_),
    .B1(_07210_),
    .B2(\reg_pc[3] ),
    .X(_07264_));
 sky130_fd_sc_hd__mux2_1 _13401_ (.A0(_04160_),
    .A1(_04251_),
    .S(_05257_),
    .X(_07265_));
 sky130_fd_sc_hd__or2_1 _13402_ (.A(_03399_),
    .B(_07265_),
    .X(_07266_));
 sky130_fd_sc_hd__a31o_1 _13403_ (.A1(_03312_),
    .A2(_04360_),
    .A3(_05259_),
    .B1(_07254_),
    .X(_07267_));
 sky130_fd_sc_hd__a22o_1 _13404_ (.A1(_07232_),
    .A2(_07264_),
    .B1(_07266_),
    .B2(_07267_),
    .X(_07268_));
 sky130_fd_sc_hd__a31o_1 _13405_ (.A1(_03276_),
    .A2(_07262_),
    .A3(_07263_),
    .B1(_07268_),
    .X(_07269_));
 sky130_fd_sc_hd__mux2_1 _13406_ (.A0(_04198_),
    .A1(_07269_),
    .S(_07225_),
    .X(_07270_));
 sky130_fd_sc_hd__clkbuf_1 _13407_ (.A(_07270_),
    .X(_00805_));
 sky130_fd_sc_hd__clkbuf_4 _13408_ (.A(_07224_),
    .X(_07271_));
 sky130_fd_sc_hd__inv_2 _13409_ (.A(_04419_),
    .Y(_07272_));
 sky130_fd_sc_hd__nand2_1 _13410_ (.A(_07272_),
    .B(_07236_),
    .Y(_07273_));
 sky130_fd_sc_hd__clkbuf_4 _13411_ (.A(_07216_),
    .X(_07274_));
 sky130_fd_sc_hd__o211a_1 _13412_ (.A1(_04037_),
    .A2(_05260_),
    .B1(_07273_),
    .C1(_07274_),
    .X(_07275_));
 sky130_fd_sc_hd__buf_2 _13413_ (.A(_05209_),
    .X(_07276_));
 sky130_fd_sc_hd__buf_2 _13414_ (.A(_07276_),
    .X(_07277_));
 sky130_fd_sc_hd__or2_1 _13415_ (.A(_04198_),
    .B(_05258_),
    .X(_07278_));
 sky130_fd_sc_hd__buf_2 _13416_ (.A(_07238_),
    .X(_07279_));
 sky130_fd_sc_hd__o211a_1 _13417_ (.A1(_04262_),
    .A2(_07277_),
    .B1(_07278_),
    .C1(_07279_),
    .X(_07280_));
 sky130_fd_sc_hd__clkbuf_4 _13418_ (.A(_07209_),
    .X(_07281_));
 sky130_fd_sc_hd__clkbuf_4 _13419_ (.A(_07211_),
    .X(_07282_));
 sky130_fd_sc_hd__clkbuf_4 _13420_ (.A(_07221_),
    .X(_07283_));
 sky130_fd_sc_hd__clkbuf_4 _13421_ (.A(_07283_),
    .X(_07284_));
 sky130_fd_sc_hd__a221o_1 _13422_ (.A1(_07281_),
    .A2(_04241_),
    .B1(_07282_),
    .B2(\reg_pc[4] ),
    .C1(_07284_),
    .X(_07285_));
 sky130_fd_sc_hd__o31a_1 _13423_ (.A1(_07191_),
    .A2(_07275_),
    .A3(_07280_),
    .B1(_07285_),
    .X(_07286_));
 sky130_fd_sc_hd__and2_1 _13424_ (.A(net93),
    .B(\decoded_imm[4] ),
    .X(_07287_));
 sky130_fd_sc_hd__nor2_1 _13425_ (.A(net93),
    .B(\decoded_imm[4] ),
    .Y(_07288_));
 sky130_fd_sc_hd__a21bo_1 _13426_ (.A1(_07260_),
    .A2(_07261_),
    .B1_N(_07259_),
    .X(_07289_));
 sky130_fd_sc_hd__o21ba_1 _13427_ (.A1(_07287_),
    .A2(_07288_),
    .B1_N(_07289_),
    .X(_07290_));
 sky130_fd_sc_hd__inv_2 _13428_ (.A(_07288_),
    .Y(_07291_));
 sky130_fd_sc_hd__and3b_1 _13429_ (.A_N(_07287_),
    .B(_07291_),
    .C(_07289_),
    .X(_07292_));
 sky130_fd_sc_hd__o31ai_1 _13430_ (.A1(_03631_),
    .A2(_07290_),
    .A3(_07292_),
    .B1(_07271_),
    .Y(_07293_));
 sky130_fd_sc_hd__o22a_1 _13431_ (.A1(_04251_),
    .A2(_07271_),
    .B1(_07286_),
    .B2(_07293_),
    .X(_00806_));
 sky130_fd_sc_hd__or2_1 _13432_ (.A(_04251_),
    .B(_05259_),
    .X(_07294_));
 sky130_fd_sc_hd__o211a_1 _13433_ (.A1(_04342_),
    .A2(_07277_),
    .B1(_07294_),
    .C1(_07279_),
    .X(_07295_));
 sky130_fd_sc_hd__or2_1 _13434_ (.A(_07287_),
    .B(_07292_),
    .X(_07296_));
 sky130_fd_sc_hd__or2_2 _13435_ (.A(_03524_),
    .B(\decoded_imm[5] ),
    .X(_07297_));
 sky130_fd_sc_hd__nand2_1 _13436_ (.A(_04262_),
    .B(\decoded_imm[5] ),
    .Y(_07298_));
 sky130_fd_sc_hd__nand3_1 _13437_ (.A(_07296_),
    .B(_07297_),
    .C(_07298_),
    .Y(_07299_));
 sky130_fd_sc_hd__a21o_1 _13438_ (.A1(_07297_),
    .A2(_07298_),
    .B1(_07296_),
    .X(_07300_));
 sky130_fd_sc_hd__or2_1 _13439_ (.A(_04456_),
    .B(_07276_),
    .X(_07301_));
 sky130_fd_sc_hd__o211a_1 _13440_ (.A1(_04040_),
    .A2(_05259_),
    .B1(_07301_),
    .C1(_07216_),
    .X(_07302_));
 sky130_fd_sc_hd__a31o_1 _13441_ (.A1(_03275_),
    .A2(_07299_),
    .A3(_07300_),
    .B1(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__clkbuf_4 _13442_ (.A(_07209_),
    .X(_07304_));
 sky130_fd_sc_hd__clkbuf_4 _13443_ (.A(_07211_),
    .X(_07305_));
 sky130_fd_sc_hd__a221o_1 _13444_ (.A1(_07304_),
    .A2(_04307_),
    .B1(_07305_),
    .B2(\reg_pc[5] ),
    .C1(_07283_),
    .X(_07306_));
 sky130_fd_sc_hd__o31a_1 _13445_ (.A1(_07191_),
    .A2(_07295_),
    .A3(_07303_),
    .B1(_07306_),
    .X(_07307_));
 sky130_fd_sc_hd__mux2_1 _13446_ (.A0(_04262_),
    .A1(_07307_),
    .S(_07225_),
    .X(_07308_));
 sky130_fd_sc_hd__clkbuf_1 _13447_ (.A(_07308_),
    .X(_00807_));
 sky130_fd_sc_hd__a221o_1 _13448_ (.A1(_03524_),
    .A2(\decoded_imm[5] ),
    .B1(_07291_),
    .B2(_07289_),
    .C1(_07287_),
    .X(_07309_));
 sky130_fd_sc_hd__nand2_1 _13449_ (.A(net95),
    .B(\decoded_imm[6] ),
    .Y(_07310_));
 sky130_fd_sc_hd__or2_1 _13450_ (.A(net95),
    .B(\decoded_imm[6] ),
    .X(_07311_));
 sky130_fd_sc_hd__and2_1 _13451_ (.A(_07310_),
    .B(_07311_),
    .X(_07312_));
 sky130_fd_sc_hd__a21oi_1 _13452_ (.A1(_07297_),
    .A2(_07309_),
    .B1(_07312_),
    .Y(_07313_));
 sky130_fd_sc_hd__a31o_1 _13453_ (.A1(_07297_),
    .A2(_07312_),
    .A3(_07309_),
    .B1(_03631_),
    .X(_07314_));
 sky130_fd_sc_hd__clkbuf_4 _13454_ (.A(_05257_),
    .X(_07315_));
 sky130_fd_sc_hd__or2_1 _13455_ (.A(_04466_),
    .B(_05209_),
    .X(_07316_));
 sky130_fd_sc_hd__o211a_1 _13456_ (.A1(_04160_),
    .A2(_07315_),
    .B1(_07316_),
    .C1(_07216_),
    .X(_07317_));
 sky130_fd_sc_hd__or2_1 _13457_ (.A(_04262_),
    .B(_05257_),
    .X(_07318_));
 sky130_fd_sc_hd__o211a_1 _13458_ (.A1(_04360_),
    .A2(_05227_),
    .B1(_07318_),
    .C1(_07237_),
    .X(_07319_));
 sky130_fd_sc_hd__or3_1 _13459_ (.A(_07190_),
    .B(_07317_),
    .C(_07319_),
    .X(_07320_));
 sky130_fd_sc_hd__nor2_1 _13460_ (.A(_03387_),
    .B(_04335_),
    .Y(_07321_));
 sky130_fd_sc_hd__a211o_1 _13461_ (.A1(\reg_pc[6] ),
    .A2(_07211_),
    .B1(_07321_),
    .C1(_07221_),
    .X(_07322_));
 sky130_fd_sc_hd__a2bb2o_1 _13462_ (.A1_N(_07313_),
    .A2_N(_07314_),
    .B1(_07320_),
    .B2(_07322_),
    .X(_07323_));
 sky130_fd_sc_hd__mux2_1 _13463_ (.A0(_04342_),
    .A1(_07323_),
    .S(_07225_),
    .X(_07324_));
 sky130_fd_sc_hd__clkbuf_1 _13464_ (.A(_07324_),
    .X(_00808_));
 sky130_fd_sc_hd__and2_1 _13465_ (.A(_03518_),
    .B(\decoded_imm[7] ),
    .X(_07325_));
 sky130_fd_sc_hd__nor2_1 _13466_ (.A(_04360_),
    .B(\decoded_imm[7] ),
    .Y(_07326_));
 sky130_fd_sc_hd__inv_2 _13467_ (.A(_07310_),
    .Y(_07327_));
 sky130_fd_sc_hd__a31o_1 _13468_ (.A1(_07297_),
    .A2(_07311_),
    .A3(_07309_),
    .B1(_07327_),
    .X(_07328_));
 sky130_fd_sc_hd__or3b_1 _13469_ (.A(_07325_),
    .B(_07326_),
    .C_N(_07328_),
    .X(_07329_));
 sky130_fd_sc_hd__o21bai_1 _13470_ (.A1(_07325_),
    .A2(_07326_),
    .B1_N(_07328_),
    .Y(_07330_));
 sky130_fd_sc_hd__or2_1 _13471_ (.A(_04342_),
    .B(_05259_),
    .X(_07331_));
 sky130_fd_sc_hd__or2_1 _13472_ (.A(_04532_),
    .B(_07276_),
    .X(_07332_));
 sky130_fd_sc_hd__a31o_1 _13473_ (.A1(_07217_),
    .A2(_07278_),
    .A3(_07332_),
    .B1(_07189_),
    .X(_07333_));
 sky130_fd_sc_hd__a31o_1 _13474_ (.A1(_07279_),
    .A2(_07273_),
    .A3(_07331_),
    .B1(_07333_),
    .X(_07334_));
 sky130_fd_sc_hd__nor2_1 _13475_ (.A(_03387_),
    .B(_04382_),
    .Y(_07335_));
 sky130_fd_sc_hd__a211o_1 _13476_ (.A1(\reg_pc[7] ),
    .A2(_07305_),
    .B1(_07335_),
    .C1(_07221_),
    .X(_07336_));
 sky130_fd_sc_hd__a32o_1 _13477_ (.A1(_03275_),
    .A2(_07329_),
    .A3(_07330_),
    .B1(_07334_),
    .B2(_07336_),
    .X(_07337_));
 sky130_fd_sc_hd__mux2_1 _13478_ (.A0(_04360_),
    .A1(_07337_),
    .S(_07225_),
    .X(_07338_));
 sky130_fd_sc_hd__clkbuf_1 _13479_ (.A(_07338_),
    .X(_00809_));
 sky130_fd_sc_hd__or2_1 _13480_ (.A(_04566_),
    .B(_07276_),
    .X(_07339_));
 sky130_fd_sc_hd__o211a_1 _13481_ (.A1(_04360_),
    .A2(_05260_),
    .B1(_07301_),
    .C1(_07279_),
    .X(_07340_));
 sky130_fd_sc_hd__a31o_1 _13482_ (.A1(_07274_),
    .A2(_07294_),
    .A3(_07339_),
    .B1(_07340_),
    .X(_07341_));
 sky130_fd_sc_hd__a221o_1 _13483_ (.A1(_07281_),
    .A2(_04415_),
    .B1(_07282_),
    .B2(\reg_pc[8] ),
    .C1(_07284_),
    .X(_07342_));
 sky130_fd_sc_hd__o21a_1 _13484_ (.A1(_07191_),
    .A2(_07341_),
    .B1(_07342_),
    .X(_07343_));
 sky130_fd_sc_hd__or2_1 _13485_ (.A(net96),
    .B(\decoded_imm[7] ),
    .X(_07344_));
 sky130_fd_sc_hd__a21oi_2 _13486_ (.A1(_07344_),
    .A2(_07328_),
    .B1(_07325_),
    .Y(_07345_));
 sky130_fd_sc_hd__xnor2_1 _13487_ (.A(_03510_),
    .B(\decoded_imm[8] ),
    .Y(_07346_));
 sky130_fd_sc_hd__nor2_1 _13488_ (.A(_07345_),
    .B(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__a21o_1 _13489_ (.A1(_07345_),
    .A2(_07346_),
    .B1(_03631_),
    .X(_07348_));
 sky130_fd_sc_hd__o21ai_1 _13490_ (.A1(_07347_),
    .A2(_07348_),
    .B1(_07271_),
    .Y(_07349_));
 sky130_fd_sc_hd__o22a_1 _13491_ (.A1(_04419_),
    .A2(_07271_),
    .B1(_07343_),
    .B2(_07349_),
    .X(_00810_));
 sky130_fd_sc_hd__and2_1 _13492_ (.A(net98),
    .B(\decoded_imm[9] ),
    .X(_07350_));
 sky130_fd_sc_hd__nor2_1 _13493_ (.A(net98),
    .B(\decoded_imm[9] ),
    .Y(_07351_));
 sky130_fd_sc_hd__nor2_1 _13494_ (.A(_07350_),
    .B(_07351_),
    .Y(_07352_));
 sky130_fd_sc_hd__a21o_1 _13495_ (.A1(_03510_),
    .A2(\decoded_imm[8] ),
    .B1(_07347_),
    .X(_07353_));
 sky130_fd_sc_hd__or2_1 _13496_ (.A(_07352_),
    .B(_07353_),
    .X(_07354_));
 sky130_fd_sc_hd__nand2_1 _13497_ (.A(_07352_),
    .B(_07353_),
    .Y(_07355_));
 sky130_fd_sc_hd__and3_1 _13498_ (.A(_03275_),
    .B(_07354_),
    .C(_07355_),
    .X(_07356_));
 sky130_fd_sc_hd__o211a_1 _13499_ (.A1(_04419_),
    .A2(_05260_),
    .B1(_07316_),
    .C1(_07279_),
    .X(_07357_));
 sky130_fd_sc_hd__or2_1 _13500_ (.A(_04602_),
    .B(_07276_),
    .X(_07358_));
 sky130_fd_sc_hd__a31o_1 _13501_ (.A1(_07274_),
    .A2(_07318_),
    .A3(_07358_),
    .B1(_07232_),
    .X(_07359_));
 sky130_fd_sc_hd__a221o_1 _13502_ (.A1(_07304_),
    .A2(_04447_),
    .B1(_07305_),
    .B2(\reg_pc[9] ),
    .C1(_07283_),
    .X(_07360_));
 sky130_fd_sc_hd__o31a_1 _13503_ (.A1(_07356_),
    .A2(_07357_),
    .A3(_07359_),
    .B1(_07360_),
    .X(_07361_));
 sky130_fd_sc_hd__mux2_1 _13504_ (.A0(_04456_),
    .A1(_07361_),
    .S(_07225_),
    .X(_07362_));
 sky130_fd_sc_hd__clkbuf_1 _13505_ (.A(_07362_),
    .X(_00811_));
 sky130_fd_sc_hd__nand2_1 _13506_ (.A(_04456_),
    .B(\decoded_imm[9] ),
    .Y(_07363_));
 sky130_fd_sc_hd__xnor2_1 _13507_ (.A(net68),
    .B(\decoded_imm[10] ),
    .Y(_07364_));
 sky130_fd_sc_hd__a21oi_1 _13508_ (.A1(_07363_),
    .A2(_07355_),
    .B1(_07364_),
    .Y(_07365_));
 sky130_fd_sc_hd__a31o_1 _13509_ (.A1(_07363_),
    .A2(_07355_),
    .A3(_07364_),
    .B1(_03311_),
    .X(_07366_));
 sky130_fd_sc_hd__nor2_1 _13510_ (.A(_07365_),
    .B(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__mux2_1 _13511_ (.A0(_04342_),
    .A1(_04611_),
    .S(_07315_),
    .X(_07368_));
 sky130_fd_sc_hd__o211a_1 _13512_ (.A1(_04456_),
    .A2(_05259_),
    .B1(_07332_),
    .C1(_07254_),
    .X(_07369_));
 sky130_fd_sc_hd__a211o_1 _13513_ (.A1(_07274_),
    .A2(_07368_),
    .B1(_07369_),
    .C1(_07190_),
    .X(_07370_));
 sky130_fd_sc_hd__inv_2 _13514_ (.A(_04493_),
    .Y(_07371_));
 sky130_fd_sc_hd__a22o_1 _13515_ (.A1(_07281_),
    .A2(_07371_),
    .B1(_07282_),
    .B2(\reg_pc[10] ),
    .X(_07372_));
 sky130_fd_sc_hd__o22a_1 _13516_ (.A1(_07367_),
    .A2(_07370_),
    .B1(_07372_),
    .B2(_07284_),
    .X(_07373_));
 sky130_fd_sc_hd__buf_4 _13517_ (.A(_07223_),
    .X(_07374_));
 sky130_fd_sc_hd__mux2_1 _13518_ (.A0(_04466_),
    .A1(_07373_),
    .S(_07374_),
    .X(_07375_));
 sky130_fd_sc_hd__clkbuf_1 _13519_ (.A(_07375_),
    .X(_00812_));
 sky130_fd_sc_hd__nand2_1 _13520_ (.A(net69),
    .B(\decoded_imm[11] ),
    .Y(_07376_));
 sky130_fd_sc_hd__or2_1 _13521_ (.A(net69),
    .B(\decoded_imm[11] ),
    .X(_07377_));
 sky130_fd_sc_hd__nand2_1 _13522_ (.A(_07376_),
    .B(_07377_),
    .Y(_07378_));
 sky130_fd_sc_hd__a21o_1 _13523_ (.A1(_04466_),
    .A2(\decoded_imm[10] ),
    .B1(_07365_),
    .X(_07379_));
 sky130_fd_sc_hd__xnor2_1 _13524_ (.A(_07378_),
    .B(_07379_),
    .Y(_07380_));
 sky130_fd_sc_hd__o211a_1 _13525_ (.A1(_04466_),
    .A2(_07315_),
    .B1(_07339_),
    .C1(_07254_),
    .X(_07381_));
 sky130_fd_sc_hd__or2_1 _13526_ (.A(_04642_),
    .B(_07276_),
    .X(_07382_));
 sky130_fd_sc_hd__o211a_1 _13527_ (.A1(_04360_),
    .A2(_07315_),
    .B1(_07382_),
    .C1(_07216_),
    .X(_07383_));
 sky130_fd_sc_hd__or3_1 _13528_ (.A(_07190_),
    .B(_07381_),
    .C(_07383_),
    .X(_07384_));
 sky130_fd_sc_hd__a221o_1 _13529_ (.A1(_07304_),
    .A2(_04526_),
    .B1(_07211_),
    .B2(\reg_pc[11] ),
    .C1(_07221_),
    .X(_07385_));
 sky130_fd_sc_hd__a22o_1 _13530_ (.A1(_03276_),
    .A2(_07380_),
    .B1(_07384_),
    .B2(_07385_),
    .X(_07386_));
 sky130_fd_sc_hd__mux2_1 _13531_ (.A0(_04532_),
    .A1(_07386_),
    .S(_07374_),
    .X(_07387_));
 sky130_fd_sc_hd__clkbuf_1 _13532_ (.A(_07387_),
    .X(_00813_));
 sky130_fd_sc_hd__o211a_1 _13533_ (.A1(_04532_),
    .A2(_07315_),
    .B1(_07358_),
    .C1(_07254_),
    .X(_07388_));
 sky130_fd_sc_hd__or2_1 _13534_ (.A(_04708_),
    .B(_07276_),
    .X(_07389_));
 sky130_fd_sc_hd__o211a_1 _13535_ (.A1(_04419_),
    .A2(_07315_),
    .B1(_07389_),
    .C1(_07216_),
    .X(_07390_));
 sky130_fd_sc_hd__or3_1 _13536_ (.A(_07190_),
    .B(_07388_),
    .C(_07390_),
    .X(_07391_));
 sky130_fd_sc_hd__a221o_1 _13537_ (.A1(_07209_),
    .A2(_04562_),
    .B1(_07211_),
    .B2(\reg_pc[12] ),
    .C1(_07221_),
    .X(_07392_));
 sky130_fd_sc_hd__nor2_1 _13538_ (.A(_07364_),
    .B(_07378_),
    .Y(_07393_));
 sky130_fd_sc_hd__or4bb_1 _13539_ (.A(_07345_),
    .B(_07346_),
    .C_N(_07352_),
    .D_N(_07393_),
    .X(_07394_));
 sky130_fd_sc_hd__a31o_1 _13540_ (.A1(_03510_),
    .A2(\decoded_imm[8] ),
    .A3(_07352_),
    .B1(_07350_),
    .X(_07395_));
 sky130_fd_sc_hd__and3_1 _13541_ (.A(net68),
    .B(\decoded_imm[10] ),
    .C(_07377_),
    .X(_07396_));
 sky130_fd_sc_hd__a221oi_2 _13542_ (.A1(net69),
    .A2(\decoded_imm[11] ),
    .B1(_07393_),
    .B2(_07395_),
    .C1(_07396_),
    .Y(_07397_));
 sky130_fd_sc_hd__nand2_1 _13543_ (.A(net70),
    .B(\decoded_imm[12] ),
    .Y(_07398_));
 sky130_fd_sc_hd__or2_1 _13544_ (.A(net70),
    .B(\decoded_imm[12] ),
    .X(_07399_));
 sky130_fd_sc_hd__nand2_1 _13545_ (.A(_07398_),
    .B(_07399_),
    .Y(_07400_));
 sky130_fd_sc_hd__a21o_1 _13546_ (.A1(_07394_),
    .A2(_07397_),
    .B1(_07400_),
    .X(_07401_));
 sky130_fd_sc_hd__a31oi_1 _13547_ (.A1(_07394_),
    .A2(_07397_),
    .A3(_07400_),
    .B1(_03631_),
    .Y(_07402_));
 sky130_fd_sc_hd__a22o_1 _13548_ (.A1(_07391_),
    .A2(_07392_),
    .B1(_07401_),
    .B2(_07402_),
    .X(_07403_));
 sky130_fd_sc_hd__mux2_1 _13549_ (.A0(_04566_),
    .A1(_07403_),
    .S(_07374_),
    .X(_07404_));
 sky130_fd_sc_hd__clkbuf_1 _13550_ (.A(_07404_),
    .X(_00814_));
 sky130_fd_sc_hd__a22o_1 _13551_ (.A1(_07281_),
    .A2(_04593_),
    .B1(_07282_),
    .B2(\reg_pc[13] ),
    .X(_07405_));
 sky130_fd_sc_hd__or2_1 _13552_ (.A(net71),
    .B(\decoded_imm[13] ),
    .X(_07406_));
 sky130_fd_sc_hd__nand2_1 _13553_ (.A(net71),
    .B(\decoded_imm[13] ),
    .Y(_07407_));
 sky130_fd_sc_hd__nand2_1 _13554_ (.A(_07406_),
    .B(_07407_),
    .Y(_07408_));
 sky130_fd_sc_hd__nand2_1 _13555_ (.A(_07398_),
    .B(_07401_),
    .Y(_07409_));
 sky130_fd_sc_hd__xnor2_1 _13556_ (.A(_07408_),
    .B(_07409_),
    .Y(_07410_));
 sky130_fd_sc_hd__mux2_1 _13557_ (.A0(_04611_),
    .A1(_04566_),
    .S(_05227_),
    .X(_07411_));
 sky130_fd_sc_hd__nand2_1 _13558_ (.A(_03566_),
    .B(_05258_),
    .Y(_07412_));
 sky130_fd_sc_hd__o211a_1 _13559_ (.A1(_04456_),
    .A2(_05258_),
    .B1(_07412_),
    .C1(_07216_),
    .X(_07413_));
 sky130_fd_sc_hd__a211o_1 _13560_ (.A1(_07238_),
    .A2(_07411_),
    .B1(_07413_),
    .C1(_07190_),
    .X(_07414_));
 sky130_fd_sc_hd__a21o_1 _13561_ (.A1(_03275_),
    .A2(_07410_),
    .B1(_07414_),
    .X(_07415_));
 sky130_fd_sc_hd__o21a_1 _13562_ (.A1(_07284_),
    .A2(_07405_),
    .B1(_07415_),
    .X(_07416_));
 sky130_fd_sc_hd__mux2_1 _13563_ (.A0(_04602_),
    .A1(_07416_),
    .S(_07374_),
    .X(_07417_));
 sky130_fd_sc_hd__clkbuf_1 _13564_ (.A(_07417_),
    .X(_00815_));
 sky130_fd_sc_hd__nand2_1 _13565_ (.A(net72),
    .B(\decoded_imm[14] ),
    .Y(_07418_));
 sky130_fd_sc_hd__or2_1 _13566_ (.A(net72),
    .B(\decoded_imm[14] ),
    .X(_07419_));
 sky130_fd_sc_hd__and2_1 _13567_ (.A(_07418_),
    .B(_07419_),
    .X(_07420_));
 sky130_fd_sc_hd__a21bo_1 _13568_ (.A1(_07406_),
    .A2(_07409_),
    .B1_N(_07407_),
    .X(_07421_));
 sky130_fd_sc_hd__nand2_1 _13569_ (.A(_07420_),
    .B(_07421_),
    .Y(_07422_));
 sky130_fd_sc_hd__o21a_1 _13570_ (.A1(_07420_),
    .A2(_07421_),
    .B1(_03275_),
    .X(_07423_));
 sky130_fd_sc_hd__o211a_1 _13571_ (.A1(_04602_),
    .A2(_07315_),
    .B1(_07382_),
    .C1(_07254_),
    .X(_07424_));
 sky130_fd_sc_hd__or2_1 _13572_ (.A(_04754_),
    .B(_07276_),
    .X(_07425_));
 sky130_fd_sc_hd__o211a_1 _13573_ (.A1(_04466_),
    .A2(_07315_),
    .B1(_07425_),
    .C1(_07216_),
    .X(_07426_));
 sky130_fd_sc_hd__or3_1 _13574_ (.A(_07190_),
    .B(_07424_),
    .C(_07426_),
    .X(_07427_));
 sky130_fd_sc_hd__nor2_1 _13575_ (.A(_03387_),
    .B(_04631_),
    .Y(_07428_));
 sky130_fd_sc_hd__a211o_1 _13576_ (.A1(\reg_pc[14] ),
    .A2(_07211_),
    .B1(_07428_),
    .C1(_07221_),
    .X(_07429_));
 sky130_fd_sc_hd__a22o_1 _13577_ (.A1(_07422_),
    .A2(_07423_),
    .B1(_07427_),
    .B2(_07429_),
    .X(_07430_));
 sky130_fd_sc_hd__mux2_1 _13578_ (.A0(_04611_),
    .A1(_07430_),
    .S(_07374_),
    .X(_07431_));
 sky130_fd_sc_hd__clkbuf_1 _13579_ (.A(_07431_),
    .X(_00816_));
 sky130_fd_sc_hd__or2_1 _13580_ (.A(net73),
    .B(\decoded_imm[15] ),
    .X(_07432_));
 sky130_fd_sc_hd__nand2_1 _13581_ (.A(net73),
    .B(\decoded_imm[15] ),
    .Y(_07433_));
 sky130_fd_sc_hd__nand2_1 _13582_ (.A(_07418_),
    .B(_07422_),
    .Y(_07434_));
 sky130_fd_sc_hd__a21oi_1 _13583_ (.A1(_07432_),
    .A2(_07433_),
    .B1(_07434_),
    .Y(_07435_));
 sky130_fd_sc_hd__a31o_1 _13584_ (.A1(_07432_),
    .A2(_07433_),
    .A3(_07434_),
    .B1(_03311_),
    .X(_07436_));
 sky130_fd_sc_hd__nor2_1 _13585_ (.A(_07435_),
    .B(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__mux2_1 _13586_ (.A0(_04532_),
    .A1(_04810_),
    .S(_07315_),
    .X(_07438_));
 sky130_fd_sc_hd__o211a_1 _13587_ (.A1(_04611_),
    .A2(_05259_),
    .B1(_07389_),
    .C1(_07254_),
    .X(_07439_));
 sky130_fd_sc_hd__a211o_1 _13588_ (.A1(_07217_),
    .A2(_07438_),
    .B1(_07439_),
    .C1(_07190_),
    .X(_07440_));
 sky130_fd_sc_hd__inv_2 _13589_ (.A(_04659_),
    .Y(_07441_));
 sky130_fd_sc_hd__a22o_1 _13590_ (.A1(_07281_),
    .A2(_07441_),
    .B1(_07305_),
    .B2(\reg_pc[15] ),
    .X(_07442_));
 sky130_fd_sc_hd__o22a_1 _13591_ (.A1(_07437_),
    .A2(_07440_),
    .B1(_07442_),
    .B2(_07284_),
    .X(_07443_));
 sky130_fd_sc_hd__mux2_1 _13592_ (.A0(_04642_),
    .A1(_07443_),
    .S(_07374_),
    .X(_07444_));
 sky130_fd_sc_hd__clkbuf_1 _13593_ (.A(_07444_),
    .X(_00817_));
 sky130_fd_sc_hd__nand2_1 _13594_ (.A(net74),
    .B(\decoded_imm[16] ),
    .Y(_07445_));
 sky130_fd_sc_hd__or2_1 _13595_ (.A(net74),
    .B(\decoded_imm[16] ),
    .X(_07446_));
 sky130_fd_sc_hd__nand2_1 _13596_ (.A(_07445_),
    .B(_07446_),
    .Y(_07447_));
 sky130_fd_sc_hd__a21bo_1 _13597_ (.A1(_07418_),
    .A2(_07422_),
    .B1_N(_07432_),
    .X(_07448_));
 sky130_fd_sc_hd__nand3_1 _13598_ (.A(_07433_),
    .B(_07447_),
    .C(_07448_),
    .Y(_07449_));
 sky130_fd_sc_hd__a21o_1 _13599_ (.A1(_07433_),
    .A2(_07448_),
    .B1(_07447_),
    .X(_07450_));
 sky130_fd_sc_hd__or2_1 _13600_ (.A(_04848_),
    .B(_05227_),
    .X(_07451_));
 sky130_fd_sc_hd__o211a_1 _13601_ (.A1(_04566_),
    .A2(_05259_),
    .B1(_07451_),
    .C1(_07217_),
    .X(_07452_));
 sky130_fd_sc_hd__or2_1 _13602_ (.A(_04642_),
    .B(_05258_),
    .X(_07453_));
 sky130_fd_sc_hd__a31o_1 _13603_ (.A1(_07254_),
    .A2(_07412_),
    .A3(_07453_),
    .B1(_07189_),
    .X(_07454_));
 sky130_fd_sc_hd__a2bb2o_1 _13604_ (.A1_N(_03387_),
    .A2_N(_04702_),
    .B1(_07210_),
    .B2(\reg_pc[16] ),
    .X(_07455_));
 sky130_fd_sc_hd__o22a_1 _13605_ (.A1(_07452_),
    .A2(_07454_),
    .B1(_07455_),
    .B2(_07283_),
    .X(_07456_));
 sky130_fd_sc_hd__a31o_1 _13606_ (.A1(_03276_),
    .A2(_07449_),
    .A3(_07450_),
    .B1(_07456_),
    .X(_07457_));
 sky130_fd_sc_hd__mux2_1 _13607_ (.A0(_04708_),
    .A1(_07457_),
    .S(_07374_),
    .X(_07458_));
 sky130_fd_sc_hd__clkbuf_1 _13608_ (.A(_07458_),
    .X(_00818_));
 sky130_fd_sc_hd__nand2_1 _13609_ (.A(net75),
    .B(\decoded_imm[17] ),
    .Y(_07459_));
 sky130_fd_sc_hd__or2_1 _13610_ (.A(net75),
    .B(\decoded_imm[17] ),
    .X(_07460_));
 sky130_fd_sc_hd__nand2_1 _13611_ (.A(_07459_),
    .B(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__a31o_1 _13612_ (.A1(_07445_),
    .A2(_07450_),
    .A3(_07461_),
    .B1(_03311_),
    .X(_07462_));
 sky130_fd_sc_hd__a21o_1 _13613_ (.A1(_07445_),
    .A2(_07450_),
    .B1(_07461_),
    .X(_07463_));
 sky130_fd_sc_hd__and2b_1 _13614_ (.A_N(_07462_),
    .B(_07463_),
    .X(_07464_));
 sky130_fd_sc_hd__nand2_1 _13615_ (.A(_03575_),
    .B(_07236_),
    .Y(_07465_));
 sky130_fd_sc_hd__o211a_1 _13616_ (.A1(_04602_),
    .A2(_07236_),
    .B1(_07465_),
    .C1(_07217_),
    .X(_07466_));
 sky130_fd_sc_hd__o211a_1 _13617_ (.A1(_04708_),
    .A2(_05260_),
    .B1(_07425_),
    .C1(_07238_),
    .X(_07467_));
 sky130_fd_sc_hd__a221o_1 _13618_ (.A1(_07304_),
    .A2(_04738_),
    .B1(_07305_),
    .B2(\reg_pc[17] ),
    .C1(_07283_),
    .X(_07468_));
 sky130_fd_sc_hd__o41a_1 _13619_ (.A1(_07191_),
    .A2(_07464_),
    .A3(_07466_),
    .A4(_07467_),
    .B1(_07468_),
    .X(_07469_));
 sky130_fd_sc_hd__mux2_1 _13620_ (.A0(_04744_),
    .A1(_07469_),
    .S(_07374_),
    .X(_07470_));
 sky130_fd_sc_hd__clkbuf_1 _13621_ (.A(_07470_),
    .X(_00819_));
 sky130_fd_sc_hd__a22o_1 _13622_ (.A1(_07281_),
    .A2(_04777_),
    .B1(_07282_),
    .B2(\reg_pc[18] ),
    .X(_07471_));
 sky130_fd_sc_hd__nand2_1 _13623_ (.A(net76),
    .B(\decoded_imm[18] ),
    .Y(_07472_));
 sky130_fd_sc_hd__or2_1 _13624_ (.A(net76),
    .B(\decoded_imm[18] ),
    .X(_07473_));
 sky130_fd_sc_hd__nand2_1 _13625_ (.A(_07472_),
    .B(_07473_),
    .Y(_07474_));
 sky130_fd_sc_hd__nand2_1 _13626_ (.A(_07459_),
    .B(_07463_),
    .Y(_07475_));
 sky130_fd_sc_hd__xnor2_1 _13627_ (.A(_07474_),
    .B(_07475_),
    .Y(_07476_));
 sky130_fd_sc_hd__mux2_1 _13628_ (.A0(_04810_),
    .A1(_04744_),
    .S(_07276_),
    .X(_07477_));
 sky130_fd_sc_hd__mux2_1 _13629_ (.A0(_04611_),
    .A1(_04913_),
    .S(_05258_),
    .X(_07478_));
 sky130_fd_sc_hd__a22o_1 _13630_ (.A1(_07254_),
    .A2(_07477_),
    .B1(_07478_),
    .B2(_07217_),
    .X(_07479_));
 sky130_fd_sc_hd__a211o_1 _13631_ (.A1(_03275_),
    .A2(_07476_),
    .B1(_07479_),
    .C1(_07232_),
    .X(_07480_));
 sky130_fd_sc_hd__o21a_1 _13632_ (.A1(_07284_),
    .A2(_07471_),
    .B1(_07480_),
    .X(_07481_));
 sky130_fd_sc_hd__mux2_1 _13633_ (.A0(_04754_),
    .A1(_07481_),
    .S(_07374_),
    .X(_07482_));
 sky130_fd_sc_hd__clkbuf_1 _13634_ (.A(_07482_),
    .X(_00820_));
 sky130_fd_sc_hd__o211a_1 _13635_ (.A1(_04754_),
    .A2(_05261_),
    .B1(_07451_),
    .C1(_07279_),
    .X(_07483_));
 sky130_fd_sc_hd__mux2_1 _13636_ (.A0(_04642_),
    .A1(_04945_),
    .S(_07236_),
    .X(_07484_));
 sky130_fd_sc_hd__a21o_1 _13637_ (.A1(_07274_),
    .A2(_07484_),
    .B1(_07191_),
    .X(_07485_));
 sky130_fd_sc_hd__a22o_1 _13638_ (.A1(_07281_),
    .A2(_04806_),
    .B1(_07282_),
    .B2(\reg_pc[19] ),
    .X(_07486_));
 sky130_fd_sc_hd__o22a_1 _13639_ (.A1(_07483_),
    .A2(_07485_),
    .B1(_07486_),
    .B2(_07284_),
    .X(_07487_));
 sky130_fd_sc_hd__nand2_1 _13640_ (.A(net77),
    .B(\decoded_imm[19] ),
    .Y(_07488_));
 sky130_fd_sc_hd__or2_1 _13641_ (.A(net77),
    .B(\decoded_imm[19] ),
    .X(_07489_));
 sky130_fd_sc_hd__nand2_1 _13642_ (.A(_07488_),
    .B(_07489_),
    .Y(_07490_));
 sky130_fd_sc_hd__a21boi_1 _13643_ (.A1(_07473_),
    .A2(_07475_),
    .B1_N(_07472_),
    .Y(_07491_));
 sky130_fd_sc_hd__xnor2_1 _13644_ (.A(_07490_),
    .B(_07491_),
    .Y(_07492_));
 sky130_fd_sc_hd__o21ai_1 _13645_ (.A1(_03631_),
    .A2(_07492_),
    .B1(_07271_),
    .Y(_07493_));
 sky130_fd_sc_hd__o22a_1 _13646_ (.A1(_04810_),
    .A2(_07271_),
    .B1(_07487_),
    .B2(_07493_),
    .X(_00821_));
 sky130_fd_sc_hd__o211a_1 _13647_ (.A1(_04810_),
    .A2(_05260_),
    .B1(_07465_),
    .C1(_07279_),
    .X(_07494_));
 sky130_fd_sc_hd__or2_1 _13648_ (.A(_04959_),
    .B(_07277_),
    .X(_07495_));
 sky130_fd_sc_hd__o211a_1 _13649_ (.A1(_04708_),
    .A2(_05261_),
    .B1(_07495_),
    .C1(_07274_),
    .X(_07496_));
 sky130_fd_sc_hd__a221o_1 _13650_ (.A1(_07281_),
    .A2(_04842_),
    .B1(_07282_),
    .B2(\reg_pc[20] ),
    .C1(_07283_),
    .X(_07497_));
 sky130_fd_sc_hd__o31a_1 _13651_ (.A1(_07191_),
    .A2(_07494_),
    .A3(_07496_),
    .B1(_07497_),
    .X(_07498_));
 sky130_fd_sc_hd__nand2_1 _13652_ (.A(net79),
    .B(\decoded_imm[20] ),
    .Y(_07499_));
 sky130_fd_sc_hd__or2_1 _13653_ (.A(net79),
    .B(\decoded_imm[20] ),
    .X(_07500_));
 sky130_fd_sc_hd__nand2_1 _13654_ (.A(_07499_),
    .B(_07500_),
    .Y(_07501_));
 sky130_fd_sc_hd__or4_1 _13655_ (.A(_07450_),
    .B(_07461_),
    .C(_07474_),
    .D(_07490_),
    .X(_07502_));
 sky130_fd_sc_hd__or2b_1 _13656_ (.A(_07445_),
    .B_N(_07460_),
    .X(_07503_));
 sky130_fd_sc_hd__a211o_1 _13657_ (.A1(_07459_),
    .A2(_07503_),
    .B1(_07490_),
    .C1(_07474_),
    .X(_07504_));
 sky130_fd_sc_hd__or2b_1 _13658_ (.A(_07472_),
    .B_N(_07489_),
    .X(_07505_));
 sky130_fd_sc_hd__and4_1 _13659_ (.A(_07488_),
    .B(_07502_),
    .C(_07504_),
    .D(_07505_),
    .X(_07506_));
 sky130_fd_sc_hd__nand2_1 _13660_ (.A(_07501_),
    .B(_07506_),
    .Y(_07507_));
 sky130_fd_sc_hd__a41o_1 _13661_ (.A1(_07488_),
    .A2(_07502_),
    .A3(_07504_),
    .A4(_07505_),
    .B1(_07501_),
    .X(_07508_));
 sky130_fd_sc_hd__and2_1 _13662_ (.A(_03276_),
    .B(_07508_),
    .X(_07509_));
 sky130_fd_sc_hd__a21bo_1 _13663_ (.A1(_07507_),
    .A2(_07509_),
    .B1_N(_07225_),
    .X(_07510_));
 sky130_fd_sc_hd__o22a_1 _13664_ (.A1(_04848_),
    .A2(_07271_),
    .B1(_07498_),
    .B2(_07510_),
    .X(_00822_));
 sky130_fd_sc_hd__nand2_1 _13665_ (.A(_04880_),
    .B(\decoded_imm[21] ),
    .Y(_07511_));
 sky130_fd_sc_hd__or2_1 _13666_ (.A(net80),
    .B(\decoded_imm[21] ),
    .X(_07512_));
 sky130_fd_sc_hd__nand2_1 _13667_ (.A(_07511_),
    .B(_07512_),
    .Y(_07513_));
 sky130_fd_sc_hd__a31o_1 _13668_ (.A1(_07499_),
    .A2(_07508_),
    .A3(_07513_),
    .B1(_03311_),
    .X(_07514_));
 sky130_fd_sc_hd__a21o_1 _13669_ (.A1(_07499_),
    .A2(_07508_),
    .B1(_07513_),
    .X(_07515_));
 sky130_fd_sc_hd__and2b_1 _13670_ (.A_N(_07514_),
    .B(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__nand2_1 _13671_ (.A(_03584_),
    .B(_05257_),
    .Y(_07517_));
 sky130_fd_sc_hd__o211a_1 _13672_ (.A1(_04744_),
    .A2(_07236_),
    .B1(_07517_),
    .C1(_07217_),
    .X(_07518_));
 sky130_fd_sc_hd__or2_1 _13673_ (.A(_04848_),
    .B(_05258_),
    .X(_07519_));
 sky130_fd_sc_hd__o211a_1 _13674_ (.A1(_04913_),
    .A2(_07277_),
    .B1(_07519_),
    .C1(_07238_),
    .X(_07520_));
 sky130_fd_sc_hd__a221o_1 _13675_ (.A1(_07304_),
    .A2(_04871_),
    .B1(_07305_),
    .B2(\reg_pc[21] ),
    .C1(_07283_),
    .X(_07521_));
 sky130_fd_sc_hd__o41a_1 _13676_ (.A1(_07191_),
    .A2(_07516_),
    .A3(_07518_),
    .A4(_07520_),
    .B1(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__mux2_1 _13677_ (.A0(_04880_),
    .A1(_07522_),
    .S(_07374_),
    .X(_07523_));
 sky130_fd_sc_hd__clkbuf_1 _13678_ (.A(_07523_),
    .X(_00823_));
 sky130_fd_sc_hd__nand2_1 _13679_ (.A(net81),
    .B(\decoded_imm[22] ),
    .Y(_07524_));
 sky130_fd_sc_hd__or2_1 _13680_ (.A(net81),
    .B(\decoded_imm[22] ),
    .X(_07525_));
 sky130_fd_sc_hd__nand2_1 _13681_ (.A(_07524_),
    .B(_07525_),
    .Y(_07526_));
 sky130_fd_sc_hd__a21oi_1 _13682_ (.A1(_07511_),
    .A2(_07515_),
    .B1(_07526_),
    .Y(_07527_));
 sky130_fd_sc_hd__a31o_1 _13683_ (.A1(_07511_),
    .A2(_07515_),
    .A3(_07526_),
    .B1(_03311_),
    .X(_07528_));
 sky130_fd_sc_hd__nor2_1 _13684_ (.A(_07527_),
    .B(_07528_),
    .Y(_07529_));
 sky130_fd_sc_hd__or2_1 _13685_ (.A(_05044_),
    .B(_07277_),
    .X(_07530_));
 sky130_fd_sc_hd__o211a_1 _13686_ (.A1(_04754_),
    .A2(_07236_),
    .B1(_07530_),
    .C1(_07217_),
    .X(_07531_));
 sky130_fd_sc_hd__nand2_1 _13687_ (.A(_03575_),
    .B(_07277_),
    .Y(_07532_));
 sky130_fd_sc_hd__o211a_1 _13688_ (.A1(_04945_),
    .A2(_07277_),
    .B1(_07532_),
    .C1(_07238_),
    .X(_07533_));
 sky130_fd_sc_hd__a221o_1 _13689_ (.A1(_07304_),
    .A2(_04909_),
    .B1(_07305_),
    .B2(\reg_pc[22] ),
    .C1(_07283_),
    .X(_07534_));
 sky130_fd_sc_hd__o41a_1 _13690_ (.A1(_07232_),
    .A2(_07529_),
    .A3(_07531_),
    .A4(_07533_),
    .B1(_07534_),
    .X(_07535_));
 sky130_fd_sc_hd__mux2_1 _13691_ (.A0(_04913_),
    .A1(_07535_),
    .S(_07224_),
    .X(_07536_));
 sky130_fd_sc_hd__clkbuf_1 _13692_ (.A(_07536_),
    .X(_00824_));
 sky130_fd_sc_hd__o211a_1 _13693_ (.A1(_04913_),
    .A2(_05261_),
    .B1(_07495_),
    .C1(_07279_),
    .X(_07537_));
 sky130_fd_sc_hd__mux2_1 _13694_ (.A0(_05076_),
    .A1(_04810_),
    .S(_07277_),
    .X(_07538_));
 sky130_fd_sc_hd__a21o_1 _13695_ (.A1(_07274_),
    .A2(_07538_),
    .B1(_07191_),
    .X(_07539_));
 sky130_fd_sc_hd__a22o_1 _13696_ (.A1(_07281_),
    .A2(_04941_),
    .B1(_07282_),
    .B2(\reg_pc[23] ),
    .X(_07540_));
 sky130_fd_sc_hd__o22a_1 _13697_ (.A1(_07537_),
    .A2(_07539_),
    .B1(_07540_),
    .B2(_07284_),
    .X(_07541_));
 sky130_fd_sc_hd__nand2_1 _13698_ (.A(net82),
    .B(\decoded_imm[23] ),
    .Y(_07542_));
 sky130_fd_sc_hd__or2_1 _13699_ (.A(net82),
    .B(\decoded_imm[23] ),
    .X(_07543_));
 sky130_fd_sc_hd__nand2_1 _13700_ (.A(_07542_),
    .B(_07543_),
    .Y(_07544_));
 sky130_fd_sc_hd__a21oi_1 _13701_ (.A1(_04913_),
    .A2(\decoded_imm[22] ),
    .B1(_07527_),
    .Y(_07545_));
 sky130_fd_sc_hd__xnor2_1 _13702_ (.A(_07544_),
    .B(_07545_),
    .Y(_07546_));
 sky130_fd_sc_hd__o21ai_1 _13703_ (.A1(_03631_),
    .A2(_07546_),
    .B1(_07271_),
    .Y(_07547_));
 sky130_fd_sc_hd__o22a_1 _13704_ (.A1(_04945_),
    .A2(_07271_),
    .B1(_07541_),
    .B2(_07547_),
    .X(_00825_));
 sky130_fd_sc_hd__or3_1 _13705_ (.A(_07513_),
    .B(_07526_),
    .C(_07544_),
    .X(_07548_));
 sky130_fd_sc_hd__nor2_1 _13706_ (.A(net82),
    .B(\decoded_imm[23] ),
    .Y(_07549_));
 sky130_fd_sc_hd__nor2_1 _13707_ (.A(_04880_),
    .B(\decoded_imm[21] ),
    .Y(_07550_));
 sky130_fd_sc_hd__o21a_1 _13708_ (.A1(_07499_),
    .A2(_07550_),
    .B1(_07511_),
    .X(_07551_));
 sky130_fd_sc_hd__or2_1 _13709_ (.A(_07524_),
    .B(_07549_),
    .X(_07552_));
 sky130_fd_sc_hd__o311a_1 _13710_ (.A1(_07526_),
    .A2(_07549_),
    .A3(_07551_),
    .B1(_07552_),
    .C1(_07542_),
    .X(_07553_));
 sky130_fd_sc_hd__o21ai_1 _13711_ (.A1(_07508_),
    .A2(_07548_),
    .B1(_07553_),
    .Y(_07554_));
 sky130_fd_sc_hd__nand2_1 _13712_ (.A(net83),
    .B(\decoded_imm[24] ),
    .Y(_07555_));
 sky130_fd_sc_hd__or2_1 _13713_ (.A(net83),
    .B(\decoded_imm[24] ),
    .X(_07556_));
 sky130_fd_sc_hd__and2_1 _13714_ (.A(_07555_),
    .B(_07556_),
    .X(_07557_));
 sky130_fd_sc_hd__nand2_1 _13715_ (.A(_07554_),
    .B(_07557_),
    .Y(_07558_));
 sky130_fd_sc_hd__or2_1 _13716_ (.A(_07554_),
    .B(_07557_),
    .X(_07559_));
 sky130_fd_sc_hd__or2_1 _13717_ (.A(_05086_),
    .B(_05227_),
    .X(_07560_));
 sky130_fd_sc_hd__o211a_1 _13718_ (.A1(_04945_),
    .A2(_05258_),
    .B1(_07517_),
    .C1(_07237_),
    .X(_07561_));
 sky130_fd_sc_hd__a31o_1 _13719_ (.A1(_07217_),
    .A2(_07519_),
    .A3(_07560_),
    .B1(_07561_),
    .X(_07562_));
 sky130_fd_sc_hd__a221o_1 _13720_ (.A1(_07209_),
    .A2(_04979_),
    .B1(_07211_),
    .B2(\reg_pc[24] ),
    .C1(_07221_),
    .X(_07563_));
 sky130_fd_sc_hd__o21a_1 _13721_ (.A1(_07232_),
    .A2(_07562_),
    .B1(_07563_),
    .X(_07564_));
 sky130_fd_sc_hd__a31o_1 _13722_ (.A1(_03276_),
    .A2(_07558_),
    .A3(_07559_),
    .B1(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__mux2_1 _13723_ (.A0(_04959_),
    .A1(_07565_),
    .S(_07224_),
    .X(_07566_));
 sky130_fd_sc_hd__clkbuf_1 _13724_ (.A(_07566_),
    .X(_00826_));
 sky130_fd_sc_hd__or2_1 _13725_ (.A(net84),
    .B(\decoded_imm[25] ),
    .X(_07567_));
 sky130_fd_sc_hd__nand2_1 _13726_ (.A(_05013_),
    .B(\decoded_imm[25] ),
    .Y(_07568_));
 sky130_fd_sc_hd__nand2_1 _13727_ (.A(_07567_),
    .B(_07568_),
    .Y(_07569_));
 sky130_fd_sc_hd__nand3_1 _13728_ (.A(_07555_),
    .B(_07558_),
    .C(_07569_),
    .Y(_07570_));
 sky130_fd_sc_hd__a21o_1 _13729_ (.A1(_07555_),
    .A2(_07558_),
    .B1(_07569_),
    .X(_07571_));
 sky130_fd_sc_hd__and3_1 _13730_ (.A(_03275_),
    .B(_07570_),
    .C(_07571_),
    .X(_07572_));
 sky130_fd_sc_hd__o211a_1 _13731_ (.A1(_05143_),
    .A2(_07277_),
    .B1(_07532_),
    .C1(_07217_),
    .X(_07573_));
 sky130_fd_sc_hd__o211a_1 _13732_ (.A1(_04959_),
    .A2(_07236_),
    .B1(_07530_),
    .C1(_07238_),
    .X(_07574_));
 sky130_fd_sc_hd__a221o_1 _13733_ (.A1(_07304_),
    .A2(_05009_),
    .B1(_07305_),
    .B2(\reg_pc[25] ),
    .C1(_07283_),
    .X(_07575_));
 sky130_fd_sc_hd__o41a_1 _13734_ (.A1(_07232_),
    .A2(_07572_),
    .A3(_07573_),
    .A4(_07574_),
    .B1(_07575_),
    .X(_07576_));
 sky130_fd_sc_hd__mux2_1 _13735_ (.A0(_05013_),
    .A1(_07576_),
    .S(_07224_),
    .X(_07577_));
 sky130_fd_sc_hd__clkbuf_1 _13736_ (.A(_07577_),
    .X(_00827_));
 sky130_fd_sc_hd__nand2_1 _13737_ (.A(net85),
    .B(\decoded_imm[26] ),
    .Y(_07578_));
 sky130_fd_sc_hd__or2_1 _13738_ (.A(net85),
    .B(\decoded_imm[26] ),
    .X(_07579_));
 sky130_fd_sc_hd__nand2_1 _13739_ (.A(_07578_),
    .B(_07579_),
    .Y(_07580_));
 sky130_fd_sc_hd__a21o_1 _13740_ (.A1(_07568_),
    .A2(_07571_),
    .B1(_07580_),
    .X(_07581_));
 sky130_fd_sc_hd__nand3_1 _13741_ (.A(_07568_),
    .B(_07571_),
    .C(_07580_),
    .Y(_07582_));
 sky130_fd_sc_hd__nor2_1 _13742_ (.A(_05013_),
    .B(_05258_),
    .Y(_07583_));
 sky130_fd_sc_hd__a21oi_1 _13743_ (.A1(_03583_),
    .A2(_07315_),
    .B1(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__mux2_1 _13744_ (.A0(_05174_),
    .A1(_04913_),
    .S(_07276_),
    .X(_07585_));
 sky130_fd_sc_hd__a22o_1 _13745_ (.A1(_07254_),
    .A2(_07584_),
    .B1(_07585_),
    .B2(_07216_),
    .X(_07586_));
 sky130_fd_sc_hd__inv_2 _13746_ (.A(_05037_),
    .Y(_07587_));
 sky130_fd_sc_hd__a22o_1 _13747_ (.A1(_07209_),
    .A2(_07587_),
    .B1(_07210_),
    .B2(\reg_pc[26] ),
    .X(_07588_));
 sky130_fd_sc_hd__mux2_1 _13748_ (.A0(_07586_),
    .A1(_07588_),
    .S(_07190_),
    .X(_07589_));
 sky130_fd_sc_hd__a31o_1 _13749_ (.A1(_03276_),
    .A2(_07581_),
    .A3(_07582_),
    .B1(_07589_),
    .X(_07590_));
 sky130_fd_sc_hd__mux2_1 _13750_ (.A0(_05044_),
    .A1(_07590_),
    .S(_07224_),
    .X(_07591_));
 sky130_fd_sc_hd__clkbuf_1 _13751_ (.A(_07591_),
    .X(_00828_));
 sky130_fd_sc_hd__o211a_1 _13752_ (.A1(_05044_),
    .A2(_05260_),
    .B1(_07560_),
    .C1(_07279_),
    .X(_07592_));
 sky130_fd_sc_hd__or2_1 _13753_ (.A(_05205_),
    .B(_05227_),
    .X(_07593_));
 sky130_fd_sc_hd__o211a_1 _13754_ (.A1(_04945_),
    .A2(_05261_),
    .B1(_07593_),
    .C1(_07274_),
    .X(_07594_));
 sky130_fd_sc_hd__inv_2 _13755_ (.A(_05069_),
    .Y(_07595_));
 sky130_fd_sc_hd__a221o_1 _13756_ (.A1(_07281_),
    .A2(_07595_),
    .B1(_07282_),
    .B2(\reg_pc[27] ),
    .C1(_07283_),
    .X(_07596_));
 sky130_fd_sc_hd__o31a_1 _13757_ (.A1(_07191_),
    .A2(_07592_),
    .A3(_07594_),
    .B1(_07596_),
    .X(_07597_));
 sky130_fd_sc_hd__xnor2_1 _13758_ (.A(net86),
    .B(\decoded_imm[27] ),
    .Y(_07598_));
 sky130_fd_sc_hd__and3_1 _13759_ (.A(_07578_),
    .B(_07581_),
    .C(_07598_),
    .X(_07599_));
 sky130_fd_sc_hd__a21oi_1 _13760_ (.A1(_07578_),
    .A2(_07581_),
    .B1(_07598_),
    .Y(_07600_));
 sky130_fd_sc_hd__o31ai_1 _13761_ (.A1(_03631_),
    .A2(_07599_),
    .A3(_07600_),
    .B1(_07225_),
    .Y(_07601_));
 sky130_fd_sc_hd__o22a_1 _13762_ (.A1(_05076_),
    .A2(_07271_),
    .B1(_07597_),
    .B2(_07601_),
    .X(_00829_));
 sky130_fd_sc_hd__nor2_1 _13763_ (.A(_07580_),
    .B(_07598_),
    .Y(_07602_));
 sky130_fd_sc_hd__inv_2 _13764_ (.A(_07602_),
    .Y(_07603_));
 sky130_fd_sc_hd__or2b_1 _13765_ (.A(_07555_),
    .B_N(_07567_),
    .X(_07604_));
 sky130_fd_sc_hd__a21o_1 _13766_ (.A1(_07568_),
    .A2(_07604_),
    .B1(_07603_),
    .X(_07605_));
 sky130_fd_sc_hd__o211a_1 _13767_ (.A1(net86),
    .A2(\decoded_imm[27] ),
    .B1(\decoded_imm[26] ),
    .C1(net85),
    .X(_07606_));
 sky130_fd_sc_hd__a21oi_1 _13768_ (.A1(net86),
    .A2(\decoded_imm[27] ),
    .B1(_07606_),
    .Y(_07607_));
 sky130_fd_sc_hd__o311a_1 _13769_ (.A1(_07558_),
    .A2(_07569_),
    .A3(_07603_),
    .B1(_07605_),
    .C1(_07607_),
    .X(_07608_));
 sky130_fd_sc_hd__and2_1 _13770_ (.A(net87),
    .B(\decoded_imm[28] ),
    .X(_07609_));
 sky130_fd_sc_hd__nor2_1 _13771_ (.A(net87),
    .B(\decoded_imm[28] ),
    .Y(_07610_));
 sky130_fd_sc_hd__or3_1 _13772_ (.A(_07608_),
    .B(_07609_),
    .C(_07610_),
    .X(_07611_));
 sky130_fd_sc_hd__o21ai_1 _13773_ (.A1(_07609_),
    .A2(_07610_),
    .B1(_07608_),
    .Y(_07612_));
 sky130_fd_sc_hd__mux2_1 _13774_ (.A0(_05143_),
    .A1(_05076_),
    .S(_05227_),
    .X(_07613_));
 sky130_fd_sc_hd__o21ai_1 _13775_ (.A1(_05227_),
    .A2(_05334_),
    .B1(_07216_),
    .Y(_07614_));
 sky130_fd_sc_hd__o21ba_1 _13776_ (.A1(_04959_),
    .A2(_07236_),
    .B1_N(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__a211o_1 _13777_ (.A1(_07238_),
    .A2(_07613_),
    .B1(_07615_),
    .C1(_07232_),
    .X(_07616_));
 sky130_fd_sc_hd__a221o_1 _13778_ (.A1(_07304_),
    .A2(_05107_),
    .B1(_07211_),
    .B2(\reg_pc[28] ),
    .C1(_07221_),
    .X(_07617_));
 sky130_fd_sc_hd__a32o_1 _13779_ (.A1(_03275_),
    .A2(_07611_),
    .A3(_07612_),
    .B1(_07616_),
    .B2(_07617_),
    .X(_07618_));
 sky130_fd_sc_hd__mux2_1 _13780_ (.A0(_05086_),
    .A1(_07618_),
    .S(_07224_),
    .X(_07619_));
 sky130_fd_sc_hd__clkbuf_1 _13781_ (.A(_07619_),
    .X(_00830_));
 sky130_fd_sc_hd__nand2_1 _13782_ (.A(net88),
    .B(\decoded_imm[29] ),
    .Y(_07620_));
 sky130_fd_sc_hd__or2_1 _13783_ (.A(net88),
    .B(\decoded_imm[29] ),
    .X(_07621_));
 sky130_fd_sc_hd__nand2_1 _13784_ (.A(_07620_),
    .B(_07621_),
    .Y(_07622_));
 sky130_fd_sc_hd__nand2_1 _13785_ (.A(_07611_),
    .B(_07622_),
    .Y(_07623_));
 sky130_fd_sc_hd__nand2_1 _13786_ (.A(_05086_),
    .B(\decoded_imm[28] ),
    .Y(_07624_));
 sky130_fd_sc_hd__a21o_1 _13787_ (.A1(_07624_),
    .A2(_07611_),
    .B1(_07622_),
    .X(_07625_));
 sky130_fd_sc_hd__o211a_1 _13788_ (.A1(_07609_),
    .A2(_07623_),
    .B1(_07625_),
    .C1(_03275_),
    .X(_07626_));
 sky130_fd_sc_hd__mux2_1 _13789_ (.A0(_05174_),
    .A1(_05086_),
    .S(_05227_),
    .X(_07627_));
 sky130_fd_sc_hd__nor2_1 _13790_ (.A(_07583_),
    .B(_07614_),
    .Y(_07628_));
 sky130_fd_sc_hd__a211o_1 _13791_ (.A1(_07238_),
    .A2(_07627_),
    .B1(_07628_),
    .C1(_07190_),
    .X(_07629_));
 sky130_fd_sc_hd__a22o_1 _13792_ (.A1(_07304_),
    .A2(_05139_),
    .B1(_07305_),
    .B2(\reg_pc[29] ),
    .X(_07630_));
 sky130_fd_sc_hd__o22a_1 _13793_ (.A1(_07626_),
    .A2(_07629_),
    .B1(_07630_),
    .B2(_07284_),
    .X(_07631_));
 sky130_fd_sc_hd__mux2_1 _13794_ (.A0(_05143_),
    .A1(_07631_),
    .S(_07224_),
    .X(_07632_));
 sky130_fd_sc_hd__clkbuf_1 _13795_ (.A(_07632_),
    .X(_00831_));
 sky130_fd_sc_hd__and2_1 _13796_ (.A(_05174_),
    .B(\decoded_imm[30] ),
    .X(_07633_));
 sky130_fd_sc_hd__nor2_1 _13797_ (.A(_05174_),
    .B(\decoded_imm[30] ),
    .Y(_07634_));
 sky130_fd_sc_hd__o211a_1 _13798_ (.A1(_07633_),
    .A2(_07634_),
    .B1(_07620_),
    .C1(_07625_),
    .X(_07635_));
 sky130_fd_sc_hd__a211oi_2 _13799_ (.A1(_07620_),
    .A2(_07625_),
    .B1(_07633_),
    .C1(_07634_),
    .Y(_07636_));
 sky130_fd_sc_hd__nor3_1 _13800_ (.A(_03631_),
    .B(_07635_),
    .C(_07636_),
    .Y(_07637_));
 sky130_fd_sc_hd__o211a_1 _13801_ (.A1(_05143_),
    .A2(_07236_),
    .B1(_07593_),
    .C1(_07238_),
    .X(_07638_));
 sky130_fd_sc_hd__o21ba_1 _13802_ (.A1(_05044_),
    .A2(_05260_),
    .B1_N(_07614_),
    .X(_07639_));
 sky130_fd_sc_hd__a221o_1 _13803_ (.A1(_07304_),
    .A2(_05170_),
    .B1(_07305_),
    .B2(\reg_pc[30] ),
    .C1(_07221_),
    .X(_07640_));
 sky130_fd_sc_hd__o41a_1 _13804_ (.A1(_07232_),
    .A2(_07637_),
    .A3(_07638_),
    .A4(_07639_),
    .B1(_07640_),
    .X(_07641_));
 sky130_fd_sc_hd__mux2_1 _13805_ (.A0(_05174_),
    .A1(_07641_),
    .S(_07224_),
    .X(_07642_));
 sky130_fd_sc_hd__clkbuf_1 _13806_ (.A(_07642_),
    .X(_00832_));
 sky130_fd_sc_hd__clkbuf_1 _13807_ (.A(\cpuregs.regs[0][0] ),
    .X(_07643_));
 sky130_fd_sc_hd__clkbuf_1 _13808_ (.A(_07643_),
    .X(_00833_));
 sky130_fd_sc_hd__clkbuf_1 _13809_ (.A(\cpuregs.regs[0][1] ),
    .X(_07644_));
 sky130_fd_sc_hd__clkbuf_1 _13810_ (.A(_07644_),
    .X(_00834_));
 sky130_fd_sc_hd__clkbuf_1 _13811_ (.A(\cpuregs.regs[0][2] ),
    .X(_07645_));
 sky130_fd_sc_hd__clkbuf_1 _13812_ (.A(_07645_),
    .X(_00835_));
 sky130_fd_sc_hd__clkbuf_1 _13813_ (.A(\cpuregs.regs[0][3] ),
    .X(_07646_));
 sky130_fd_sc_hd__clkbuf_1 _13814_ (.A(_07646_),
    .X(_00836_));
 sky130_fd_sc_hd__clkbuf_1 _13815_ (.A(\cpuregs.regs[0][4] ),
    .X(_07647_));
 sky130_fd_sc_hd__clkbuf_1 _13816_ (.A(_07647_),
    .X(_00837_));
 sky130_fd_sc_hd__clkbuf_1 _13817_ (.A(\cpuregs.regs[0][5] ),
    .X(_07648_));
 sky130_fd_sc_hd__clkbuf_1 _13818_ (.A(_07648_),
    .X(_00838_));
 sky130_fd_sc_hd__clkbuf_1 _13819_ (.A(\cpuregs.regs[0][6] ),
    .X(_07649_));
 sky130_fd_sc_hd__clkbuf_1 _13820_ (.A(_07649_),
    .X(_00839_));
 sky130_fd_sc_hd__clkbuf_1 _13821_ (.A(\cpuregs.regs[0][7] ),
    .X(_07650_));
 sky130_fd_sc_hd__clkbuf_1 _13822_ (.A(_07650_),
    .X(_00840_));
 sky130_fd_sc_hd__clkbuf_1 _13823_ (.A(\cpuregs.regs[0][8] ),
    .X(_07651_));
 sky130_fd_sc_hd__clkbuf_1 _13824_ (.A(_07651_),
    .X(_00841_));
 sky130_fd_sc_hd__clkbuf_1 _13825_ (.A(\cpuregs.regs[0][9] ),
    .X(_07652_));
 sky130_fd_sc_hd__clkbuf_1 _13826_ (.A(_07652_),
    .X(_00842_));
 sky130_fd_sc_hd__clkbuf_1 _13827_ (.A(\cpuregs.regs[0][10] ),
    .X(_07653_));
 sky130_fd_sc_hd__clkbuf_1 _13828_ (.A(_07653_),
    .X(_00843_));
 sky130_fd_sc_hd__clkbuf_1 _13829_ (.A(\cpuregs.regs[0][11] ),
    .X(_07654_));
 sky130_fd_sc_hd__clkbuf_1 _13830_ (.A(_07654_),
    .X(_00844_));
 sky130_fd_sc_hd__clkbuf_1 _13831_ (.A(\cpuregs.regs[0][12] ),
    .X(_07655_));
 sky130_fd_sc_hd__clkbuf_1 _13832_ (.A(_07655_),
    .X(_00845_));
 sky130_fd_sc_hd__clkbuf_1 _13833_ (.A(\cpuregs.regs[0][13] ),
    .X(_07656_));
 sky130_fd_sc_hd__clkbuf_1 _13834_ (.A(_07656_),
    .X(_00846_));
 sky130_fd_sc_hd__clkbuf_1 _13835_ (.A(\cpuregs.regs[0][14] ),
    .X(_07657_));
 sky130_fd_sc_hd__clkbuf_1 _13836_ (.A(_07657_),
    .X(_00847_));
 sky130_fd_sc_hd__clkbuf_1 _13837_ (.A(\cpuregs.regs[0][15] ),
    .X(_07658_));
 sky130_fd_sc_hd__clkbuf_1 _13838_ (.A(_07658_),
    .X(_00848_));
 sky130_fd_sc_hd__clkbuf_1 _13839_ (.A(\cpuregs.regs[0][16] ),
    .X(_07659_));
 sky130_fd_sc_hd__clkbuf_1 _13840_ (.A(_07659_),
    .X(_00849_));
 sky130_fd_sc_hd__clkbuf_1 _13841_ (.A(\cpuregs.regs[0][17] ),
    .X(_07660_));
 sky130_fd_sc_hd__clkbuf_1 _13842_ (.A(_07660_),
    .X(_00850_));
 sky130_fd_sc_hd__clkbuf_1 _13843_ (.A(\cpuregs.regs[0][18] ),
    .X(_07661_));
 sky130_fd_sc_hd__clkbuf_1 _13844_ (.A(_07661_),
    .X(_00851_));
 sky130_fd_sc_hd__clkbuf_1 _13845_ (.A(\cpuregs.regs[0][19] ),
    .X(_07662_));
 sky130_fd_sc_hd__clkbuf_1 _13846_ (.A(_07662_),
    .X(_00852_));
 sky130_fd_sc_hd__clkbuf_1 _13847_ (.A(\cpuregs.regs[0][20] ),
    .X(_07663_));
 sky130_fd_sc_hd__clkbuf_1 _13848_ (.A(_07663_),
    .X(_00853_));
 sky130_fd_sc_hd__clkbuf_1 _13849_ (.A(\cpuregs.regs[0][21] ),
    .X(_07664_));
 sky130_fd_sc_hd__clkbuf_1 _13850_ (.A(_07664_),
    .X(_00854_));
 sky130_fd_sc_hd__clkbuf_1 _13851_ (.A(\cpuregs.regs[0][22] ),
    .X(_07665_));
 sky130_fd_sc_hd__clkbuf_1 _13852_ (.A(_07665_),
    .X(_00855_));
 sky130_fd_sc_hd__clkbuf_1 _13853_ (.A(\cpuregs.regs[0][23] ),
    .X(_07666_));
 sky130_fd_sc_hd__clkbuf_1 _13854_ (.A(_07666_),
    .X(_00856_));
 sky130_fd_sc_hd__clkbuf_1 _13855_ (.A(\cpuregs.regs[0][24] ),
    .X(_07667_));
 sky130_fd_sc_hd__clkbuf_1 _13856_ (.A(_07667_),
    .X(_00857_));
 sky130_fd_sc_hd__clkbuf_1 _13857_ (.A(\cpuregs.regs[0][25] ),
    .X(_07668_));
 sky130_fd_sc_hd__clkbuf_1 _13858_ (.A(_07668_),
    .X(_00858_));
 sky130_fd_sc_hd__clkbuf_1 _13859_ (.A(\cpuregs.regs[0][26] ),
    .X(_07669_));
 sky130_fd_sc_hd__clkbuf_1 _13860_ (.A(_07669_),
    .X(_00859_));
 sky130_fd_sc_hd__clkbuf_1 _13861_ (.A(\cpuregs.regs[0][27] ),
    .X(_07670_));
 sky130_fd_sc_hd__clkbuf_1 _13862_ (.A(_07670_),
    .X(_00860_));
 sky130_fd_sc_hd__clkbuf_1 _13863_ (.A(\cpuregs.regs[0][28] ),
    .X(_07671_));
 sky130_fd_sc_hd__clkbuf_1 _13864_ (.A(_07671_),
    .X(_00861_));
 sky130_fd_sc_hd__clkbuf_1 _13865_ (.A(\cpuregs.regs[0][29] ),
    .X(_07672_));
 sky130_fd_sc_hd__clkbuf_1 _13866_ (.A(_07672_),
    .X(_00862_));
 sky130_fd_sc_hd__clkbuf_1 _13867_ (.A(\cpuregs.regs[0][30] ),
    .X(_07673_));
 sky130_fd_sc_hd__clkbuf_1 _13868_ (.A(_07673_),
    .X(_00863_));
 sky130_fd_sc_hd__clkbuf_1 _13869_ (.A(\cpuregs.regs[0][31] ),
    .X(_07674_));
 sky130_fd_sc_hd__clkbuf_1 _13870_ (.A(_07674_),
    .X(_00864_));
 sky130_fd_sc_hd__buf_4 _13871_ (.A(_06053_),
    .X(_07675_));
 sky130_fd_sc_hd__nand2_1 _13872_ (.A(_06072_),
    .B(_03298_),
    .Y(_07676_));
 sky130_fd_sc_hd__nor2_2 _13873_ (.A(_03301_),
    .B(_07676_),
    .Y(_07677_));
 sky130_fd_sc_hd__buf_2 _13874_ (.A(_07677_),
    .X(_07678_));
 sky130_fd_sc_hd__nand2_2 _13875_ (.A(_03292_),
    .B(\cpu_state[2] ),
    .Y(_07679_));
 sky130_fd_sc_hd__nor2_1 _13876_ (.A(_03271_),
    .B(instr_retirq),
    .Y(_07680_));
 sky130_fd_sc_hd__a21o_2 _13877_ (.A1(_07676_),
    .A2(_07679_),
    .B1(_07680_),
    .X(_07681_));
 sky130_fd_sc_hd__buf_2 _13878_ (.A(_07681_),
    .X(_07682_));
 sky130_fd_sc_hd__a22o_1 _13879_ (.A1(_03338_),
    .A2(_07678_),
    .B1(_07682_),
    .B2(net131),
    .X(_07683_));
 sky130_fd_sc_hd__and2_1 _13880_ (.A(_07675_),
    .B(_07683_),
    .X(_07684_));
 sky130_fd_sc_hd__clkbuf_1 _13881_ (.A(_07684_),
    .X(_00866_));
 sky130_fd_sc_hd__a22o_1 _13882_ (.A1(_03351_),
    .A2(_07678_),
    .B1(_07682_),
    .B2(net142),
    .X(_07685_));
 sky130_fd_sc_hd__and2_1 _13883_ (.A(_07675_),
    .B(_07685_),
    .X(_07686_));
 sky130_fd_sc_hd__clkbuf_1 _13884_ (.A(_07686_),
    .X(_00867_));
 sky130_fd_sc_hd__a22o_1 _13885_ (.A1(_03326_),
    .A2(_07678_),
    .B1(_07682_),
    .B2(net153),
    .X(_07687_));
 sky130_fd_sc_hd__and2_1 _13886_ (.A(_07675_),
    .B(_07687_),
    .X(_07688_));
 sky130_fd_sc_hd__clkbuf_1 _13887_ (.A(_07688_),
    .X(_00868_));
 sky130_fd_sc_hd__a22o_1 _13888_ (.A1(_03344_),
    .A2(_07678_),
    .B1(_07682_),
    .B2(net156),
    .X(_07689_));
 sky130_fd_sc_hd__and2_1 _13889_ (.A(_07675_),
    .B(_07689_),
    .X(_07690_));
 sky130_fd_sc_hd__clkbuf_1 _13890_ (.A(_07690_),
    .X(_00869_));
 sky130_fd_sc_hd__clkbuf_2 _13891_ (.A(_06053_),
    .X(_07691_));
 sky130_fd_sc_hd__a22o_1 _13892_ (.A1(_03327_),
    .A2(_07678_),
    .B1(_07682_),
    .B2(net157),
    .X(_07692_));
 sky130_fd_sc_hd__and2_1 _13893_ (.A(_07691_),
    .B(_07692_),
    .X(_07693_));
 sky130_fd_sc_hd__clkbuf_1 _13894_ (.A(_07693_),
    .X(_00870_));
 sky130_fd_sc_hd__a22o_1 _13895_ (.A1(_03322_),
    .A2(_07678_),
    .B1(_07682_),
    .B2(net158),
    .X(_07694_));
 sky130_fd_sc_hd__and2_1 _13896_ (.A(_07691_),
    .B(_07694_),
    .X(_07695_));
 sky130_fd_sc_hd__clkbuf_1 _13897_ (.A(_07695_),
    .X(_00871_));
 sky130_fd_sc_hd__a22o_1 _13898_ (.A1(_03321_),
    .A2(_07678_),
    .B1(_07682_),
    .B2(net159),
    .X(_07696_));
 sky130_fd_sc_hd__and2_1 _13899_ (.A(_07691_),
    .B(_07696_),
    .X(_07697_));
 sky130_fd_sc_hd__clkbuf_1 _13900_ (.A(_07697_),
    .X(_00872_));
 sky130_fd_sc_hd__a22o_1 _13901_ (.A1(_03349_),
    .A2(_07678_),
    .B1(_07682_),
    .B2(net160),
    .X(_07698_));
 sky130_fd_sc_hd__and2_1 _13902_ (.A(_07691_),
    .B(_07698_),
    .X(_07699_));
 sky130_fd_sc_hd__clkbuf_1 _13903_ (.A(_07699_),
    .X(_00873_));
 sky130_fd_sc_hd__a22o_1 _13904_ (.A1(_03359_),
    .A2(_07678_),
    .B1(_07682_),
    .B2(net161),
    .X(_07700_));
 sky130_fd_sc_hd__and2_1 _13905_ (.A(_07691_),
    .B(_07700_),
    .X(_07701_));
 sky130_fd_sc_hd__clkbuf_1 _13906_ (.A(_07701_),
    .X(_00874_));
 sky130_fd_sc_hd__a22o_1 _13907_ (.A1(_03323_),
    .A2(_07678_),
    .B1(_07682_),
    .B2(net162),
    .X(_07702_));
 sky130_fd_sc_hd__and2_1 _13908_ (.A(_07691_),
    .B(_07702_),
    .X(_07703_));
 sky130_fd_sc_hd__clkbuf_1 _13909_ (.A(_07703_),
    .X(_00875_));
 sky130_fd_sc_hd__buf_2 _13910_ (.A(_07677_),
    .X(_07704_));
 sky130_fd_sc_hd__buf_2 _13911_ (.A(_07681_),
    .X(_07705_));
 sky130_fd_sc_hd__a22o_1 _13912_ (.A1(_03333_),
    .A2(_07704_),
    .B1(_07705_),
    .B2(net132),
    .X(_07706_));
 sky130_fd_sc_hd__and2_1 _13913_ (.A(_07691_),
    .B(_07706_),
    .X(_07707_));
 sky130_fd_sc_hd__clkbuf_1 _13914_ (.A(_07707_),
    .X(_00876_));
 sky130_fd_sc_hd__a22o_1 _13915_ (.A1(_03335_),
    .A2(_07704_),
    .B1(_07705_),
    .B2(net133),
    .X(_07708_));
 sky130_fd_sc_hd__and2_1 _13916_ (.A(_07691_),
    .B(_07708_),
    .X(_07709_));
 sky130_fd_sc_hd__clkbuf_1 _13917_ (.A(_07709_),
    .X(_00877_));
 sky130_fd_sc_hd__a22o_1 _13918_ (.A1(_03357_),
    .A2(_07704_),
    .B1(_07705_),
    .B2(net134),
    .X(_07710_));
 sky130_fd_sc_hd__and2_1 _13919_ (.A(_07691_),
    .B(_07710_),
    .X(_07711_));
 sky130_fd_sc_hd__clkbuf_1 _13920_ (.A(_07711_),
    .X(_00878_));
 sky130_fd_sc_hd__a22o_1 _13921_ (.A1(_03352_),
    .A2(_07704_),
    .B1(_07705_),
    .B2(net135),
    .X(_07712_));
 sky130_fd_sc_hd__and2_1 _13922_ (.A(_07691_),
    .B(_07712_),
    .X(_07713_));
 sky130_fd_sc_hd__clkbuf_1 _13923_ (.A(_07713_),
    .X(_00879_));
 sky130_fd_sc_hd__clkbuf_2 _13924_ (.A(_06053_),
    .X(_07714_));
 sky130_fd_sc_hd__a22o_1 _13925_ (.A1(_03353_),
    .A2(_07704_),
    .B1(_07705_),
    .B2(net136),
    .X(_07715_));
 sky130_fd_sc_hd__and2_1 _13926_ (.A(_07714_),
    .B(_07715_),
    .X(_07716_));
 sky130_fd_sc_hd__clkbuf_1 _13927_ (.A(_07716_),
    .X(_00880_));
 sky130_fd_sc_hd__a22o_1 _13928_ (.A1(_03356_),
    .A2(_07704_),
    .B1(_07705_),
    .B2(net137),
    .X(_07717_));
 sky130_fd_sc_hd__and2_1 _13929_ (.A(_07714_),
    .B(_07717_),
    .X(_07718_));
 sky130_fd_sc_hd__clkbuf_1 _13930_ (.A(_07718_),
    .X(_00881_));
 sky130_fd_sc_hd__a22o_1 _13931_ (.A1(_03330_),
    .A2(_07704_),
    .B1(_07705_),
    .B2(net138),
    .X(_07719_));
 sky130_fd_sc_hd__and2_1 _13932_ (.A(_07714_),
    .B(_07719_),
    .X(_07720_));
 sky130_fd_sc_hd__clkbuf_1 _13933_ (.A(_07720_),
    .X(_00882_));
 sky130_fd_sc_hd__a22o_1 _13934_ (.A1(_03348_),
    .A2(_07704_),
    .B1(_07705_),
    .B2(net139),
    .X(_07721_));
 sky130_fd_sc_hd__and2_1 _13935_ (.A(_07714_),
    .B(_07721_),
    .X(_07722_));
 sky130_fd_sc_hd__clkbuf_1 _13936_ (.A(_07722_),
    .X(_00883_));
 sky130_fd_sc_hd__a22o_1 _13937_ (.A1(_03336_),
    .A2(_07704_),
    .B1(_07705_),
    .B2(net140),
    .X(_07723_));
 sky130_fd_sc_hd__and2_1 _13938_ (.A(_07714_),
    .B(_07723_),
    .X(_07724_));
 sky130_fd_sc_hd__clkbuf_1 _13939_ (.A(_07724_),
    .X(_00884_));
 sky130_fd_sc_hd__a22o_1 _13940_ (.A1(_03358_),
    .A2(_07704_),
    .B1(_07705_),
    .B2(net141),
    .X(_07725_));
 sky130_fd_sc_hd__and2_1 _13941_ (.A(_07714_),
    .B(_07725_),
    .X(_07726_));
 sky130_fd_sc_hd__clkbuf_1 _13942_ (.A(_07726_),
    .X(_00885_));
 sky130_fd_sc_hd__buf_2 _13943_ (.A(_07677_),
    .X(_07727_));
 sky130_fd_sc_hd__buf_2 _13944_ (.A(_07681_),
    .X(_07728_));
 sky130_fd_sc_hd__a22o_1 _13945_ (.A1(_03332_),
    .A2(_07727_),
    .B1(_07728_),
    .B2(net143),
    .X(_07729_));
 sky130_fd_sc_hd__and2_1 _13946_ (.A(_07714_),
    .B(_07729_),
    .X(_07730_));
 sky130_fd_sc_hd__clkbuf_1 _13947_ (.A(_07730_),
    .X(_00886_));
 sky130_fd_sc_hd__a22o_1 _13948_ (.A1(_03346_),
    .A2(_07727_),
    .B1(_07728_),
    .B2(net144),
    .X(_07731_));
 sky130_fd_sc_hd__and2_1 _13949_ (.A(_07714_),
    .B(_07731_),
    .X(_07732_));
 sky130_fd_sc_hd__clkbuf_1 _13950_ (.A(_07732_),
    .X(_00887_));
 sky130_fd_sc_hd__a22o_1 _13951_ (.A1(_03320_),
    .A2(_07727_),
    .B1(_07728_),
    .B2(net145),
    .X(_07733_));
 sky130_fd_sc_hd__and2_1 _13952_ (.A(_07714_),
    .B(_07733_),
    .X(_07734_));
 sky130_fd_sc_hd__clkbuf_1 _13953_ (.A(_07734_),
    .X(_00888_));
 sky130_fd_sc_hd__a22o_1 _13954_ (.A1(_03343_),
    .A2(_07727_),
    .B1(_07728_),
    .B2(net146),
    .X(_07735_));
 sky130_fd_sc_hd__and2_1 _13955_ (.A(_07714_),
    .B(_07735_),
    .X(_07736_));
 sky130_fd_sc_hd__clkbuf_1 _13956_ (.A(_07736_),
    .X(_00889_));
 sky130_fd_sc_hd__buf_4 _13957_ (.A(_03304_),
    .X(_07737_));
 sky130_fd_sc_hd__a22o_1 _13958_ (.A1(_03342_),
    .A2(_07727_),
    .B1(_07728_),
    .B2(net147),
    .X(_07738_));
 sky130_fd_sc_hd__and2_1 _13959_ (.A(_07737_),
    .B(_07738_),
    .X(_07739_));
 sky130_fd_sc_hd__clkbuf_1 _13960_ (.A(_07739_),
    .X(_00890_));
 sky130_fd_sc_hd__a22o_1 _13961_ (.A1(_03347_),
    .A2(_07727_),
    .B1(_07728_),
    .B2(net148),
    .X(_07740_));
 sky130_fd_sc_hd__and2_1 _13962_ (.A(_07737_),
    .B(_07740_),
    .X(_07741_));
 sky130_fd_sc_hd__clkbuf_1 _13963_ (.A(_07741_),
    .X(_00891_));
 sky130_fd_sc_hd__a22o_1 _13964_ (.A1(_03325_),
    .A2(_07727_),
    .B1(_07728_),
    .B2(net149),
    .X(_07742_));
 sky130_fd_sc_hd__and2_1 _13965_ (.A(_07737_),
    .B(_07742_),
    .X(_07743_));
 sky130_fd_sc_hd__clkbuf_1 _13966_ (.A(_07743_),
    .X(_00892_));
 sky130_fd_sc_hd__a22o_1 _13967_ (.A1(_03341_),
    .A2(_07727_),
    .B1(_07728_),
    .B2(net150),
    .X(_07744_));
 sky130_fd_sc_hd__and2_1 _13968_ (.A(_07737_),
    .B(_07744_),
    .X(_07745_));
 sky130_fd_sc_hd__clkbuf_1 _13969_ (.A(_07745_),
    .X(_00893_));
 sky130_fd_sc_hd__a22o_1 _13970_ (.A1(_03354_),
    .A2(_07727_),
    .B1(_07728_),
    .B2(net151),
    .X(_07746_));
 sky130_fd_sc_hd__and2_1 _13971_ (.A(_07737_),
    .B(_07746_),
    .X(_07747_));
 sky130_fd_sc_hd__clkbuf_1 _13972_ (.A(_07747_),
    .X(_00894_));
 sky130_fd_sc_hd__a22o_1 _13973_ (.A1(_03337_),
    .A2(_07727_),
    .B1(_07728_),
    .B2(net152),
    .X(_07748_));
 sky130_fd_sc_hd__and2_1 _13974_ (.A(_07737_),
    .B(_07748_),
    .X(_07749_));
 sky130_fd_sc_hd__clkbuf_1 _13975_ (.A(_07749_),
    .X(_00895_));
 sky130_fd_sc_hd__a22o_1 _13976_ (.A1(_03328_),
    .A2(_07677_),
    .B1(_07681_),
    .B2(net154),
    .X(_07750_));
 sky130_fd_sc_hd__and2_1 _13977_ (.A(_07737_),
    .B(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__clkbuf_1 _13978_ (.A(_07751_),
    .X(_00896_));
 sky130_fd_sc_hd__a22o_1 _13979_ (.A1(_03331_),
    .A2(_07677_),
    .B1(_07681_),
    .B2(net155),
    .X(_07752_));
 sky130_fd_sc_hd__and2_1 _13980_ (.A(_07737_),
    .B(_07752_),
    .X(_07753_));
 sky130_fd_sc_hd__clkbuf_1 _13981_ (.A(_07753_),
    .X(_00897_));
 sky130_fd_sc_hd__and2b_2 _13982_ (.A_N(instr_waitirq),
    .B(decoder_trigger),
    .X(_07754_));
 sky130_fd_sc_hd__and4b_2 _13983_ (.A_N(_03363_),
    .B(_07754_),
    .C(\cpu_state[1] ),
    .D(_03376_),
    .X(_07755_));
 sky130_fd_sc_hd__and2_1 _13984_ (.A(\count_instr[0] ),
    .B(_07755_),
    .X(_07756_));
 sky130_fd_sc_hd__o21ai_1 _13985_ (.A1(\count_instr[0] ),
    .A2(_07755_),
    .B1(_06054_),
    .Y(_07757_));
 sky130_fd_sc_hd__nor2_1 _13986_ (.A(_07756_),
    .B(_07757_),
    .Y(_00898_));
 sky130_fd_sc_hd__and3_1 _13987_ (.A(\count_instr[1] ),
    .B(\count_instr[0] ),
    .C(_07755_),
    .X(_07758_));
 sky130_fd_sc_hd__clkbuf_4 _13988_ (.A(_06053_),
    .X(_07759_));
 sky130_fd_sc_hd__o21ai_1 _13989_ (.A1(\count_instr[1] ),
    .A2(_07756_),
    .B1(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__nor2_1 _13990_ (.A(_07758_),
    .B(_07760_),
    .Y(_00899_));
 sky130_fd_sc_hd__and4_1 _13991_ (.A(\count_instr[2] ),
    .B(\count_instr[1] ),
    .C(\count_instr[0] ),
    .D(_07755_),
    .X(_07761_));
 sky130_fd_sc_hd__o21ai_1 _13992_ (.A1(\count_instr[2] ),
    .A2(_07758_),
    .B1(_07759_),
    .Y(_07762_));
 sky130_fd_sc_hd__nor2_1 _13993_ (.A(_07761_),
    .B(_07762_),
    .Y(_00900_));
 sky130_fd_sc_hd__and2_1 _13994_ (.A(\count_instr[3] ),
    .B(_07761_),
    .X(_07763_));
 sky130_fd_sc_hd__o21ai_1 _13995_ (.A1(\count_instr[3] ),
    .A2(_07761_),
    .B1(_07759_),
    .Y(_07764_));
 sky130_fd_sc_hd__nor2_1 _13996_ (.A(_07763_),
    .B(_07764_),
    .Y(_00901_));
 sky130_fd_sc_hd__and3_1 _13997_ (.A(\count_instr[4] ),
    .B(\count_instr[3] ),
    .C(_07761_),
    .X(_07765_));
 sky130_fd_sc_hd__o21ai_1 _13998_ (.A1(\count_instr[4] ),
    .A2(_07763_),
    .B1(_07759_),
    .Y(_07766_));
 sky130_fd_sc_hd__nor2_1 _13999_ (.A(_07765_),
    .B(_07766_),
    .Y(_00902_));
 sky130_fd_sc_hd__and4_1 _14000_ (.A(\count_instr[5] ),
    .B(\count_instr[4] ),
    .C(\count_instr[3] ),
    .D(_07761_),
    .X(_07767_));
 sky130_fd_sc_hd__o21ai_1 _14001_ (.A1(\count_instr[5] ),
    .A2(_07765_),
    .B1(_07759_),
    .Y(_07768_));
 sky130_fd_sc_hd__nor2_1 _14002_ (.A(_07767_),
    .B(_07768_),
    .Y(_00903_));
 sky130_fd_sc_hd__and2_1 _14003_ (.A(\count_instr[6] ),
    .B(_07767_),
    .X(_07769_));
 sky130_fd_sc_hd__o21ai_1 _14004_ (.A1(\count_instr[6] ),
    .A2(_07767_),
    .B1(_07759_),
    .Y(_07770_));
 sky130_fd_sc_hd__nor2_1 _14005_ (.A(_07769_),
    .B(_07770_),
    .Y(_00904_));
 sky130_fd_sc_hd__and3_1 _14006_ (.A(\count_instr[7] ),
    .B(\count_instr[6] ),
    .C(_07767_),
    .X(_07771_));
 sky130_fd_sc_hd__o21ai_1 _14007_ (.A1(\count_instr[7] ),
    .A2(_07769_),
    .B1(_07759_),
    .Y(_07772_));
 sky130_fd_sc_hd__nor2_1 _14008_ (.A(_07771_),
    .B(_07772_),
    .Y(_00905_));
 sky130_fd_sc_hd__and4_2 _14009_ (.A(\count_instr[8] ),
    .B(\count_instr[7] ),
    .C(\count_instr[6] ),
    .D(_07767_),
    .X(_07773_));
 sky130_fd_sc_hd__o21ai_1 _14010_ (.A1(\count_instr[8] ),
    .A2(_07771_),
    .B1(_07759_),
    .Y(_07774_));
 sky130_fd_sc_hd__nor2_1 _14011_ (.A(_07773_),
    .B(_07774_),
    .Y(_00906_));
 sky130_fd_sc_hd__buf_4 _14012_ (.A(_03239_),
    .X(_07775_));
 sky130_fd_sc_hd__a21oi_1 _14013_ (.A1(\count_instr[9] ),
    .A2(_07773_),
    .B1(_07775_),
    .Y(_07776_));
 sky130_fd_sc_hd__o21a_1 _14014_ (.A1(\count_instr[9] ),
    .A2(_07773_),
    .B1(_07776_),
    .X(_00907_));
 sky130_fd_sc_hd__and3_1 _14015_ (.A(\count_instr[10] ),
    .B(\count_instr[9] ),
    .C(_07773_),
    .X(_07777_));
 sky130_fd_sc_hd__clkbuf_8 _14016_ (.A(_03304_),
    .X(_07778_));
 sky130_fd_sc_hd__a21o_1 _14017_ (.A1(\count_instr[9] ),
    .A2(_07773_),
    .B1(\count_instr[10] ),
    .X(_07779_));
 sky130_fd_sc_hd__and3b_1 _14018_ (.A_N(_07777_),
    .B(_07778_),
    .C(_07779_),
    .X(_07780_));
 sky130_fd_sc_hd__clkbuf_1 _14019_ (.A(_07780_),
    .X(_00908_));
 sky130_fd_sc_hd__and4_2 _14020_ (.A(\count_instr[11] ),
    .B(\count_instr[10] ),
    .C(\count_instr[9] ),
    .D(_07773_),
    .X(_07781_));
 sky130_fd_sc_hd__o21ai_1 _14021_ (.A1(\count_instr[11] ),
    .A2(_07777_),
    .B1(_07759_),
    .Y(_07782_));
 sky130_fd_sc_hd__nor2_1 _14022_ (.A(_07781_),
    .B(_07782_),
    .Y(_00909_));
 sky130_fd_sc_hd__a21oi_1 _14023_ (.A1(\count_instr[12] ),
    .A2(_07781_),
    .B1(_07775_),
    .Y(_07783_));
 sky130_fd_sc_hd__o21a_1 _14024_ (.A1(\count_instr[12] ),
    .A2(_07781_),
    .B1(_07783_),
    .X(_00910_));
 sky130_fd_sc_hd__and3_1 _14025_ (.A(\count_instr[13] ),
    .B(\count_instr[12] ),
    .C(_07781_),
    .X(_07784_));
 sky130_fd_sc_hd__a21o_1 _14026_ (.A1(\count_instr[12] ),
    .A2(_07781_),
    .B1(\count_instr[13] ),
    .X(_07785_));
 sky130_fd_sc_hd__and3b_1 _14027_ (.A_N(_07784_),
    .B(_07778_),
    .C(_07785_),
    .X(_07786_));
 sky130_fd_sc_hd__clkbuf_1 _14028_ (.A(_07786_),
    .X(_00911_));
 sky130_fd_sc_hd__and4_1 _14029_ (.A(\count_instr[14] ),
    .B(\count_instr[13] ),
    .C(\count_instr[12] ),
    .D(_07781_),
    .X(_07787_));
 sky130_fd_sc_hd__o21ai_1 _14030_ (.A1(\count_instr[14] ),
    .A2(_07784_),
    .B1(_07759_),
    .Y(_07788_));
 sky130_fd_sc_hd__nor2_1 _14031_ (.A(_07787_),
    .B(_07788_),
    .Y(_00912_));
 sky130_fd_sc_hd__and2_1 _14032_ (.A(\count_instr[15] ),
    .B(_07787_),
    .X(_07789_));
 sky130_fd_sc_hd__clkbuf_4 _14033_ (.A(_06053_),
    .X(_07790_));
 sky130_fd_sc_hd__o21ai_1 _14034_ (.A1(\count_instr[15] ),
    .A2(_07787_),
    .B1(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__nor2_1 _14035_ (.A(_07789_),
    .B(_07791_),
    .Y(_00913_));
 sky130_fd_sc_hd__and3_1 _14036_ (.A(\count_instr[16] ),
    .B(\count_instr[15] ),
    .C(_07787_),
    .X(_07792_));
 sky130_fd_sc_hd__o21ai_1 _14037_ (.A1(\count_instr[16] ),
    .A2(_07789_),
    .B1(_07790_),
    .Y(_07793_));
 sky130_fd_sc_hd__nor2_1 _14038_ (.A(_07792_),
    .B(_07793_),
    .Y(_00914_));
 sky130_fd_sc_hd__o21ai_1 _14039_ (.A1(\count_instr[17] ),
    .A2(_07792_),
    .B1(_07675_),
    .Y(_07794_));
 sky130_fd_sc_hd__a21oi_1 _14040_ (.A1(\count_instr[17] ),
    .A2(_07792_),
    .B1(_07794_),
    .Y(_00915_));
 sky130_fd_sc_hd__and3_1 _14041_ (.A(\count_instr[18] ),
    .B(\count_instr[17] ),
    .C(\count_instr[16] ),
    .X(_07795_));
 sky130_fd_sc_hd__and3_1 _14042_ (.A(\count_instr[15] ),
    .B(_07787_),
    .C(_07795_),
    .X(_07796_));
 sky130_fd_sc_hd__a21o_1 _14043_ (.A1(\count_instr[17] ),
    .A2(_07792_),
    .B1(\count_instr[18] ),
    .X(_07797_));
 sky130_fd_sc_hd__and3b_1 _14044_ (.A_N(_07796_),
    .B(_07778_),
    .C(_07797_),
    .X(_07798_));
 sky130_fd_sc_hd__clkbuf_1 _14045_ (.A(_07798_),
    .X(_00916_));
 sky130_fd_sc_hd__and4_1 _14046_ (.A(\count_instr[19] ),
    .B(\count_instr[15] ),
    .C(_07787_),
    .D(_07795_),
    .X(_07799_));
 sky130_fd_sc_hd__o21ai_1 _14047_ (.A1(\count_instr[19] ),
    .A2(_07796_),
    .B1(_07790_),
    .Y(_07800_));
 sky130_fd_sc_hd__nor2_1 _14048_ (.A(_07799_),
    .B(_07800_),
    .Y(_00917_));
 sky130_fd_sc_hd__and2_1 _14049_ (.A(\count_instr[20] ),
    .B(_07799_),
    .X(_07801_));
 sky130_fd_sc_hd__o21ai_1 _14050_ (.A1(\count_instr[20] ),
    .A2(_07799_),
    .B1(_07790_),
    .Y(_07802_));
 sky130_fd_sc_hd__nor2_1 _14051_ (.A(_07801_),
    .B(_07802_),
    .Y(_00918_));
 sky130_fd_sc_hd__and3_1 _14052_ (.A(\count_instr[21] ),
    .B(\count_instr[20] ),
    .C(_07799_),
    .X(_07803_));
 sky130_fd_sc_hd__o21ai_1 _14053_ (.A1(\count_instr[21] ),
    .A2(_07801_),
    .B1(_07790_),
    .Y(_07804_));
 sky130_fd_sc_hd__nor2_1 _14054_ (.A(_07803_),
    .B(_07804_),
    .Y(_00919_));
 sky130_fd_sc_hd__and4_2 _14055_ (.A(\count_instr[22] ),
    .B(\count_instr[21] ),
    .C(\count_instr[20] ),
    .D(_07799_),
    .X(_07805_));
 sky130_fd_sc_hd__o21ai_1 _14056_ (.A1(\count_instr[22] ),
    .A2(_07803_),
    .B1(_07790_),
    .Y(_07806_));
 sky130_fd_sc_hd__nor2_1 _14057_ (.A(_07805_),
    .B(_07806_),
    .Y(_00920_));
 sky130_fd_sc_hd__a21oi_1 _14058_ (.A1(\count_instr[23] ),
    .A2(_07805_),
    .B1(_07775_),
    .Y(_07807_));
 sky130_fd_sc_hd__o21a_1 _14059_ (.A1(\count_instr[23] ),
    .A2(_07805_),
    .B1(_07807_),
    .X(_00921_));
 sky130_fd_sc_hd__and3_1 _14060_ (.A(\count_instr[24] ),
    .B(\count_instr[23] ),
    .C(_07805_),
    .X(_07808_));
 sky130_fd_sc_hd__a21o_1 _14061_ (.A1(\count_instr[23] ),
    .A2(_07805_),
    .B1(\count_instr[24] ),
    .X(_07809_));
 sky130_fd_sc_hd__and3b_1 _14062_ (.A_N(_07808_),
    .B(_07778_),
    .C(_07809_),
    .X(_07810_));
 sky130_fd_sc_hd__clkbuf_1 _14063_ (.A(_07810_),
    .X(_00922_));
 sky130_fd_sc_hd__and4_2 _14064_ (.A(\count_instr[25] ),
    .B(\count_instr[24] ),
    .C(\count_instr[23] ),
    .D(_07805_),
    .X(_07811_));
 sky130_fd_sc_hd__o21ai_1 _14065_ (.A1(\count_instr[25] ),
    .A2(_07808_),
    .B1(_07790_),
    .Y(_07812_));
 sky130_fd_sc_hd__nor2_1 _14066_ (.A(_07811_),
    .B(_07812_),
    .Y(_00923_));
 sky130_fd_sc_hd__a21oi_1 _14067_ (.A1(\count_instr[26] ),
    .A2(_07811_),
    .B1(_07775_),
    .Y(_07813_));
 sky130_fd_sc_hd__o21a_1 _14068_ (.A1(\count_instr[26] ),
    .A2(_07811_),
    .B1(_07813_),
    .X(_00924_));
 sky130_fd_sc_hd__and3_1 _14069_ (.A(\count_instr[27] ),
    .B(\count_instr[26] ),
    .C(_07811_),
    .X(_07814_));
 sky130_fd_sc_hd__clkbuf_4 _14070_ (.A(_03304_),
    .X(_07815_));
 sky130_fd_sc_hd__a21o_1 _14071_ (.A1(\count_instr[26] ),
    .A2(_07811_),
    .B1(\count_instr[27] ),
    .X(_07816_));
 sky130_fd_sc_hd__and3b_1 _14072_ (.A_N(_07814_),
    .B(_07815_),
    .C(_07816_),
    .X(_07817_));
 sky130_fd_sc_hd__clkbuf_1 _14073_ (.A(_07817_),
    .X(_00925_));
 sky130_fd_sc_hd__and4_2 _14074_ (.A(\count_instr[28] ),
    .B(\count_instr[27] ),
    .C(\count_instr[26] ),
    .D(_07811_),
    .X(_07818_));
 sky130_fd_sc_hd__o21ai_1 _14075_ (.A1(\count_instr[28] ),
    .A2(_07814_),
    .B1(_07790_),
    .Y(_07819_));
 sky130_fd_sc_hd__nor2_1 _14076_ (.A(_07818_),
    .B(_07819_),
    .Y(_00926_));
 sky130_fd_sc_hd__a21oi_1 _14077_ (.A1(\count_instr[29] ),
    .A2(_07818_),
    .B1(_07775_),
    .Y(_07820_));
 sky130_fd_sc_hd__o21a_1 _14078_ (.A1(\count_instr[29] ),
    .A2(_07818_),
    .B1(_07820_),
    .X(_00927_));
 sky130_fd_sc_hd__and3_1 _14079_ (.A(\count_instr[30] ),
    .B(\count_instr[29] ),
    .C(_07818_),
    .X(_07821_));
 sky130_fd_sc_hd__a21o_1 _14080_ (.A1(\count_instr[29] ),
    .A2(_07818_),
    .B1(\count_instr[30] ),
    .X(_07822_));
 sky130_fd_sc_hd__and3b_1 _14081_ (.A_N(_07821_),
    .B(_07815_),
    .C(_07822_),
    .X(_07823_));
 sky130_fd_sc_hd__clkbuf_1 _14082_ (.A(_07823_),
    .X(_00928_));
 sky130_fd_sc_hd__and4_2 _14083_ (.A(\count_instr[31] ),
    .B(\count_instr[30] ),
    .C(\count_instr[29] ),
    .D(_07818_),
    .X(_07824_));
 sky130_fd_sc_hd__o21ai_1 _14084_ (.A1(\count_instr[31] ),
    .A2(_07821_),
    .B1(_07790_),
    .Y(_07825_));
 sky130_fd_sc_hd__nor2_1 _14085_ (.A(_07824_),
    .B(_07825_),
    .Y(_00929_));
 sky130_fd_sc_hd__buf_4 _14086_ (.A(_03239_),
    .X(_07826_));
 sky130_fd_sc_hd__a21oi_1 _14087_ (.A1(\count_instr[32] ),
    .A2(_07824_),
    .B1(_07826_),
    .Y(_07827_));
 sky130_fd_sc_hd__o21a_1 _14088_ (.A1(\count_instr[32] ),
    .A2(_07824_),
    .B1(_07827_),
    .X(_00930_));
 sky130_fd_sc_hd__and3_1 _14089_ (.A(\count_instr[33] ),
    .B(\count_instr[32] ),
    .C(_07824_),
    .X(_07828_));
 sky130_fd_sc_hd__a21o_1 _14090_ (.A1(\count_instr[32] ),
    .A2(_07824_),
    .B1(\count_instr[33] ),
    .X(_07829_));
 sky130_fd_sc_hd__and3b_1 _14091_ (.A_N(_07828_),
    .B(_07815_),
    .C(_07829_),
    .X(_07830_));
 sky130_fd_sc_hd__clkbuf_1 _14092_ (.A(_07830_),
    .X(_00931_));
 sky130_fd_sc_hd__and4_2 _14093_ (.A(\count_instr[34] ),
    .B(\count_instr[33] ),
    .C(\count_instr[32] ),
    .D(_07824_),
    .X(_07831_));
 sky130_fd_sc_hd__o21ai_1 _14094_ (.A1(\count_instr[34] ),
    .A2(_07828_),
    .B1(_07790_),
    .Y(_07832_));
 sky130_fd_sc_hd__nor2_1 _14095_ (.A(_07831_),
    .B(_07832_),
    .Y(_00932_));
 sky130_fd_sc_hd__and2_1 _14096_ (.A(\count_instr[35] ),
    .B(_07831_),
    .X(_07833_));
 sky130_fd_sc_hd__clkbuf_4 _14097_ (.A(_06053_),
    .X(_07834_));
 sky130_fd_sc_hd__o21ai_1 _14098_ (.A1(\count_instr[35] ),
    .A2(_07831_),
    .B1(_07834_),
    .Y(_07835_));
 sky130_fd_sc_hd__nor2_1 _14099_ (.A(_07833_),
    .B(_07835_),
    .Y(_00933_));
 sky130_fd_sc_hd__and3_1 _14100_ (.A(\count_instr[36] ),
    .B(\count_instr[35] ),
    .C(_07831_),
    .X(_07836_));
 sky130_fd_sc_hd__o21ai_1 _14101_ (.A1(\count_instr[36] ),
    .A2(_07833_),
    .B1(_07834_),
    .Y(_07837_));
 sky130_fd_sc_hd__nor2_1 _14102_ (.A(_07836_),
    .B(_07837_),
    .Y(_00934_));
 sky130_fd_sc_hd__o21ai_1 _14103_ (.A1(\count_instr[37] ),
    .A2(_07836_),
    .B1(_07675_),
    .Y(_07838_));
 sky130_fd_sc_hd__a21oi_1 _14104_ (.A1(\count_instr[37] ),
    .A2(_07836_),
    .B1(_07838_),
    .Y(_00935_));
 sky130_fd_sc_hd__and3_1 _14105_ (.A(\count_instr[38] ),
    .B(\count_instr[37] ),
    .C(\count_instr[36] ),
    .X(_07839_));
 sky130_fd_sc_hd__and3_1 _14106_ (.A(\count_instr[35] ),
    .B(_07831_),
    .C(_07839_),
    .X(_07840_));
 sky130_fd_sc_hd__a21o_1 _14107_ (.A1(\count_instr[37] ),
    .A2(_07836_),
    .B1(\count_instr[38] ),
    .X(_07841_));
 sky130_fd_sc_hd__and3b_1 _14108_ (.A_N(_07840_),
    .B(_07815_),
    .C(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__clkbuf_1 _14109_ (.A(_07842_),
    .X(_00936_));
 sky130_fd_sc_hd__and4_2 _14110_ (.A(\count_instr[39] ),
    .B(\count_instr[35] ),
    .C(_07831_),
    .D(_07839_),
    .X(_07843_));
 sky130_fd_sc_hd__o21ai_1 _14111_ (.A1(\count_instr[39] ),
    .A2(_07840_),
    .B1(_07834_),
    .Y(_07844_));
 sky130_fd_sc_hd__nor2_1 _14112_ (.A(_07843_),
    .B(_07844_),
    .Y(_00937_));
 sky130_fd_sc_hd__and2_1 _14113_ (.A(\count_instr[40] ),
    .B(_07843_),
    .X(_07845_));
 sky130_fd_sc_hd__o21ai_1 _14114_ (.A1(\count_instr[40] ),
    .A2(_07843_),
    .B1(_07834_),
    .Y(_07846_));
 sky130_fd_sc_hd__nor2_1 _14115_ (.A(_07845_),
    .B(_07846_),
    .Y(_00938_));
 sky130_fd_sc_hd__o21ai_1 _14116_ (.A1(\count_instr[41] ),
    .A2(_07845_),
    .B1(_07675_),
    .Y(_07847_));
 sky130_fd_sc_hd__a21oi_1 _14117_ (.A1(\count_instr[41] ),
    .A2(_07845_),
    .B1(_07847_),
    .Y(_00939_));
 sky130_fd_sc_hd__and3_1 _14118_ (.A(\count_instr[42] ),
    .B(\count_instr[41] ),
    .C(\count_instr[40] ),
    .X(_07848_));
 sky130_fd_sc_hd__and2_1 _14119_ (.A(_07843_),
    .B(_07848_),
    .X(_07849_));
 sky130_fd_sc_hd__a31o_1 _14120_ (.A1(\count_instr[41] ),
    .A2(\count_instr[40] ),
    .A3(_07843_),
    .B1(\count_instr[42] ),
    .X(_07850_));
 sky130_fd_sc_hd__and3b_1 _14121_ (.A_N(_07849_),
    .B(_07815_),
    .C(_07850_),
    .X(_07851_));
 sky130_fd_sc_hd__clkbuf_1 _14122_ (.A(_07851_),
    .X(_00940_));
 sky130_fd_sc_hd__and3_1 _14123_ (.A(\count_instr[43] ),
    .B(_07843_),
    .C(_07848_),
    .X(_07852_));
 sky130_fd_sc_hd__o21ai_1 _14124_ (.A1(\count_instr[43] ),
    .A2(_07849_),
    .B1(_07834_),
    .Y(_07853_));
 sky130_fd_sc_hd__nor2_1 _14125_ (.A(_07852_),
    .B(_07853_),
    .Y(_00941_));
 sky130_fd_sc_hd__or2_1 _14126_ (.A(\count_instr[44] ),
    .B(_07852_),
    .X(_07854_));
 sky130_fd_sc_hd__nand2_1 _14127_ (.A(\count_instr[44] ),
    .B(_07852_),
    .Y(_07855_));
 sky130_fd_sc_hd__and3_1 _14128_ (.A(_07778_),
    .B(_07854_),
    .C(_07855_),
    .X(_07856_));
 sky130_fd_sc_hd__clkbuf_1 _14129_ (.A(_07856_),
    .X(_00942_));
 sky130_fd_sc_hd__inv_2 _14130_ (.A(\count_instr[45] ),
    .Y(_07857_));
 sky130_fd_sc_hd__and2_1 _14131_ (.A(\count_instr[45] ),
    .B(\count_instr[44] ),
    .X(_07858_));
 sky130_fd_sc_hd__and4_1 _14132_ (.A(\count_instr[43] ),
    .B(_07843_),
    .C(_07848_),
    .D(_07858_),
    .X(_07859_));
 sky130_fd_sc_hd__a211oi_1 _14133_ (.A1(_07857_),
    .A2(_07855_),
    .B1(_07859_),
    .C1(_07775_),
    .Y(_00943_));
 sky130_fd_sc_hd__and2_1 _14134_ (.A(\count_instr[46] ),
    .B(_07859_),
    .X(_07860_));
 sky130_fd_sc_hd__o21ai_1 _14135_ (.A1(\count_instr[46] ),
    .A2(_07859_),
    .B1(_07834_),
    .Y(_07861_));
 sky130_fd_sc_hd__nor2_1 _14136_ (.A(_07860_),
    .B(_07861_),
    .Y(_00944_));
 sky130_fd_sc_hd__and3_1 _14137_ (.A(\count_instr[47] ),
    .B(\count_instr[46] ),
    .C(_07859_),
    .X(_07862_));
 sky130_fd_sc_hd__o21ai_1 _14138_ (.A1(\count_instr[47] ),
    .A2(_07860_),
    .B1(_07834_),
    .Y(_07863_));
 sky130_fd_sc_hd__nor2_1 _14139_ (.A(_07862_),
    .B(_07863_),
    .Y(_00945_));
 sky130_fd_sc_hd__and4_1 _14140_ (.A(\count_instr[48] ),
    .B(\count_instr[47] ),
    .C(\count_instr[46] ),
    .D(_07859_),
    .X(_07864_));
 sky130_fd_sc_hd__clkbuf_2 _14141_ (.A(_07864_),
    .X(_07865_));
 sky130_fd_sc_hd__o21ai_1 _14142_ (.A1(\count_instr[48] ),
    .A2(_07862_),
    .B1(_07834_),
    .Y(_07866_));
 sky130_fd_sc_hd__nor2_1 _14143_ (.A(_07865_),
    .B(_07866_),
    .Y(_00946_));
 sky130_fd_sc_hd__a21oi_1 _14144_ (.A1(\count_instr[49] ),
    .A2(_07865_),
    .B1(_07826_),
    .Y(_07867_));
 sky130_fd_sc_hd__o21a_1 _14145_ (.A1(\count_instr[49] ),
    .A2(_07865_),
    .B1(_07867_),
    .X(_00947_));
 sky130_fd_sc_hd__and2_1 _14146_ (.A(\count_instr[50] ),
    .B(\count_instr[49] ),
    .X(_07868_));
 sky130_fd_sc_hd__and2_1 _14147_ (.A(_07865_),
    .B(_07868_),
    .X(_07869_));
 sky130_fd_sc_hd__a21o_1 _14148_ (.A1(\count_instr[49] ),
    .A2(_07865_),
    .B1(\count_instr[50] ),
    .X(_07870_));
 sky130_fd_sc_hd__and3b_1 _14149_ (.A_N(_07869_),
    .B(_07815_),
    .C(_07870_),
    .X(_07871_));
 sky130_fd_sc_hd__clkbuf_1 _14150_ (.A(_07871_),
    .X(_00948_));
 sky130_fd_sc_hd__and3_1 _14151_ (.A(\count_instr[51] ),
    .B(_07865_),
    .C(_07868_),
    .X(_07872_));
 sky130_fd_sc_hd__o21ai_1 _14152_ (.A1(\count_instr[51] ),
    .A2(_07869_),
    .B1(_07834_),
    .Y(_07873_));
 sky130_fd_sc_hd__nor2_1 _14153_ (.A(_07872_),
    .B(_07873_),
    .Y(_00949_));
 sky130_fd_sc_hd__and4_1 _14154_ (.A(\count_instr[52] ),
    .B(\count_instr[51] ),
    .C(_07865_),
    .D(_07868_),
    .X(_07874_));
 sky130_fd_sc_hd__o21ai_1 _14155_ (.A1(\count_instr[52] ),
    .A2(_07872_),
    .B1(_07834_),
    .Y(_07875_));
 sky130_fd_sc_hd__nor2_1 _14156_ (.A(_07874_),
    .B(_07875_),
    .Y(_00950_));
 sky130_fd_sc_hd__and2_1 _14157_ (.A(\count_instr[53] ),
    .B(_07874_),
    .X(_07876_));
 sky130_fd_sc_hd__clkbuf_4 _14158_ (.A(_06053_),
    .X(_07877_));
 sky130_fd_sc_hd__o21ai_1 _14159_ (.A1(\count_instr[53] ),
    .A2(_07874_),
    .B1(_07877_),
    .Y(_07878_));
 sky130_fd_sc_hd__nor2_1 _14160_ (.A(_07876_),
    .B(_07878_),
    .Y(_00951_));
 sky130_fd_sc_hd__and3_1 _14161_ (.A(\count_instr[54] ),
    .B(\count_instr[53] ),
    .C(_07874_),
    .X(_07879_));
 sky130_fd_sc_hd__o21ai_1 _14162_ (.A1(\count_instr[54] ),
    .A2(_07876_),
    .B1(_07877_),
    .Y(_07880_));
 sky130_fd_sc_hd__nor2_1 _14163_ (.A(_07879_),
    .B(_07880_),
    .Y(_00952_));
 sky130_fd_sc_hd__and4_2 _14164_ (.A(\count_instr[55] ),
    .B(\count_instr[54] ),
    .C(\count_instr[53] ),
    .D(_07874_),
    .X(_07881_));
 sky130_fd_sc_hd__o21ai_1 _14165_ (.A1(\count_instr[55] ),
    .A2(_07879_),
    .B1(_07877_),
    .Y(_07882_));
 sky130_fd_sc_hd__nor2_1 _14166_ (.A(_07881_),
    .B(_07882_),
    .Y(_00953_));
 sky130_fd_sc_hd__a21oi_1 _14167_ (.A1(\count_instr[56] ),
    .A2(_07881_),
    .B1(_07826_),
    .Y(_07883_));
 sky130_fd_sc_hd__o21a_1 _14168_ (.A1(\count_instr[56] ),
    .A2(_07881_),
    .B1(_07883_),
    .X(_00954_));
 sky130_fd_sc_hd__and3_1 _14169_ (.A(\count_instr[57] ),
    .B(\count_instr[56] ),
    .C(_07881_),
    .X(_07884_));
 sky130_fd_sc_hd__a21o_1 _14170_ (.A1(\count_instr[56] ),
    .A2(_07881_),
    .B1(\count_instr[57] ),
    .X(_07885_));
 sky130_fd_sc_hd__and3b_1 _14171_ (.A_N(_07884_),
    .B(_07815_),
    .C(_07885_),
    .X(_07886_));
 sky130_fd_sc_hd__clkbuf_1 _14172_ (.A(_07886_),
    .X(_00955_));
 sky130_fd_sc_hd__and4_2 _14173_ (.A(\count_instr[58] ),
    .B(\count_instr[57] ),
    .C(\count_instr[56] ),
    .D(_07881_),
    .X(_07887_));
 sky130_fd_sc_hd__o21ai_1 _14174_ (.A1(\count_instr[58] ),
    .A2(_07884_),
    .B1(_07877_),
    .Y(_07888_));
 sky130_fd_sc_hd__nor2_1 _14175_ (.A(_07887_),
    .B(_07888_),
    .Y(_00956_));
 sky130_fd_sc_hd__a21oi_1 _14176_ (.A1(\count_instr[59] ),
    .A2(_07887_),
    .B1(_07826_),
    .Y(_07889_));
 sky130_fd_sc_hd__o21a_1 _14177_ (.A1(\count_instr[59] ),
    .A2(_07887_),
    .B1(_07889_),
    .X(_00957_));
 sky130_fd_sc_hd__and3_1 _14178_ (.A(\count_instr[60] ),
    .B(\count_instr[59] ),
    .C(_07887_),
    .X(_07890_));
 sky130_fd_sc_hd__a21o_1 _14179_ (.A1(\count_instr[59] ),
    .A2(_07887_),
    .B1(\count_instr[60] ),
    .X(_07891_));
 sky130_fd_sc_hd__and3b_1 _14180_ (.A_N(_07890_),
    .B(_07815_),
    .C(_07891_),
    .X(_07892_));
 sky130_fd_sc_hd__clkbuf_1 _14181_ (.A(_07892_),
    .X(_00958_));
 sky130_fd_sc_hd__and4_2 _14182_ (.A(\count_instr[61] ),
    .B(\count_instr[60] ),
    .C(\count_instr[59] ),
    .D(_07887_),
    .X(_07893_));
 sky130_fd_sc_hd__o21ai_1 _14183_ (.A1(\count_instr[61] ),
    .A2(_07890_),
    .B1(_07877_),
    .Y(_07894_));
 sky130_fd_sc_hd__nor2_1 _14184_ (.A(_07893_),
    .B(_07894_),
    .Y(_00959_));
 sky130_fd_sc_hd__a21oi_1 _14185_ (.A1(\count_instr[62] ),
    .A2(_07893_),
    .B1(_07826_),
    .Y(_07895_));
 sky130_fd_sc_hd__o21a_1 _14186_ (.A1(\count_instr[62] ),
    .A2(_07893_),
    .B1(_07895_),
    .X(_00960_));
 sky130_fd_sc_hd__a21oi_1 _14187_ (.A1(\count_instr[62] ),
    .A2(_07893_),
    .B1(\count_instr[63] ),
    .Y(_07896_));
 sky130_fd_sc_hd__a31o_1 _14188_ (.A1(\count_instr[63] ),
    .A2(\count_instr[62] ),
    .A3(_07893_),
    .B1(_03240_),
    .X(_07897_));
 sky130_fd_sc_hd__nor2_1 _14189_ (.A(_07896_),
    .B(_07897_),
    .Y(_00961_));
 sky130_fd_sc_hd__clkbuf_4 _14190_ (.A(_03293_),
    .X(_07898_));
 sky130_fd_sc_hd__clkbuf_4 _14191_ (.A(_07898_),
    .X(_07899_));
 sky130_fd_sc_hd__or2b_1 _14192_ (.A(latched_branch),
    .B_N(\irq_state[0] ),
    .X(_07900_));
 sky130_fd_sc_hd__clkbuf_4 _14193_ (.A(_07900_),
    .X(_07901_));
 sky130_fd_sc_hd__o211a_1 _14194_ (.A1(_03188_),
    .A2(_06088_),
    .B1(_07901_),
    .C1(_03190_),
    .X(_07902_));
 sky130_fd_sc_hd__nor2_1 _14195_ (.A(_03298_),
    .B(_03196_),
    .Y(_07903_));
 sky130_fd_sc_hd__buf_4 _14196_ (.A(_07903_),
    .X(_07904_));
 sky130_fd_sc_hd__buf_4 _14197_ (.A(_07904_),
    .X(_07905_));
 sky130_fd_sc_hd__clkbuf_4 _14198_ (.A(_07905_),
    .X(_07906_));
 sky130_fd_sc_hd__a22o_1 _14199_ (.A1(_07899_),
    .A2(_07902_),
    .B1(_07906_),
    .B2(\reg_pc[1] ),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _14200_ (.A0(\reg_next_pc[2] ),
    .A1(_06099_),
    .S(_03189_),
    .X(_07907_));
 sky130_fd_sc_hd__nand2_1 _14201_ (.A(_07901_),
    .B(_07907_),
    .Y(_07908_));
 sky130_fd_sc_hd__nor2_1 _14202_ (.A(_06860_),
    .B(_07908_),
    .Y(_07909_));
 sky130_fd_sc_hd__a21o_1 _14203_ (.A1(\reg_pc[2] ),
    .A2(_07906_),
    .B1(_07909_),
    .X(_00963_));
 sky130_fd_sc_hd__or2_1 _14204_ (.A(_03188_),
    .B(_06107_),
    .X(_07910_));
 sky130_fd_sc_hd__o211a_1 _14205_ (.A1(\reg_next_pc[3] ),
    .A2(_03189_),
    .B1(_07900_),
    .C1(_07910_),
    .X(_07911_));
 sky130_fd_sc_hd__clkbuf_4 _14206_ (.A(_03294_),
    .X(_07912_));
 sky130_fd_sc_hd__a22o_1 _14207_ (.A1(\reg_pc[3] ),
    .A2(_07906_),
    .B1(_07911_),
    .B2(_07912_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _14208_ (.A0(\reg_next_pc[4] ),
    .A1(_06117_),
    .S(_03189_),
    .X(_07913_));
 sky130_fd_sc_hd__or2_1 _14209_ (.A(\irq_state[0] ),
    .B(_07913_),
    .X(_07914_));
 sky130_fd_sc_hd__buf_2 _14210_ (.A(_07914_),
    .X(_07915_));
 sky130_fd_sc_hd__a22o_1 _14211_ (.A1(\reg_pc[4] ),
    .A2(_07906_),
    .B1(_07915_),
    .B2(_07912_),
    .X(_00965_));
 sky130_fd_sc_hd__or2_1 _14212_ (.A(_05856_),
    .B(_06128_),
    .X(_07916_));
 sky130_fd_sc_hd__o211a_2 _14213_ (.A1(\reg_next_pc[5] ),
    .A2(_05834_),
    .B1(_07901_),
    .C1(_07916_),
    .X(_07917_));
 sky130_fd_sc_hd__a22o_1 _14214_ (.A1(\reg_pc[5] ),
    .A2(_07906_),
    .B1(_07917_),
    .B2(_07912_),
    .X(_00966_));
 sky130_fd_sc_hd__or2_1 _14215_ (.A(_05856_),
    .B(_06134_),
    .X(_07918_));
 sky130_fd_sc_hd__o211a_2 _14216_ (.A1(\reg_next_pc[6] ),
    .A2(_05834_),
    .B1(_07901_),
    .C1(_07918_),
    .X(_07919_));
 sky130_fd_sc_hd__a22o_1 _14217_ (.A1(\reg_pc[6] ),
    .A2(_07906_),
    .B1(_07919_),
    .B2(_07912_),
    .X(_00967_));
 sky130_fd_sc_hd__or2_1 _14218_ (.A(_05856_),
    .B(_06143_),
    .X(_07920_));
 sky130_fd_sc_hd__o211a_2 _14219_ (.A1(\reg_next_pc[7] ),
    .A2(_05834_),
    .B1(_07901_),
    .C1(_07920_),
    .X(_07921_));
 sky130_fd_sc_hd__a22o_1 _14220_ (.A1(\reg_pc[7] ),
    .A2(_07906_),
    .B1(_07921_),
    .B2(_07912_),
    .X(_00968_));
 sky130_fd_sc_hd__clkbuf_4 _14221_ (.A(_07901_),
    .X(_07922_));
 sky130_fd_sc_hd__or2_1 _14222_ (.A(_05856_),
    .B(_06153_),
    .X(_07923_));
 sky130_fd_sc_hd__o211a_2 _14223_ (.A1(\reg_next_pc[8] ),
    .A2(_05858_),
    .B1(_07922_),
    .C1(_07923_),
    .X(_07924_));
 sky130_fd_sc_hd__a22o_1 _14224_ (.A1(\reg_pc[8] ),
    .A2(_07906_),
    .B1(_07924_),
    .B2(_07912_),
    .X(_00969_));
 sky130_fd_sc_hd__o211a_2 _14225_ (.A1(_05857_),
    .A2(_06159_),
    .B1(_07922_),
    .C1(_05859_),
    .X(_07925_));
 sky130_fd_sc_hd__a22o_1 _14226_ (.A1(\reg_pc[9] ),
    .A2(_07906_),
    .B1(_07925_),
    .B2(_07912_),
    .X(_00970_));
 sky130_fd_sc_hd__clkbuf_4 _14227_ (.A(_07905_),
    .X(_07926_));
 sky130_fd_sc_hd__or2_1 _14228_ (.A(_05856_),
    .B(_06168_),
    .X(_07927_));
 sky130_fd_sc_hd__o211a_2 _14229_ (.A1(\reg_next_pc[10] ),
    .A2(_05858_),
    .B1(_07922_),
    .C1(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__a22o_1 _14230_ (.A1(\reg_pc[10] ),
    .A2(_07926_),
    .B1(_07928_),
    .B2(_07912_),
    .X(_00971_));
 sky130_fd_sc_hd__or2_1 _14231_ (.A(_05856_),
    .B(_06180_),
    .X(_07929_));
 sky130_fd_sc_hd__o211a_2 _14232_ (.A1(\reg_next_pc[11] ),
    .A2(_05834_),
    .B1(_07901_),
    .C1(_07929_),
    .X(_07930_));
 sky130_fd_sc_hd__a22o_1 _14233_ (.A1(\reg_pc[11] ),
    .A2(_07926_),
    .B1(_07930_),
    .B2(_07912_),
    .X(_00972_));
 sky130_fd_sc_hd__or2_1 _14234_ (.A(_05856_),
    .B(_06190_),
    .X(_07931_));
 sky130_fd_sc_hd__o211a_2 _14235_ (.A1(\reg_next_pc[12] ),
    .A2(_05858_),
    .B1(_07901_),
    .C1(_07931_),
    .X(_07932_));
 sky130_fd_sc_hd__a22o_1 _14236_ (.A1(\reg_pc[12] ),
    .A2(_07926_),
    .B1(_07932_),
    .B2(_07912_),
    .X(_00973_));
 sky130_fd_sc_hd__or2_1 _14237_ (.A(_05857_),
    .B(_06198_),
    .X(_07933_));
 sky130_fd_sc_hd__o211a_2 _14238_ (.A1(\reg_next_pc[13] ),
    .A2(_05876_),
    .B1(_07922_),
    .C1(_07933_),
    .X(_07934_));
 sky130_fd_sc_hd__buf_2 _14239_ (.A(_03294_),
    .X(_07935_));
 sky130_fd_sc_hd__a22o_1 _14240_ (.A1(\reg_pc[13] ),
    .A2(_07926_),
    .B1(_07934_),
    .B2(_07935_),
    .X(_00974_));
 sky130_fd_sc_hd__or2_1 _14241_ (.A(_05857_),
    .B(_06205_),
    .X(_07936_));
 sky130_fd_sc_hd__o211a_2 _14242_ (.A1(\reg_next_pc[14] ),
    .A2(_05876_),
    .B1(_07922_),
    .C1(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__a22o_1 _14243_ (.A1(\reg_pc[14] ),
    .A2(_07926_),
    .B1(_07937_),
    .B2(_07935_),
    .X(_00975_));
 sky130_fd_sc_hd__or2_1 _14244_ (.A(_05857_),
    .B(_06213_),
    .X(_07938_));
 sky130_fd_sc_hd__o211a_2 _14245_ (.A1(\reg_next_pc[15] ),
    .A2(_05858_),
    .B1(_07922_),
    .C1(_07938_),
    .X(_07939_));
 sky130_fd_sc_hd__a22o_1 _14246_ (.A1(\reg_pc[15] ),
    .A2(_07926_),
    .B1(_07939_),
    .B2(_07935_),
    .X(_00976_));
 sky130_fd_sc_hd__or2_1 _14247_ (.A(_05856_),
    .B(_06221_),
    .X(_07940_));
 sky130_fd_sc_hd__o211a_2 _14248_ (.A1(\reg_next_pc[16] ),
    .A2(_05858_),
    .B1(_07922_),
    .C1(_07940_),
    .X(_07941_));
 sky130_fd_sc_hd__a22o_1 _14249_ (.A1(\reg_pc[16] ),
    .A2(_07926_),
    .B1(_07941_),
    .B2(_07935_),
    .X(_00977_));
 sky130_fd_sc_hd__clkbuf_4 _14250_ (.A(_07922_),
    .X(_07942_));
 sky130_fd_sc_hd__o211a_2 _14251_ (.A1(_05909_),
    .A2(_06229_),
    .B1(_07942_),
    .C1(_05893_),
    .X(_07943_));
 sky130_fd_sc_hd__a22o_1 _14252_ (.A1(\reg_pc[17] ),
    .A2(_07926_),
    .B1(_07943_),
    .B2(_07935_),
    .X(_00978_));
 sky130_fd_sc_hd__buf_4 _14253_ (.A(_07942_),
    .X(_07944_));
 sky130_fd_sc_hd__o21a_1 _14254_ (.A1(latched_branch),
    .A2(\irq_state[0] ),
    .B1(latched_store),
    .X(_07945_));
 sky130_fd_sc_hd__o22a_2 _14255_ (.A1(_05909_),
    .A2(_06237_),
    .B1(_07945_),
    .B2(\reg_next_pc[18] ),
    .X(_07946_));
 sky130_fd_sc_hd__clkbuf_4 _14256_ (.A(_07904_),
    .X(_07947_));
 sky130_fd_sc_hd__clkbuf_4 _14257_ (.A(_07947_),
    .X(_07948_));
 sky130_fd_sc_hd__a32o_1 _14258_ (.A1(_07899_),
    .A2(_07944_),
    .A3(_07946_),
    .B1(_07948_),
    .B2(\reg_pc[18] ),
    .X(_00979_));
 sky130_fd_sc_hd__or2_1 _14259_ (.A(_05857_),
    .B(_06245_),
    .X(_07949_));
 sky130_fd_sc_hd__o211a_2 _14260_ (.A1(\reg_next_pc[19] ),
    .A2(_05876_),
    .B1(_07922_),
    .C1(_07949_),
    .X(_07950_));
 sky130_fd_sc_hd__a22o_1 _14261_ (.A1(\reg_pc[19] ),
    .A2(_07926_),
    .B1(_07950_),
    .B2(_07935_),
    .X(_00980_));
 sky130_fd_sc_hd__or2_1 _14262_ (.A(_05857_),
    .B(_06254_),
    .X(_07951_));
 sky130_fd_sc_hd__o211a_2 _14263_ (.A1(\reg_next_pc[20] ),
    .A2(_05876_),
    .B1(_07922_),
    .C1(_07951_),
    .X(_07952_));
 sky130_fd_sc_hd__a22o_1 _14264_ (.A1(\reg_pc[20] ),
    .A2(_07926_),
    .B1(_07952_),
    .B2(_07935_),
    .X(_00981_));
 sky130_fd_sc_hd__clkbuf_4 _14265_ (.A(_07905_),
    .X(_07953_));
 sky130_fd_sc_hd__o211a_2 _14266_ (.A1(_05909_),
    .A2(_06263_),
    .B1(_07942_),
    .C1(_05910_),
    .X(_07954_));
 sky130_fd_sc_hd__a22o_1 _14267_ (.A1(\reg_pc[21] ),
    .A2(_07953_),
    .B1(_07954_),
    .B2(_07935_),
    .X(_00982_));
 sky130_fd_sc_hd__or2_1 _14268_ (.A(_05909_),
    .B(_06271_),
    .X(_07955_));
 sky130_fd_sc_hd__o211a_2 _14269_ (.A1(\reg_next_pc[22] ),
    .A2(_05898_),
    .B1(_07942_),
    .C1(_07955_),
    .X(_07956_));
 sky130_fd_sc_hd__a22o_1 _14270_ (.A1(\reg_pc[22] ),
    .A2(_07953_),
    .B1(_07956_),
    .B2(_07935_),
    .X(_00983_));
 sky130_fd_sc_hd__or2_1 _14271_ (.A(_05857_),
    .B(_06278_),
    .X(_07957_));
 sky130_fd_sc_hd__o211a_2 _14272_ (.A1(\reg_next_pc[23] ),
    .A2(_05898_),
    .B1(_07942_),
    .C1(_07957_),
    .X(_07958_));
 sky130_fd_sc_hd__a22o_1 _14273_ (.A1(\reg_pc[23] ),
    .A2(_07953_),
    .B1(_07958_),
    .B2(_07935_),
    .X(_00984_));
 sky130_fd_sc_hd__o211a_2 _14274_ (.A1(_05909_),
    .A2(_06286_),
    .B1(_07942_),
    .C1(_05922_),
    .X(_07959_));
 sky130_fd_sc_hd__buf_4 _14275_ (.A(_03294_),
    .X(_07960_));
 sky130_fd_sc_hd__a22o_1 _14276_ (.A1(\reg_pc[24] ),
    .A2(_07953_),
    .B1(_07959_),
    .B2(_07960_),
    .X(_00985_));
 sky130_fd_sc_hd__o22a_1 _14277_ (.A1(_05909_),
    .A2(_06294_),
    .B1(_07945_),
    .B2(\reg_next_pc[25] ),
    .X(_07961_));
 sky130_fd_sc_hd__and3_1 _14278_ (.A(_03293_),
    .B(_07944_),
    .C(_07961_),
    .X(_07962_));
 sky130_fd_sc_hd__a21o_1 _14279_ (.A1(\reg_pc[25] ),
    .A2(_07906_),
    .B1(_07962_),
    .X(_00986_));
 sky130_fd_sc_hd__or2_1 _14280_ (.A(_05909_),
    .B(_06301_),
    .X(_07963_));
 sky130_fd_sc_hd__o211a_2 _14281_ (.A1(\reg_next_pc[26] ),
    .A2(_05928_),
    .B1(_07942_),
    .C1(_07963_),
    .X(_07964_));
 sky130_fd_sc_hd__a22o_1 _14282_ (.A1(\reg_pc[26] ),
    .A2(_07953_),
    .B1(_07964_),
    .B2(_07960_),
    .X(_00987_));
 sky130_fd_sc_hd__or2_1 _14283_ (.A(_05941_),
    .B(_06309_),
    .X(_07965_));
 sky130_fd_sc_hd__o211a_2 _14284_ (.A1(\reg_next_pc[27] ),
    .A2(_05928_),
    .B1(_07944_),
    .C1(_07965_),
    .X(_07966_));
 sky130_fd_sc_hd__a22o_1 _14285_ (.A1(\reg_pc[27] ),
    .A2(_07953_),
    .B1(_07966_),
    .B2(_07960_),
    .X(_00988_));
 sky130_fd_sc_hd__o211a_2 _14286_ (.A1(_05941_),
    .A2(_06317_),
    .B1(_07944_),
    .C1(_05942_),
    .X(_07967_));
 sky130_fd_sc_hd__a22o_1 _14287_ (.A1(\reg_pc[28] ),
    .A2(_07953_),
    .B1(_07967_),
    .B2(_07960_),
    .X(_00989_));
 sky130_fd_sc_hd__o211a_2 _14288_ (.A1(_05941_),
    .A2(_06325_),
    .B1(_07944_),
    .C1(_05947_),
    .X(_07968_));
 sky130_fd_sc_hd__a22o_1 _14289_ (.A1(\reg_pc[29] ),
    .A2(_07953_),
    .B1(_07968_),
    .B2(_07960_),
    .X(_00990_));
 sky130_fd_sc_hd__o211a_2 _14290_ (.A1(_05941_),
    .A2(_06333_),
    .B1(_07944_),
    .C1(_05951_),
    .X(_07969_));
 sky130_fd_sc_hd__a22o_1 _14291_ (.A1(\reg_pc[30] ),
    .A2(_07953_),
    .B1(_07969_),
    .B2(_07960_),
    .X(_00991_));
 sky130_fd_sc_hd__or2_1 _14292_ (.A(_05941_),
    .B(_06340_),
    .X(_07970_));
 sky130_fd_sc_hd__o211a_2 _14293_ (.A1(\reg_next_pc[31] ),
    .A2(_05928_),
    .B1(_07944_),
    .C1(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__a22o_1 _14294_ (.A1(\reg_pc[31] ),
    .A2(_07953_),
    .B1(_07971_),
    .B2(_07960_),
    .X(_00992_));
 sky130_fd_sc_hd__and2_2 _14295_ (.A(_06863_),
    .B(_03368_),
    .X(_07972_));
 sky130_fd_sc_hd__or4_1 _14296_ (.A(\irq_pending[20] ),
    .B(\irq_pending[21] ),
    .C(\irq_pending[22] ),
    .D(\irq_pending[23] ),
    .X(_07973_));
 sky130_fd_sc_hd__or4_1 _14297_ (.A(\irq_pending[16] ),
    .B(\irq_pending[17] ),
    .C(\irq_pending[18] ),
    .D(\irq_pending[19] ),
    .X(_07974_));
 sky130_fd_sc_hd__or4_1 _14298_ (.A(\irq_pending[28] ),
    .B(\irq_pending[29] ),
    .C(\irq_pending[30] ),
    .D(\irq_pending[31] ),
    .X(_07975_));
 sky130_fd_sc_hd__or4_1 _14299_ (.A(\irq_pending[24] ),
    .B(\irq_pending[25] ),
    .C(\irq_pending[26] ),
    .D(\irq_pending[27] ),
    .X(_07976_));
 sky130_fd_sc_hd__or4_1 _14300_ (.A(_07973_),
    .B(_07974_),
    .C(_07975_),
    .D(_07976_),
    .X(_07977_));
 sky130_fd_sc_hd__or4_1 _14301_ (.A(\irq_pending[8] ),
    .B(\irq_pending[9] ),
    .C(\irq_pending[10] ),
    .D(\irq_pending[11] ),
    .X(_07978_));
 sky130_fd_sc_hd__or4_1 _14302_ (.A(\irq_pending[12] ),
    .B(\irq_pending[13] ),
    .C(\irq_pending[14] ),
    .D(\irq_pending[15] ),
    .X(_07979_));
 sky130_fd_sc_hd__or4_1 _14303_ (.A(\irq_pending[4] ),
    .B(\irq_pending[5] ),
    .C(\irq_pending[6] ),
    .D(\irq_pending[7] ),
    .X(_07980_));
 sky130_fd_sc_hd__or4_1 _14304_ (.A(\irq_pending[0] ),
    .B(\irq_pending[1] ),
    .C(\irq_pending[2] ),
    .D(\irq_pending[3] ),
    .X(_07981_));
 sky130_fd_sc_hd__or3_1 _14305_ (.A(_07979_),
    .B(_07980_),
    .C(_07981_),
    .X(_07982_));
 sky130_fd_sc_hd__or3_2 _14306_ (.A(_07977_),
    .B(_07978_),
    .C(_07982_),
    .X(_07983_));
 sky130_fd_sc_hd__and2_2 _14307_ (.A(_03319_),
    .B(_07983_),
    .X(_07984_));
 sky130_fd_sc_hd__or2_1 _14308_ (.A(_03379_),
    .B(_07984_),
    .X(_07985_));
 sky130_fd_sc_hd__clkbuf_4 _14309_ (.A(_07985_),
    .X(_07986_));
 sky130_fd_sc_hd__and2_1 _14310_ (.A(_03364_),
    .B(_07986_),
    .X(_07987_));
 sky130_fd_sc_hd__buf_2 _14311_ (.A(_07987_),
    .X(_07988_));
 sky130_fd_sc_hd__o211ai_2 _14312_ (.A1(_05856_),
    .A2(_06088_),
    .B1(_07901_),
    .C1(_03190_),
    .Y(_07989_));
 sky130_fd_sc_hd__a211o_1 _14313_ (.A1(compressed_instr),
    .A2(_07988_),
    .B1(_07989_),
    .C1(_06860_),
    .X(_07990_));
 sky130_fd_sc_hd__a21oi_1 _14314_ (.A1(\decoded_imm_j[1] ),
    .A2(_07972_),
    .B1(_07990_),
    .Y(_07991_));
 sky130_fd_sc_hd__o21ai_4 _14315_ (.A1(decoder_trigger),
    .A2(_03319_),
    .B1(_03364_),
    .Y(_07992_));
 sky130_fd_sc_hd__or2_1 _14316_ (.A(_03369_),
    .B(_07983_),
    .X(_07993_));
 sky130_fd_sc_hd__inv_2 _14317_ (.A(_07993_),
    .Y(_07994_));
 sky130_fd_sc_hd__or2_2 _14318_ (.A(_07992_),
    .B(_07994_),
    .X(_07995_));
 sky130_fd_sc_hd__nor2_1 _14319_ (.A(_06860_),
    .B(_07995_),
    .Y(_07996_));
 sky130_fd_sc_hd__clkbuf_4 _14320_ (.A(_07996_),
    .X(_07997_));
 sky130_fd_sc_hd__nor2_4 _14321_ (.A(_03366_),
    .B(_03319_),
    .Y(_07998_));
 sky130_fd_sc_hd__mux2_1 _14322_ (.A0(compressed_instr),
    .A1(\decoded_imm_j[1] ),
    .S(_07998_),
    .X(_07999_));
 sky130_fd_sc_hd__a32o_1 _14323_ (.A1(_07989_),
    .A2(_07997_),
    .A3(_07999_),
    .B1(_07904_),
    .B2(\reg_next_pc[1] ),
    .X(_08000_));
 sky130_fd_sc_hd__or2_1 _14324_ (.A(_07991_),
    .B(_08000_),
    .X(_08001_));
 sky130_fd_sc_hd__clkbuf_1 _14325_ (.A(_08001_),
    .X(_00993_));
 sky130_fd_sc_hd__or2_1 _14326_ (.A(_07909_),
    .B(_07997_),
    .X(_08002_));
 sky130_fd_sc_hd__and2_1 _14327_ (.A(compressed_instr),
    .B(_07989_),
    .X(_08003_));
 sky130_fd_sc_hd__nor2_1 _14328_ (.A(_07908_),
    .B(_08003_),
    .Y(_08004_));
 sky130_fd_sc_hd__and2_1 _14329_ (.A(_07908_),
    .B(_08003_),
    .X(_08005_));
 sky130_fd_sc_hd__o21ai_1 _14330_ (.A1(_08004_),
    .A2(_08005_),
    .B1(_07988_),
    .Y(_08006_));
 sky130_fd_sc_hd__and3_1 _14331_ (.A(\decoded_imm_j[2] ),
    .B(_07900_),
    .C(_07907_),
    .X(_08007_));
 sky130_fd_sc_hd__a21oi_1 _14332_ (.A1(_07901_),
    .A2(_07907_),
    .B1(\decoded_imm_j[2] ),
    .Y(_08008_));
 sky130_fd_sc_hd__nor2_1 _14333_ (.A(_08007_),
    .B(_08008_),
    .Y(_08009_));
 sky130_fd_sc_hd__and3_1 _14334_ (.A(\decoded_imm_j[1] ),
    .B(_07902_),
    .C(_08009_),
    .X(_08010_));
 sky130_fd_sc_hd__a21oi_1 _14335_ (.A1(\decoded_imm_j[1] ),
    .A2(_07902_),
    .B1(_08009_),
    .Y(_08011_));
 sky130_fd_sc_hd__clkbuf_4 _14336_ (.A(_07972_),
    .X(_08012_));
 sky130_fd_sc_hd__o21ai_1 _14337_ (.A1(_08010_),
    .A2(_08011_),
    .B1(_08012_),
    .Y(_08013_));
 sky130_fd_sc_hd__a32o_1 _14338_ (.A1(_08002_),
    .A2(_08006_),
    .A3(_08013_),
    .B1(_07905_),
    .B2(\reg_next_pc[2] ),
    .X(_00994_));
 sky130_fd_sc_hd__or2_1 _14339_ (.A(_07998_),
    .B(_08004_),
    .X(_08014_));
 sky130_fd_sc_hd__a22o_1 _14340_ (.A1(_03294_),
    .A2(_07911_),
    .B1(_07997_),
    .B2(_08014_),
    .X(_08015_));
 sky130_fd_sc_hd__and2_1 _14341_ (.A(_07911_),
    .B(_08004_),
    .X(_08016_));
 sky130_fd_sc_hd__and2_1 _14342_ (.A(\decoded_imm_j[3] ),
    .B(_07911_),
    .X(_08017_));
 sky130_fd_sc_hd__nor2_1 _14343_ (.A(\decoded_imm_j[3] ),
    .B(_07911_),
    .Y(_08018_));
 sky130_fd_sc_hd__or2_1 _14344_ (.A(_08017_),
    .B(_08018_),
    .X(_08019_));
 sky130_fd_sc_hd__nor2_1 _14345_ (.A(_08007_),
    .B(_08010_),
    .Y(_08020_));
 sky130_fd_sc_hd__xnor2_1 _14346_ (.A(_08019_),
    .B(_08020_),
    .Y(_08021_));
 sky130_fd_sc_hd__a22oi_1 _14347_ (.A1(_07988_),
    .A2(_08016_),
    .B1(_08021_),
    .B2(_08012_),
    .Y(_08022_));
 sky130_fd_sc_hd__a22o_1 _14348_ (.A1(\reg_next_pc[3] ),
    .A2(_07948_),
    .B1(_08015_),
    .B2(_08022_),
    .X(_00995_));
 sky130_fd_sc_hd__o21ba_1 _14349_ (.A1(_08007_),
    .A2(_08010_),
    .B1_N(_08019_),
    .X(_08023_));
 sky130_fd_sc_hd__nand2_1 _14350_ (.A(\decoded_imm_j[4] ),
    .B(_07915_),
    .Y(_08024_));
 sky130_fd_sc_hd__or2_1 _14351_ (.A(\decoded_imm_j[4] ),
    .B(_07915_),
    .X(_08025_));
 sky130_fd_sc_hd__and2_1 _14352_ (.A(_08024_),
    .B(_08025_),
    .X(_08026_));
 sky130_fd_sc_hd__or3_1 _14353_ (.A(_08017_),
    .B(_08023_),
    .C(_08026_),
    .X(_08027_));
 sky130_fd_sc_hd__o21ai_2 _14354_ (.A1(_08017_),
    .A2(_08023_),
    .B1(_08026_),
    .Y(_08028_));
 sky130_fd_sc_hd__nand2_1 _14355_ (.A(_07915_),
    .B(_08016_),
    .Y(_08029_));
 sky130_fd_sc_hd__or2_1 _14356_ (.A(_07915_),
    .B(_08016_),
    .X(_08030_));
 sky130_fd_sc_hd__a32o_1 _14357_ (.A1(_07986_),
    .A2(_08029_),
    .A3(_08030_),
    .B1(_07994_),
    .B2(_07915_),
    .X(_08031_));
 sky130_fd_sc_hd__a31o_1 _14358_ (.A1(_03368_),
    .A2(_08027_),
    .A3(_08028_),
    .B1(_08031_),
    .X(_08032_));
 sky130_fd_sc_hd__clkbuf_4 _14359_ (.A(_03378_),
    .X(_08033_));
 sky130_fd_sc_hd__a22o_1 _14360_ (.A1(\reg_next_pc[4] ),
    .A2(_07947_),
    .B1(_08032_),
    .B2(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__a31o_1 _14361_ (.A1(_07960_),
    .A2(_07915_),
    .A3(_07992_),
    .B1(_08034_),
    .X(_00996_));
 sky130_fd_sc_hd__nor2_4 _14362_ (.A(_03379_),
    .B(_07984_),
    .Y(_08035_));
 sky130_fd_sc_hd__and3_1 _14363_ (.A(_07915_),
    .B(_07917_),
    .C(_08016_),
    .X(_08036_));
 sky130_fd_sc_hd__a21oi_1 _14364_ (.A1(_07915_),
    .A2(_08016_),
    .B1(_07917_),
    .Y(_08037_));
 sky130_fd_sc_hd__nand2_1 _14365_ (.A(\decoded_imm_j[5] ),
    .B(_07917_),
    .Y(_08038_));
 sky130_fd_sc_hd__or2_1 _14366_ (.A(\decoded_imm_j[5] ),
    .B(_07917_),
    .X(_08039_));
 sky130_fd_sc_hd__nand2_1 _14367_ (.A(_08038_),
    .B(_08039_),
    .Y(_08040_));
 sky130_fd_sc_hd__a21o_1 _14368_ (.A1(_08024_),
    .A2(_08028_),
    .B1(_08040_),
    .X(_08041_));
 sky130_fd_sc_hd__nand2_1 _14369_ (.A(_03368_),
    .B(_08041_),
    .Y(_08042_));
 sky130_fd_sc_hd__a31o_1 _14370_ (.A1(_08024_),
    .A2(_08028_),
    .A3(_08040_),
    .B1(_08042_),
    .X(_08043_));
 sky130_fd_sc_hd__o31ai_1 _14371_ (.A1(_08035_),
    .A2(_08036_),
    .A3(_08037_),
    .B1(_08043_),
    .Y(_08044_));
 sky130_fd_sc_hd__a21o_1 _14372_ (.A1(_07917_),
    .A2(_07994_),
    .B1(_08044_),
    .X(_08045_));
 sky130_fd_sc_hd__a22o_1 _14373_ (.A1(\reg_next_pc[5] ),
    .A2(_07947_),
    .B1(_08045_),
    .B2(_08033_),
    .X(_08046_));
 sky130_fd_sc_hd__a31o_1 _14374_ (.A1(_07899_),
    .A2(_07917_),
    .A3(_07992_),
    .B1(_08046_),
    .X(_00997_));
 sky130_fd_sc_hd__a21o_1 _14375_ (.A1(_06863_),
    .A2(_08036_),
    .B1(_07919_),
    .X(_08047_));
 sky130_fd_sc_hd__and2_1 _14376_ (.A(_07919_),
    .B(_08036_),
    .X(_08048_));
 sky130_fd_sc_hd__inv_2 _14377_ (.A(_08048_),
    .Y(_08049_));
 sky130_fd_sc_hd__clkbuf_4 _14378_ (.A(_07995_),
    .X(_08050_));
 sky130_fd_sc_hd__a32o_1 _14379_ (.A1(_07986_),
    .A2(_08047_),
    .A3(_08049_),
    .B1(_08050_),
    .B2(_07919_),
    .X(_08051_));
 sky130_fd_sc_hd__nand2_1 _14380_ (.A(\decoded_imm_j[6] ),
    .B(_07919_),
    .Y(_08052_));
 sky130_fd_sc_hd__or2_1 _14381_ (.A(\decoded_imm_j[6] ),
    .B(_07919_),
    .X(_08053_));
 sky130_fd_sc_hd__nand2_1 _14382_ (.A(_08052_),
    .B(_08053_),
    .Y(_08054_));
 sky130_fd_sc_hd__nand2_2 _14383_ (.A(_03368_),
    .B(_03378_),
    .Y(_08055_));
 sky130_fd_sc_hd__a31o_1 _14384_ (.A1(_08038_),
    .A2(_08041_),
    .A3(_08054_),
    .B1(_08055_),
    .X(_08056_));
 sky130_fd_sc_hd__a211o_1 _14385_ (.A1(_08024_),
    .A2(_08028_),
    .B1(_08040_),
    .C1(_08054_),
    .X(_08057_));
 sky130_fd_sc_hd__or2_1 _14386_ (.A(_08038_),
    .B(_08054_),
    .X(_08058_));
 sky130_fd_sc_hd__and3b_1 _14387_ (.A_N(_08056_),
    .B(_08057_),
    .C(_08058_),
    .X(_08059_));
 sky130_fd_sc_hd__a221o_1 _14388_ (.A1(\reg_next_pc[6] ),
    .A2(_07905_),
    .B1(_08051_),
    .B2(_07899_),
    .C1(_08059_),
    .X(_00998_));
 sky130_fd_sc_hd__nand2_1 _14389_ (.A(\decoded_imm_j[7] ),
    .B(_07921_),
    .Y(_08060_));
 sky130_fd_sc_hd__or2_1 _14390_ (.A(\decoded_imm_j[7] ),
    .B(_07921_),
    .X(_08061_));
 sky130_fd_sc_hd__nand2_1 _14391_ (.A(_08060_),
    .B(_08061_),
    .Y(_08062_));
 sky130_fd_sc_hd__and4_1 _14392_ (.A(_08052_),
    .B(_08058_),
    .C(_08057_),
    .D(_08062_),
    .X(_08063_));
 sky130_fd_sc_hd__a31o_1 _14393_ (.A1(_08052_),
    .A2(_08058_),
    .A3(_08057_),
    .B1(_08062_),
    .X(_08064_));
 sky130_fd_sc_hd__nand2_1 _14394_ (.A(_03368_),
    .B(_08064_),
    .Y(_08065_));
 sky130_fd_sc_hd__xnor2_1 _14395_ (.A(_07921_),
    .B(_08048_),
    .Y(_08066_));
 sky130_fd_sc_hd__o22a_1 _14396_ (.A1(_08063_),
    .A2(_08065_),
    .B1(_08066_),
    .B2(_08035_),
    .X(_08067_));
 sky130_fd_sc_hd__a21bo_1 _14397_ (.A1(_07921_),
    .A2(_07994_),
    .B1_N(_08067_),
    .X(_08068_));
 sky130_fd_sc_hd__a22o_1 _14398_ (.A1(\reg_next_pc[7] ),
    .A2(_07947_),
    .B1(_08068_),
    .B2(_08033_),
    .X(_08069_));
 sky130_fd_sc_hd__a31o_1 _14399_ (.A1(_07899_),
    .A2(_07921_),
    .A3(_07992_),
    .B1(_08069_),
    .X(_00999_));
 sky130_fd_sc_hd__and2_1 _14400_ (.A(_03368_),
    .B(_03378_),
    .X(_08070_));
 sky130_fd_sc_hd__buf_2 _14401_ (.A(_08070_),
    .X(_08071_));
 sky130_fd_sc_hd__and2_1 _14402_ (.A(\decoded_imm_j[8] ),
    .B(_07924_),
    .X(_08072_));
 sky130_fd_sc_hd__nor2_1 _14403_ (.A(\decoded_imm_j[8] ),
    .B(_07924_),
    .Y(_08073_));
 sky130_fd_sc_hd__a211o_1 _14404_ (.A1(_08060_),
    .A2(_08064_),
    .B1(_08072_),
    .C1(_08073_),
    .X(_08074_));
 sky130_fd_sc_hd__o211ai_1 _14405_ (.A1(_08072_),
    .A2(_08073_),
    .B1(_08060_),
    .C1(_08064_),
    .Y(_08075_));
 sky130_fd_sc_hd__and3_1 _14406_ (.A(_07921_),
    .B(_07924_),
    .C(_08048_),
    .X(_08076_));
 sky130_fd_sc_hd__a2bb2o_1 _14407_ (.A1_N(_08035_),
    .A2_N(_08076_),
    .B1(_07995_),
    .B2(_07924_),
    .X(_08077_));
 sky130_fd_sc_hd__a32o_1 _14408_ (.A1(_03378_),
    .A2(_07921_),
    .A3(_08048_),
    .B1(_07924_),
    .B2(_03293_),
    .X(_08078_));
 sky130_fd_sc_hd__a22o_1 _14409_ (.A1(\reg_next_pc[8] ),
    .A2(_07947_),
    .B1(_08077_),
    .B2(_08078_),
    .X(_08079_));
 sky130_fd_sc_hd__a31o_1 _14410_ (.A1(_08071_),
    .A2(_08074_),
    .A3(_08075_),
    .B1(_08079_),
    .X(_01000_));
 sky130_fd_sc_hd__or2_1 _14411_ (.A(_07998_),
    .B(_08076_),
    .X(_08080_));
 sky130_fd_sc_hd__a22o_1 _14412_ (.A1(_03294_),
    .A2(_07925_),
    .B1(_07997_),
    .B2(_08080_),
    .X(_08081_));
 sky130_fd_sc_hd__nand2_1 _14413_ (.A(\decoded_imm_j[9] ),
    .B(_07925_),
    .Y(_08082_));
 sky130_fd_sc_hd__or2_1 _14414_ (.A(\decoded_imm_j[9] ),
    .B(_07925_),
    .X(_08083_));
 sky130_fd_sc_hd__nand2_1 _14415_ (.A(_08082_),
    .B(_08083_),
    .Y(_08084_));
 sky130_fd_sc_hd__nand2_1 _14416_ (.A(\decoded_imm_j[8] ),
    .B(_07924_),
    .Y(_08085_));
 sky130_fd_sc_hd__a31o_1 _14417_ (.A1(_08060_),
    .A2(_08064_),
    .A3(_08085_),
    .B1(_08073_),
    .X(_08086_));
 sky130_fd_sc_hd__or2_1 _14418_ (.A(_08084_),
    .B(_08086_),
    .X(_08087_));
 sky130_fd_sc_hd__nand2_1 _14419_ (.A(_08084_),
    .B(_08086_),
    .Y(_08088_));
 sky130_fd_sc_hd__nand2_1 _14420_ (.A(_08087_),
    .B(_08088_),
    .Y(_08089_));
 sky130_fd_sc_hd__and3_1 _14421_ (.A(_07925_),
    .B(_07988_),
    .C(_08076_),
    .X(_08090_));
 sky130_fd_sc_hd__a21oi_1 _14422_ (.A1(_08012_),
    .A2(_08089_),
    .B1(_08090_),
    .Y(_08091_));
 sky130_fd_sc_hd__a22o_1 _14423_ (.A1(\reg_next_pc[9] ),
    .A2(_07948_),
    .B1(_08081_),
    .B2(_08091_),
    .X(_01001_));
 sky130_fd_sc_hd__and3_1 _14424_ (.A(_07925_),
    .B(_07928_),
    .C(_08076_),
    .X(_08092_));
 sky130_fd_sc_hd__a21oi_1 _14425_ (.A1(_07925_),
    .A2(_08076_),
    .B1(_07928_),
    .Y(_08093_));
 sky130_fd_sc_hd__xnor2_2 _14426_ (.A(\decoded_imm_j[10] ),
    .B(_07928_),
    .Y(_08094_));
 sky130_fd_sc_hd__nor2_1 _14427_ (.A(_08087_),
    .B(_08094_),
    .Y(_08095_));
 sky130_fd_sc_hd__nor2_1 _14428_ (.A(_08082_),
    .B(_08094_),
    .Y(_08096_));
 sky130_fd_sc_hd__nand2_2 _14429_ (.A(instr_jal),
    .B(_07754_),
    .Y(_08097_));
 sky130_fd_sc_hd__a311o_1 _14430_ (.A1(_08082_),
    .A2(_08087_),
    .A3(_08094_),
    .B1(_08096_),
    .C1(_08097_),
    .X(_08098_));
 sky130_fd_sc_hd__o32a_1 _14431_ (.A1(_08035_),
    .A2(_08092_),
    .A3(_08093_),
    .B1(_08095_),
    .B2(_08098_),
    .X(_08099_));
 sky130_fd_sc_hd__inv_2 _14432_ (.A(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__a22o_1 _14433_ (.A1(\reg_next_pc[10] ),
    .A2(_07947_),
    .B1(_08100_),
    .B2(_08033_),
    .X(_08101_));
 sky130_fd_sc_hd__a31o_1 _14434_ (.A1(_07899_),
    .A2(_07928_),
    .A3(_08050_),
    .B1(_08101_),
    .X(_01002_));
 sky130_fd_sc_hd__and2_1 _14435_ (.A(_07930_),
    .B(_08092_),
    .X(_08102_));
 sky130_fd_sc_hd__o21ai_1 _14436_ (.A1(_07930_),
    .A2(_08092_),
    .B1(_07986_),
    .Y(_08103_));
 sky130_fd_sc_hd__nand2_1 _14437_ (.A(\decoded_imm_j[11] ),
    .B(_07930_),
    .Y(_08104_));
 sky130_fd_sc_hd__or2_1 _14438_ (.A(\decoded_imm_j[11] ),
    .B(_07930_),
    .X(_08105_));
 sky130_fd_sc_hd__nand2_1 _14439_ (.A(_08104_),
    .B(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__a21oi_1 _14440_ (.A1(\decoded_imm_j[10] ),
    .A2(_07928_),
    .B1(_08096_),
    .Y(_08107_));
 sky130_fd_sc_hd__o21a_1 _14441_ (.A1(_08087_),
    .A2(_08094_),
    .B1(_08107_),
    .X(_08108_));
 sky130_fd_sc_hd__o21a_1 _14442_ (.A1(_08106_),
    .A2(_08108_),
    .B1(_03368_),
    .X(_08109_));
 sky130_fd_sc_hd__nand2_1 _14443_ (.A(_08106_),
    .B(_08108_),
    .Y(_08110_));
 sky130_fd_sc_hd__a2bb2o_1 _14444_ (.A1_N(_08102_),
    .A2_N(_08103_),
    .B1(_08109_),
    .B2(_08110_),
    .X(_08111_));
 sky130_fd_sc_hd__a22o_1 _14445_ (.A1(\reg_next_pc[11] ),
    .A2(_07947_),
    .B1(_08111_),
    .B2(_08033_),
    .X(_08112_));
 sky130_fd_sc_hd__a31o_1 _14446_ (.A1(_07899_),
    .A2(_07930_),
    .A3(_08050_),
    .B1(_08112_),
    .X(_01003_));
 sky130_fd_sc_hd__and2_1 _14447_ (.A(\decoded_imm_j[12] ),
    .B(_07932_),
    .X(_08113_));
 sky130_fd_sc_hd__nor2_1 _14448_ (.A(\decoded_imm_j[12] ),
    .B(_07932_),
    .Y(_08114_));
 sky130_fd_sc_hd__nor2_1 _14449_ (.A(_08113_),
    .B(_08114_),
    .Y(_08115_));
 sky130_fd_sc_hd__o21a_1 _14450_ (.A1(_08106_),
    .A2(_08108_),
    .B1(_08104_),
    .X(_08116_));
 sky130_fd_sc_hd__xnor2_1 _14451_ (.A(_08115_),
    .B(_08116_),
    .Y(_08117_));
 sky130_fd_sc_hd__a32o_1 _14452_ (.A1(_07898_),
    .A2(_07932_),
    .A3(_08050_),
    .B1(_07947_),
    .B2(\reg_next_pc[12] ),
    .X(_08118_));
 sky130_fd_sc_hd__and3_2 _14453_ (.A(_07930_),
    .B(_07932_),
    .C(_08092_),
    .X(_08119_));
 sky130_fd_sc_hd__nand2_2 _14454_ (.A(_03364_),
    .B(_07986_),
    .Y(_08120_));
 sky130_fd_sc_hd__nor2_2 _14455_ (.A(_06860_),
    .B(_08120_),
    .Y(_08121_));
 sky130_fd_sc_hd__o21ai_1 _14456_ (.A1(_07932_),
    .A2(_08102_),
    .B1(_08121_),
    .Y(_08122_));
 sky130_fd_sc_hd__nor2_1 _14457_ (.A(_08119_),
    .B(_08122_),
    .Y(_08123_));
 sky130_fd_sc_hd__a211o_1 _14458_ (.A1(_08071_),
    .A2(_08117_),
    .B1(_08118_),
    .C1(_08123_),
    .X(_01004_));
 sky130_fd_sc_hd__or3_1 _14459_ (.A(_08106_),
    .B(_08113_),
    .C(_08114_),
    .X(_08124_));
 sky130_fd_sc_hd__nand2_1 _14460_ (.A(\decoded_imm_j[12] ),
    .B(_07932_),
    .Y(_08125_));
 sky130_fd_sc_hd__o221a_1 _14461_ (.A1(_08104_),
    .A2(_08114_),
    .B1(_08124_),
    .B2(_08107_),
    .C1(_08125_),
    .X(_08126_));
 sky130_fd_sc_hd__or4_1 _14462_ (.A(_08084_),
    .B(_08086_),
    .C(_08094_),
    .D(_08124_),
    .X(_08127_));
 sky130_fd_sc_hd__and2_1 _14463_ (.A(\decoded_imm_j[13] ),
    .B(_07934_),
    .X(_08128_));
 sky130_fd_sc_hd__nor2_1 _14464_ (.A(\decoded_imm_j[13] ),
    .B(_07934_),
    .Y(_08129_));
 sky130_fd_sc_hd__or2_1 _14465_ (.A(_08128_),
    .B(_08129_),
    .X(_08130_));
 sky130_fd_sc_hd__a21oi_2 _14466_ (.A1(_08126_),
    .A2(_08127_),
    .B1(_08130_),
    .Y(_08131_));
 sky130_fd_sc_hd__and3_1 _14467_ (.A(_08130_),
    .B(_08126_),
    .C(_08127_),
    .X(_08132_));
 sky130_fd_sc_hd__o21ai_1 _14468_ (.A1(_08131_),
    .A2(_08132_),
    .B1(_08012_),
    .Y(_08133_));
 sky130_fd_sc_hd__o21a_1 _14469_ (.A1(_07998_),
    .A2(_08119_),
    .B1(_07996_),
    .X(_08134_));
 sky130_fd_sc_hd__a21o_1 _14470_ (.A1(_07898_),
    .A2(_07934_),
    .B1(_08134_),
    .X(_08135_));
 sky130_fd_sc_hd__nand2_1 _14471_ (.A(_07934_),
    .B(_08119_),
    .Y(_08136_));
 sky130_fd_sc_hd__nor2_1 _14472_ (.A(_08035_),
    .B(_08136_),
    .Y(_08137_));
 sky130_fd_sc_hd__nand2_1 _14473_ (.A(_06863_),
    .B(_08137_),
    .Y(_08138_));
 sky130_fd_sc_hd__a32o_1 _14474_ (.A1(_08133_),
    .A2(_08135_),
    .A3(_08138_),
    .B1(_07905_),
    .B2(\reg_next_pc[13] ),
    .X(_01005_));
 sky130_fd_sc_hd__and2_1 _14475_ (.A(\decoded_imm_j[14] ),
    .B(_07937_),
    .X(_08139_));
 sky130_fd_sc_hd__nor2_1 _14476_ (.A(\decoded_imm_j[14] ),
    .B(_07937_),
    .Y(_08140_));
 sky130_fd_sc_hd__or2_1 _14477_ (.A(_08139_),
    .B(_08140_),
    .X(_08141_));
 sky130_fd_sc_hd__o21bai_1 _14478_ (.A1(_08128_),
    .A2(_08131_),
    .B1_N(_08141_),
    .Y(_08142_));
 sky130_fd_sc_hd__or3b_1 _14479_ (.A(_08128_),
    .B(_08131_),
    .C_N(_08141_),
    .X(_08143_));
 sky130_fd_sc_hd__a21o_1 _14480_ (.A1(_07986_),
    .A2(_08136_),
    .B1(_07994_),
    .X(_08144_));
 sky130_fd_sc_hd__mux2_1 _14481_ (.A0(_08137_),
    .A1(_08144_),
    .S(_07937_),
    .X(_08145_));
 sky130_fd_sc_hd__a22o_1 _14482_ (.A1(_07937_),
    .A2(_07992_),
    .B1(_08145_),
    .B2(_06863_),
    .X(_08146_));
 sky130_fd_sc_hd__a31o_1 _14483_ (.A1(_08012_),
    .A2(_08142_),
    .A3(_08143_),
    .B1(_08146_),
    .X(_08147_));
 sky130_fd_sc_hd__a22o_1 _14484_ (.A1(\reg_next_pc[14] ),
    .A2(_07948_),
    .B1(_08147_),
    .B2(_07960_),
    .X(_01006_));
 sky130_fd_sc_hd__nand2_1 _14485_ (.A(\decoded_imm_j[15] ),
    .B(_07939_),
    .Y(_08148_));
 sky130_fd_sc_hd__or2_1 _14486_ (.A(\decoded_imm_j[15] ),
    .B(_07939_),
    .X(_08149_));
 sky130_fd_sc_hd__nand2_1 _14487_ (.A(_08148_),
    .B(_08149_),
    .Y(_08150_));
 sky130_fd_sc_hd__nor2_1 _14488_ (.A(_08128_),
    .B(_08139_),
    .Y(_08151_));
 sky130_fd_sc_hd__and2b_1 _14489_ (.A_N(_08131_),
    .B(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__or3_1 _14490_ (.A(_08140_),
    .B(_08150_),
    .C(_08152_),
    .X(_08153_));
 sky130_fd_sc_hd__o21ai_1 _14491_ (.A1(_08140_),
    .A2(_08152_),
    .B1(_08150_),
    .Y(_08154_));
 sky130_fd_sc_hd__a31o_1 _14492_ (.A1(_07934_),
    .A2(_07937_),
    .A3(_08119_),
    .B1(_07939_),
    .X(_08155_));
 sky130_fd_sc_hd__nand4_2 _14493_ (.A(_07934_),
    .B(_07937_),
    .C(_07939_),
    .D(_08119_),
    .Y(_08156_));
 sky130_fd_sc_hd__a32o_1 _14494_ (.A1(_07986_),
    .A2(_08155_),
    .A3(_08156_),
    .B1(_07994_),
    .B2(_07939_),
    .X(_08157_));
 sky130_fd_sc_hd__a31o_1 _14495_ (.A1(_03368_),
    .A2(_08153_),
    .A3(_08154_),
    .B1(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__a22o_1 _14496_ (.A1(\reg_next_pc[15] ),
    .A2(_07947_),
    .B1(_08158_),
    .B2(_08033_),
    .X(_08159_));
 sky130_fd_sc_hd__a31o_1 _14497_ (.A1(_07899_),
    .A2(_07939_),
    .A3(_07992_),
    .B1(_08159_),
    .X(_01007_));
 sky130_fd_sc_hd__inv_2 _14498_ (.A(_07941_),
    .Y(_08160_));
 sky130_fd_sc_hd__nand2_1 _14499_ (.A(_08160_),
    .B(_08156_),
    .Y(_08161_));
 sky130_fd_sc_hd__nor2_1 _14500_ (.A(_08160_),
    .B(_08156_),
    .Y(_08162_));
 sky130_fd_sc_hd__nor2_1 _14501_ (.A(_08120_),
    .B(_08162_),
    .Y(_08163_));
 sky130_fd_sc_hd__and2_1 _14502_ (.A(\decoded_imm_j[16] ),
    .B(_07941_),
    .X(_08164_));
 sky130_fd_sc_hd__nor2_1 _14503_ (.A(\decoded_imm_j[16] ),
    .B(_07941_),
    .Y(_08165_));
 sky130_fd_sc_hd__or2_1 _14504_ (.A(_08164_),
    .B(_08165_),
    .X(_08166_));
 sky130_fd_sc_hd__and2_1 _14505_ (.A(_08148_),
    .B(_08153_),
    .X(_08167_));
 sky130_fd_sc_hd__nand2_1 _14506_ (.A(_08166_),
    .B(_08167_),
    .Y(_08168_));
 sky130_fd_sc_hd__or2_1 _14507_ (.A(_08166_),
    .B(_08167_),
    .X(_08169_));
 sky130_fd_sc_hd__a32o_1 _14508_ (.A1(_07972_),
    .A2(_08168_),
    .A3(_08169_),
    .B1(_08050_),
    .B2(_07941_),
    .X(_08170_));
 sky130_fd_sc_hd__a21o_1 _14509_ (.A1(_08161_),
    .A2(_08163_),
    .B1(_08170_),
    .X(_08171_));
 sky130_fd_sc_hd__a22o_1 _14510_ (.A1(\reg_next_pc[16] ),
    .A2(_07948_),
    .B1(_08171_),
    .B2(_07960_),
    .X(_01008_));
 sky130_fd_sc_hd__or2_1 _14511_ (.A(_08150_),
    .B(_08166_),
    .X(_08172_));
 sky130_fd_sc_hd__or3_1 _14512_ (.A(_08140_),
    .B(_08151_),
    .C(_08172_),
    .X(_08173_));
 sky130_fd_sc_hd__nor2_1 _14513_ (.A(_08141_),
    .B(_08172_),
    .Y(_08174_));
 sky130_fd_sc_hd__a22oi_1 _14514_ (.A1(\decoded_imm_j[16] ),
    .A2(_07941_),
    .B1(_08131_),
    .B2(_08174_),
    .Y(_08175_));
 sky130_fd_sc_hd__o211a_1 _14515_ (.A1(_08148_),
    .A2(_08165_),
    .B1(_08173_),
    .C1(_08175_),
    .X(_08176_));
 sky130_fd_sc_hd__nand2_1 _14516_ (.A(\decoded_imm_j[17] ),
    .B(_07943_),
    .Y(_08177_));
 sky130_fd_sc_hd__or2_1 _14517_ (.A(\decoded_imm_j[17] ),
    .B(_07943_),
    .X(_08178_));
 sky130_fd_sc_hd__nand2_1 _14518_ (.A(_08177_),
    .B(_08178_),
    .Y(_08179_));
 sky130_fd_sc_hd__or2_2 _14519_ (.A(_08176_),
    .B(_08179_),
    .X(_08180_));
 sky130_fd_sc_hd__nand2_1 _14520_ (.A(_08176_),
    .B(_08179_),
    .Y(_08181_));
 sky130_fd_sc_hd__a21bo_1 _14521_ (.A1(_08180_),
    .A2(_08181_),
    .B1_N(_08012_),
    .X(_08182_));
 sky130_fd_sc_hd__or2_1 _14522_ (.A(_07998_),
    .B(_08162_),
    .X(_08183_));
 sky130_fd_sc_hd__a22o_1 _14523_ (.A1(_07898_),
    .A2(_07943_),
    .B1(_07997_),
    .B2(_08183_),
    .X(_08184_));
 sky130_fd_sc_hd__nand2_1 _14524_ (.A(_07943_),
    .B(_08162_),
    .Y(_08185_));
 sky130_fd_sc_hd__or2_1 _14525_ (.A(_08120_),
    .B(_08185_),
    .X(_08186_));
 sky130_fd_sc_hd__a32o_1 _14526_ (.A1(_08182_),
    .A2(_08184_),
    .A3(_08186_),
    .B1(_07905_),
    .B2(\reg_next_pc[17] ),
    .X(_01009_));
 sky130_fd_sc_hd__a21oi_1 _14527_ (.A1(_07942_),
    .A2(_07946_),
    .B1(\decoded_imm_j[18] ),
    .Y(_08187_));
 sky130_fd_sc_hd__nand3_1 _14528_ (.A(\decoded_imm_j[18] ),
    .B(_07942_),
    .C(_07946_),
    .Y(_08188_));
 sky130_fd_sc_hd__or2b_1 _14529_ (.A(_08187_),
    .B_N(_08188_),
    .X(_08189_));
 sky130_fd_sc_hd__a21o_1 _14530_ (.A1(_08177_),
    .A2(_08180_),
    .B1(_08189_),
    .X(_08190_));
 sky130_fd_sc_hd__nand3_1 _14531_ (.A(_08177_),
    .B(_08180_),
    .C(_08189_),
    .Y(_08191_));
 sky130_fd_sc_hd__nor2_1 _14532_ (.A(_07946_),
    .B(_08185_),
    .Y(_08192_));
 sky130_fd_sc_hd__a21o_1 _14533_ (.A1(_07986_),
    .A2(_08185_),
    .B1(_07995_),
    .X(_08193_));
 sky130_fd_sc_hd__and4_1 _14534_ (.A(_03293_),
    .B(_07944_),
    .C(_07946_),
    .D(_08193_),
    .X(_08194_));
 sky130_fd_sc_hd__a221o_1 _14535_ (.A1(\reg_next_pc[18] ),
    .A2(_07904_),
    .B1(_08121_),
    .B2(_08192_),
    .C1(_08194_),
    .X(_08195_));
 sky130_fd_sc_hd__a31o_1 _14536_ (.A1(_08071_),
    .A2(_08190_),
    .A3(_08191_),
    .B1(_08195_),
    .X(_01010_));
 sky130_fd_sc_hd__nand2_1 _14537_ (.A(\decoded_imm_j[19] ),
    .B(_07950_),
    .Y(_08196_));
 sky130_fd_sc_hd__or2_1 _14538_ (.A(\decoded_imm_j[19] ),
    .B(_07950_),
    .X(_08197_));
 sky130_fd_sc_hd__nand2_1 _14539_ (.A(_08196_),
    .B(_08197_),
    .Y(_08198_));
 sky130_fd_sc_hd__and2_1 _14540_ (.A(_08177_),
    .B(_08188_),
    .X(_08199_));
 sky130_fd_sc_hd__a21o_1 _14541_ (.A1(_08180_),
    .A2(_08199_),
    .B1(_08187_),
    .X(_08200_));
 sky130_fd_sc_hd__or2_1 _14542_ (.A(_08198_),
    .B(_08200_),
    .X(_08201_));
 sky130_fd_sc_hd__nand2_1 _14543_ (.A(_08198_),
    .B(_08200_),
    .Y(_08202_));
 sky130_fd_sc_hd__a21bo_1 _14544_ (.A1(_08201_),
    .A2(_08202_),
    .B1_N(_07972_),
    .X(_08203_));
 sky130_fd_sc_hd__a31o_1 _14545_ (.A1(_07943_),
    .A2(_07946_),
    .A3(_08162_),
    .B1(_07998_),
    .X(_08204_));
 sky130_fd_sc_hd__a22o_1 _14546_ (.A1(_07898_),
    .A2(_07950_),
    .B1(_07997_),
    .B2(_08204_),
    .X(_08205_));
 sky130_fd_sc_hd__and4_1 _14547_ (.A(_07943_),
    .B(_07946_),
    .C(_07950_),
    .D(_08162_),
    .X(_08206_));
 sky130_fd_sc_hd__nand2_1 _14548_ (.A(_07988_),
    .B(_08206_),
    .Y(_08207_));
 sky130_fd_sc_hd__a32o_1 _14549_ (.A1(_08203_),
    .A2(_08205_),
    .A3(_08207_),
    .B1(_07905_),
    .B2(\reg_next_pc[19] ),
    .X(_01011_));
 sky130_fd_sc_hd__nor2_1 _14550_ (.A(_07952_),
    .B(_08206_),
    .Y(_08208_));
 sky130_fd_sc_hd__and2_1 _14551_ (.A(_07952_),
    .B(_08206_),
    .X(_08209_));
 sky130_fd_sc_hd__nor2_1 _14552_ (.A(_08208_),
    .B(_08209_),
    .Y(_08210_));
 sky130_fd_sc_hd__a32o_1 _14553_ (.A1(_07898_),
    .A2(_07952_),
    .A3(_08050_),
    .B1(_07904_),
    .B2(\reg_next_pc[20] ),
    .X(_08211_));
 sky130_fd_sc_hd__buf_2 _14554_ (.A(\decoded_imm_j[20] ),
    .X(_08212_));
 sky130_fd_sc_hd__xnor2_1 _14555_ (.A(_08212_),
    .B(_07952_),
    .Y(_08213_));
 sky130_fd_sc_hd__a21oi_1 _14556_ (.A1(_08196_),
    .A2(_08201_),
    .B1(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__a31o_1 _14557_ (.A1(_08196_),
    .A2(_08201_),
    .A3(_08213_),
    .B1(_08055_),
    .X(_08215_));
 sky130_fd_sc_hd__nor2_1 _14558_ (.A(_08214_),
    .B(_08215_),
    .Y(_08216_));
 sky130_fd_sc_hd__a211o_1 _14559_ (.A1(_08121_),
    .A2(_08210_),
    .B1(_08211_),
    .C1(_08216_),
    .X(_01012_));
 sky130_fd_sc_hd__or2_1 _14560_ (.A(_07998_),
    .B(_08209_),
    .X(_08217_));
 sky130_fd_sc_hd__a22o_1 _14561_ (.A1(_03294_),
    .A2(_07954_),
    .B1(_07997_),
    .B2(_08217_),
    .X(_08218_));
 sky130_fd_sc_hd__xnor2_1 _14562_ (.A(_08212_),
    .B(_07954_),
    .Y(_08219_));
 sky130_fd_sc_hd__or2_1 _14563_ (.A(_08198_),
    .B(_08213_),
    .X(_08220_));
 sky130_fd_sc_hd__clkbuf_4 _14564_ (.A(_08212_),
    .X(_08221_));
 sky130_fd_sc_hd__a22o_1 _14565_ (.A1(\decoded_imm_j[19] ),
    .A2(_07950_),
    .B1(_07952_),
    .B2(_08212_),
    .X(_08222_));
 sky130_fd_sc_hd__o21ai_1 _14566_ (.A1(_08221_),
    .A2(_07952_),
    .B1(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__o31a_1 _14567_ (.A1(_08187_),
    .A2(_08199_),
    .A3(_08220_),
    .B1(_08223_),
    .X(_08224_));
 sky130_fd_sc_hd__o31a_1 _14568_ (.A1(_08180_),
    .A2(_08189_),
    .A3(_08220_),
    .B1(_08224_),
    .X(_08225_));
 sky130_fd_sc_hd__or2_1 _14569_ (.A(_08219_),
    .B(_08225_),
    .X(_08226_));
 sky130_fd_sc_hd__nand2_1 _14570_ (.A(_08219_),
    .B(_08225_),
    .Y(_08227_));
 sky130_fd_sc_hd__nand2_1 _14571_ (.A(_08226_),
    .B(_08227_),
    .Y(_08228_));
 sky130_fd_sc_hd__and3_1 _14572_ (.A(_07954_),
    .B(_07988_),
    .C(_08209_),
    .X(_08229_));
 sky130_fd_sc_hd__a21oi_1 _14573_ (.A1(_08012_),
    .A2(_08228_),
    .B1(_08229_),
    .Y(_08230_));
 sky130_fd_sc_hd__a22o_1 _14574_ (.A1(\reg_next_pc[21] ),
    .A2(_07948_),
    .B1(_08218_),
    .B2(_08230_),
    .X(_01013_));
 sky130_fd_sc_hd__xnor2_1 _14575_ (.A(_08212_),
    .B(_07956_),
    .Y(_08231_));
 sky130_fd_sc_hd__buf_4 _14576_ (.A(_08221_),
    .X(_08232_));
 sky130_fd_sc_hd__a21bo_1 _14577_ (.A1(_08232_),
    .A2(_07954_),
    .B1_N(_08226_),
    .X(_08233_));
 sky130_fd_sc_hd__xnor2_1 _14578_ (.A(_08231_),
    .B(_08233_),
    .Y(_08234_));
 sky130_fd_sc_hd__a32o_1 _14579_ (.A1(_07898_),
    .A2(_07956_),
    .A3(_08050_),
    .B1(_07904_),
    .B2(\reg_next_pc[22] ),
    .X(_08235_));
 sky130_fd_sc_hd__and3_1 _14580_ (.A(_07954_),
    .B(_07956_),
    .C(_08209_),
    .X(_08236_));
 sky130_fd_sc_hd__a31o_1 _14581_ (.A1(_07952_),
    .A2(_07954_),
    .A3(_08206_),
    .B1(_07956_),
    .X(_08237_));
 sky130_fd_sc_hd__and3b_1 _14582_ (.A_N(_08236_),
    .B(_08121_),
    .C(_08237_),
    .X(_08238_));
 sky130_fd_sc_hd__a211o_1 _14583_ (.A1(_08071_),
    .A2(_08234_),
    .B1(_08235_),
    .C1(_08238_),
    .X(_01014_));
 sky130_fd_sc_hd__nand2_1 _14584_ (.A(_08212_),
    .B(_07958_),
    .Y(_08239_));
 sky130_fd_sc_hd__or2_1 _14585_ (.A(_08212_),
    .B(_07958_),
    .X(_08240_));
 sky130_fd_sc_hd__nand2_1 _14586_ (.A(_08239_),
    .B(_08240_),
    .Y(_08241_));
 sky130_fd_sc_hd__o21ai_1 _14587_ (.A1(_07954_),
    .A2(_07956_),
    .B1(_08221_),
    .Y(_08242_));
 sky130_fd_sc_hd__o21a_1 _14588_ (.A1(_08226_),
    .A2(_08231_),
    .B1(_08242_),
    .X(_08243_));
 sky130_fd_sc_hd__o21ai_1 _14589_ (.A1(_08241_),
    .A2(_08243_),
    .B1(_08071_),
    .Y(_08244_));
 sky130_fd_sc_hd__a21oi_1 _14590_ (.A1(_08241_),
    .A2(_08243_),
    .B1(_08244_),
    .Y(_08245_));
 sky130_fd_sc_hd__nand2_1 _14591_ (.A(_07958_),
    .B(_08236_),
    .Y(_08246_));
 sky130_fd_sc_hd__or2_1 _14592_ (.A(_07958_),
    .B(_08236_),
    .X(_08247_));
 sky130_fd_sc_hd__and2_1 _14593_ (.A(_08246_),
    .B(_08247_),
    .X(_08248_));
 sky130_fd_sc_hd__a22o_1 _14594_ (.A1(_07958_),
    .A2(_07994_),
    .B1(_08248_),
    .B2(_07984_),
    .X(_08249_));
 sky130_fd_sc_hd__a21o_1 _14595_ (.A1(_03379_),
    .A2(_08248_),
    .B1(_08249_),
    .X(_08250_));
 sky130_fd_sc_hd__and3_1 _14596_ (.A(_03293_),
    .B(_07958_),
    .C(_07992_),
    .X(_08251_));
 sky130_fd_sc_hd__a221o_1 _14597_ (.A1(\reg_next_pc[23] ),
    .A2(_07903_),
    .B1(_08250_),
    .B2(_03378_),
    .C1(_08251_),
    .X(_08252_));
 sky130_fd_sc_hd__or2_1 _14598_ (.A(_08245_),
    .B(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__clkbuf_1 _14599_ (.A(_08253_),
    .X(_01015_));
 sky130_fd_sc_hd__xnor2_1 _14600_ (.A(_08212_),
    .B(_07959_),
    .Y(_08254_));
 sky130_fd_sc_hd__o21ai_1 _14601_ (.A1(_08241_),
    .A2(_08243_),
    .B1(_08239_),
    .Y(_08255_));
 sky130_fd_sc_hd__xnor2_1 _14602_ (.A(_08254_),
    .B(_08255_),
    .Y(_08256_));
 sky130_fd_sc_hd__o211ai_4 _14603_ (.A1(_05941_),
    .A2(_06286_),
    .B1(_07944_),
    .C1(_05922_),
    .Y(_08257_));
 sky130_fd_sc_hd__nor2_1 _14604_ (.A(_08257_),
    .B(_08246_),
    .Y(_08258_));
 sky130_fd_sc_hd__o32a_1 _14605_ (.A1(_07754_),
    .A2(_08257_),
    .A3(_07984_),
    .B1(_08035_),
    .B2(_08258_),
    .X(_08259_));
 sky130_fd_sc_hd__a21oi_1 _14606_ (.A1(_08257_),
    .A2(_08246_),
    .B1(_08259_),
    .Y(_08260_));
 sky130_fd_sc_hd__o211a_1 _14607_ (.A1(_03195_),
    .A2(_03363_),
    .B1(_07959_),
    .C1(_07898_),
    .X(_08261_));
 sky130_fd_sc_hd__a221o_1 _14608_ (.A1(\reg_next_pc[24] ),
    .A2(_07904_),
    .B1(_08260_),
    .B2(_03378_),
    .C1(_08261_),
    .X(_08262_));
 sky130_fd_sc_hd__a21o_1 _14609_ (.A1(_08071_),
    .A2(_08256_),
    .B1(_08262_),
    .X(_01016_));
 sky130_fd_sc_hd__and2_1 _14610_ (.A(_07961_),
    .B(_08258_),
    .X(_08263_));
 sky130_fd_sc_hd__nand2_1 _14611_ (.A(_07988_),
    .B(_08263_),
    .Y(_08264_));
 sky130_fd_sc_hd__or4_1 _14612_ (.A(_08219_),
    .B(_08231_),
    .C(_08241_),
    .D(_08254_),
    .X(_08265_));
 sky130_fd_sc_hd__o21ai_1 _14613_ (.A1(_07958_),
    .A2(_07959_),
    .B1(_08221_),
    .Y(_08266_));
 sky130_fd_sc_hd__o211a_1 _14614_ (.A1(_08225_),
    .A2(_08265_),
    .B1(_08266_),
    .C1(_08242_),
    .X(_08267_));
 sky130_fd_sc_hd__and2_1 _14615_ (.A(_07942_),
    .B(_07961_),
    .X(_08268_));
 sky130_fd_sc_hd__nand2_1 _14616_ (.A(_08221_),
    .B(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__or2_1 _14617_ (.A(_08221_),
    .B(_08268_),
    .X(_08270_));
 sky130_fd_sc_hd__nand2_1 _14618_ (.A(_08269_),
    .B(_08270_),
    .Y(_08271_));
 sky130_fd_sc_hd__or2_2 _14619_ (.A(_08267_),
    .B(_08271_),
    .X(_08272_));
 sky130_fd_sc_hd__nand2_1 _14620_ (.A(_08267_),
    .B(_08271_),
    .Y(_08273_));
 sky130_fd_sc_hd__nand2_1 _14621_ (.A(_08272_),
    .B(_08273_),
    .Y(_08274_));
 sky130_fd_sc_hd__o21a_1 _14622_ (.A1(_07998_),
    .A2(_08258_),
    .B1(_07997_),
    .X(_08275_));
 sky130_fd_sc_hd__o2bb2a_1 _14623_ (.A1_N(_08012_),
    .A2_N(_08274_),
    .B1(_08275_),
    .B2(_07962_),
    .X(_08276_));
 sky130_fd_sc_hd__a22o_1 _14624_ (.A1(\reg_next_pc[25] ),
    .A2(_07948_),
    .B1(_08264_),
    .B2(_08276_),
    .X(_01017_));
 sky130_fd_sc_hd__and3_1 _14625_ (.A(_07961_),
    .B(_07964_),
    .C(_08258_),
    .X(_08277_));
 sky130_fd_sc_hd__nor2_1 _14626_ (.A(_08035_),
    .B(_08277_),
    .Y(_08278_));
 sky130_fd_sc_hd__or2_1 _14627_ (.A(_08050_),
    .B(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__xnor2_2 _14628_ (.A(_08221_),
    .B(_07964_),
    .Y(_08280_));
 sky130_fd_sc_hd__a21oi_1 _14629_ (.A1(_08269_),
    .A2(_08272_),
    .B1(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__a31o_1 _14630_ (.A1(_08269_),
    .A2(_08272_),
    .A3(_08280_),
    .B1(_08097_),
    .X(_08282_));
 sky130_fd_sc_hd__a2bb2o_1 _14631_ (.A1_N(_08281_),
    .A2_N(_08282_),
    .B1(_08278_),
    .B2(_08263_),
    .X(_08283_));
 sky130_fd_sc_hd__a22o_1 _14632_ (.A1(\reg_next_pc[26] ),
    .A2(_07947_),
    .B1(_08283_),
    .B2(_08033_),
    .X(_08284_));
 sky130_fd_sc_hd__a31o_1 _14633_ (.A1(_07899_),
    .A2(_07964_),
    .A3(_08279_),
    .B1(_08284_),
    .X(_01018_));
 sky130_fd_sc_hd__or2_1 _14634_ (.A(_07998_),
    .B(_08277_),
    .X(_08285_));
 sky130_fd_sc_hd__a22o_1 _14635_ (.A1(_03294_),
    .A2(_07966_),
    .B1(_07997_),
    .B2(_08285_),
    .X(_08286_));
 sky130_fd_sc_hd__xnor2_1 _14636_ (.A(_08221_),
    .B(_07966_),
    .Y(_08287_));
 sky130_fd_sc_hd__o21ai_2 _14637_ (.A1(_08268_),
    .A2(_07964_),
    .B1(_08232_),
    .Y(_08288_));
 sky130_fd_sc_hd__o21a_1 _14638_ (.A1(_08272_),
    .A2(_08280_),
    .B1(_08288_),
    .X(_08289_));
 sky130_fd_sc_hd__nor2_1 _14639_ (.A(_08287_),
    .B(_08289_),
    .Y(_08290_));
 sky130_fd_sc_hd__and2_1 _14640_ (.A(_08287_),
    .B(_08289_),
    .X(_08291_));
 sky130_fd_sc_hd__or2_1 _14641_ (.A(_08290_),
    .B(_08291_),
    .X(_08292_));
 sky130_fd_sc_hd__and3_1 _14642_ (.A(_07966_),
    .B(_07988_),
    .C(_08277_),
    .X(_08293_));
 sky130_fd_sc_hd__a21oi_1 _14643_ (.A1(_08012_),
    .A2(_08292_),
    .B1(_08293_),
    .Y(_08294_));
 sky130_fd_sc_hd__a22o_1 _14644_ (.A1(\reg_next_pc[27] ),
    .A2(_07948_),
    .B1(_08286_),
    .B2(_08294_),
    .X(_01019_));
 sky130_fd_sc_hd__xnor2_1 _14645_ (.A(_08221_),
    .B(_07967_),
    .Y(_08295_));
 sky130_fd_sc_hd__a21oi_1 _14646_ (.A1(_08232_),
    .A2(_07966_),
    .B1(_08290_),
    .Y(_08296_));
 sky130_fd_sc_hd__a21oi_1 _14647_ (.A1(_08295_),
    .A2(_08296_),
    .B1(_08055_),
    .Y(_08297_));
 sky130_fd_sc_hd__o21a_1 _14648_ (.A1(_08295_),
    .A2(_08296_),
    .B1(_08297_),
    .X(_08298_));
 sky130_fd_sc_hd__a32o_1 _14649_ (.A1(_03293_),
    .A2(_07967_),
    .A3(_07995_),
    .B1(_07904_),
    .B2(\reg_next_pc[28] ),
    .X(_08299_));
 sky130_fd_sc_hd__a21oi_1 _14650_ (.A1(_07966_),
    .A2(_08277_),
    .B1(_07967_),
    .Y(_08300_));
 sky130_fd_sc_hd__and3_1 _14651_ (.A(_07966_),
    .B(_07967_),
    .C(_08277_),
    .X(_08301_));
 sky130_fd_sc_hd__or3b_1 _14652_ (.A(_08300_),
    .B(_08301_),
    .C_N(_08121_),
    .X(_08302_));
 sky130_fd_sc_hd__or3b_1 _14653_ (.A(_08298_),
    .B(_08299_),
    .C_N(_08302_),
    .X(_08303_));
 sky130_fd_sc_hd__clkbuf_1 _14654_ (.A(_08303_),
    .X(_01020_));
 sky130_fd_sc_hd__or2_1 _14655_ (.A(_07998_),
    .B(_08301_),
    .X(_08304_));
 sky130_fd_sc_hd__a22o_1 _14656_ (.A1(_03294_),
    .A2(_07968_),
    .B1(_07997_),
    .B2(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__or4_1 _14657_ (.A(_08272_),
    .B(_08280_),
    .C(_08287_),
    .D(_08295_),
    .X(_08306_));
 sky130_fd_sc_hd__o21ai_1 _14658_ (.A1(_07966_),
    .A2(_07967_),
    .B1(_08232_),
    .Y(_08307_));
 sky130_fd_sc_hd__and3_1 _14659_ (.A(_08288_),
    .B(_08306_),
    .C(_08307_),
    .X(_08308_));
 sky130_fd_sc_hd__nand2_1 _14660_ (.A(_08232_),
    .B(_07968_),
    .Y(_08309_));
 sky130_fd_sc_hd__or2_1 _14661_ (.A(_08221_),
    .B(_07968_),
    .X(_08310_));
 sky130_fd_sc_hd__nand2_1 _14662_ (.A(_08309_),
    .B(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__xnor2_1 _14663_ (.A(_08308_),
    .B(_08311_),
    .Y(_08312_));
 sky130_fd_sc_hd__nand2_1 _14664_ (.A(_07968_),
    .B(_08301_),
    .Y(_08313_));
 sky130_fd_sc_hd__o2bb2a_1 _14665_ (.A1_N(_08012_),
    .A2_N(_08312_),
    .B1(_08313_),
    .B2(_08120_),
    .X(_08314_));
 sky130_fd_sc_hd__a22o_1 _14666_ (.A1(\reg_next_pc[29] ),
    .A2(_07948_),
    .B1(_08305_),
    .B2(_08314_),
    .X(_01021_));
 sky130_fd_sc_hd__a31o_1 _14667_ (.A1(_08288_),
    .A2(_08306_),
    .A3(_08307_),
    .B1(_08311_),
    .X(_08315_));
 sky130_fd_sc_hd__nand2_1 _14668_ (.A(_08232_),
    .B(_07969_),
    .Y(_08316_));
 sky130_fd_sc_hd__or2_1 _14669_ (.A(_08232_),
    .B(_07969_),
    .X(_08317_));
 sky130_fd_sc_hd__nand2_1 _14670_ (.A(_08316_),
    .B(_08317_),
    .Y(_08318_));
 sky130_fd_sc_hd__a21oi_1 _14671_ (.A1(_08309_),
    .A2(_08315_),
    .B1(_08318_),
    .Y(_08319_));
 sky130_fd_sc_hd__a31o_1 _14672_ (.A1(_08309_),
    .A2(_08315_),
    .A3(_08318_),
    .B1(_08055_),
    .X(_08320_));
 sky130_fd_sc_hd__a21oi_1 _14673_ (.A1(_07968_),
    .A2(_08301_),
    .B1(_07969_),
    .Y(_08321_));
 sky130_fd_sc_hd__and3_1 _14674_ (.A(_07968_),
    .B(_07969_),
    .C(_08301_),
    .X(_08322_));
 sky130_fd_sc_hd__nor2_1 _14675_ (.A(_08321_),
    .B(_08322_),
    .Y(_08323_));
 sky130_fd_sc_hd__a32o_1 _14676_ (.A1(_07898_),
    .A2(_07969_),
    .A3(_08050_),
    .B1(_07904_),
    .B2(\reg_next_pc[30] ),
    .X(_08324_));
 sky130_fd_sc_hd__a21oi_1 _14677_ (.A1(_08121_),
    .A2(_08323_),
    .B1(_08324_),
    .Y(_08325_));
 sky130_fd_sc_hd__o21ai_1 _14678_ (.A1(_08319_),
    .A2(_08320_),
    .B1(_08325_),
    .Y(_01022_));
 sky130_fd_sc_hd__a21o_1 _14679_ (.A1(_03294_),
    .A2(_07971_),
    .B1(_08033_),
    .X(_08326_));
 sky130_fd_sc_hd__nand2_1 _14680_ (.A(_07971_),
    .B(_08322_),
    .Y(_08327_));
 sky130_fd_sc_hd__o21a_1 _14681_ (.A1(_07971_),
    .A2(_08322_),
    .B1(_07986_),
    .X(_08328_));
 sky130_fd_sc_hd__o31a_1 _14682_ (.A1(_03195_),
    .A2(_03363_),
    .A3(_07971_),
    .B1(_08050_),
    .X(_08329_));
 sky130_fd_sc_hd__o211a_1 _14683_ (.A1(_08315_),
    .A2(_08318_),
    .B1(_08316_),
    .C1(_08309_),
    .X(_08330_));
 sky130_fd_sc_hd__xnor2_1 _14684_ (.A(_08232_),
    .B(_07971_),
    .Y(_08331_));
 sky130_fd_sc_hd__a21oi_1 _14685_ (.A1(_08330_),
    .A2(_08331_),
    .B1(_08097_),
    .Y(_08332_));
 sky130_fd_sc_hd__o21a_1 _14686_ (.A1(_08330_),
    .A2(_08331_),
    .B1(_08332_),
    .X(_08333_));
 sky130_fd_sc_hd__a211o_1 _14687_ (.A1(_08327_),
    .A2(_08328_),
    .B1(_08329_),
    .C1(_08333_),
    .X(_08334_));
 sky130_fd_sc_hd__a22o_1 _14688_ (.A1(\reg_next_pc[31] ),
    .A2(_07948_),
    .B1(_08326_),
    .B2(_08334_),
    .X(_01023_));
 sky130_fd_sc_hd__clkbuf_4 _14689_ (.A(_03240_),
    .X(_08335_));
 sky130_fd_sc_hd__nor2_1 _14690_ (.A(_08335_),
    .B(\count_cycle[0] ),
    .Y(_01024_));
 sky130_fd_sc_hd__o21ai_1 _14691_ (.A1(\count_cycle[0] ),
    .A2(\count_cycle[1] ),
    .B1(_07675_),
    .Y(_08336_));
 sky130_fd_sc_hd__a21oi_1 _14692_ (.A1(\count_cycle[0] ),
    .A2(\count_cycle[1] ),
    .B1(_08336_),
    .Y(_01025_));
 sky130_fd_sc_hd__and3_1 _14693_ (.A(\count_cycle[0] ),
    .B(\count_cycle[1] ),
    .C(\count_cycle[2] ),
    .X(_08337_));
 sky130_fd_sc_hd__a21o_1 _14694_ (.A1(\count_cycle[0] ),
    .A2(\count_cycle[1] ),
    .B1(\count_cycle[2] ),
    .X(_08338_));
 sky130_fd_sc_hd__and3b_1 _14695_ (.A_N(_08337_),
    .B(_07815_),
    .C(_08338_),
    .X(_08339_));
 sky130_fd_sc_hd__clkbuf_1 _14696_ (.A(_08339_),
    .X(_01026_));
 sky130_fd_sc_hd__and4_2 _14697_ (.A(\count_cycle[0] ),
    .B(\count_cycle[1] ),
    .C(\count_cycle[2] ),
    .D(\count_cycle[3] ),
    .X(_08340_));
 sky130_fd_sc_hd__o21ai_1 _14698_ (.A1(\count_cycle[3] ),
    .A2(_08337_),
    .B1(_07877_),
    .Y(_08341_));
 sky130_fd_sc_hd__nor2_1 _14699_ (.A(_08340_),
    .B(_08341_),
    .Y(_01027_));
 sky130_fd_sc_hd__a21oi_1 _14700_ (.A1(\count_cycle[4] ),
    .A2(_08340_),
    .B1(_07826_),
    .Y(_08342_));
 sky130_fd_sc_hd__o21a_1 _14701_ (.A1(\count_cycle[4] ),
    .A2(_08340_),
    .B1(_08342_),
    .X(_01028_));
 sky130_fd_sc_hd__and3_1 _14702_ (.A(\count_cycle[4] ),
    .B(\count_cycle[5] ),
    .C(_08340_),
    .X(_08343_));
 sky130_fd_sc_hd__a21o_1 _14703_ (.A1(\count_cycle[4] ),
    .A2(_08340_),
    .B1(\count_cycle[5] ),
    .X(_08344_));
 sky130_fd_sc_hd__and3b_1 _14704_ (.A_N(_08343_),
    .B(_07815_),
    .C(_08344_),
    .X(_08345_));
 sky130_fd_sc_hd__clkbuf_1 _14705_ (.A(_08345_),
    .X(_01029_));
 sky130_fd_sc_hd__and4_2 _14706_ (.A(\count_cycle[4] ),
    .B(\count_cycle[5] ),
    .C(\count_cycle[6] ),
    .D(_08340_),
    .X(_08346_));
 sky130_fd_sc_hd__o21ai_1 _14707_ (.A1(\count_cycle[6] ),
    .A2(_08343_),
    .B1(_07877_),
    .Y(_08347_));
 sky130_fd_sc_hd__nor2_1 _14708_ (.A(_08346_),
    .B(_08347_),
    .Y(_01030_));
 sky130_fd_sc_hd__a21oi_1 _14709_ (.A1(\count_cycle[7] ),
    .A2(_08346_),
    .B1(_07826_),
    .Y(_08348_));
 sky130_fd_sc_hd__o21a_1 _14710_ (.A1(\count_cycle[7] ),
    .A2(_08346_),
    .B1(_08348_),
    .X(_01031_));
 sky130_fd_sc_hd__and3_1 _14711_ (.A(\count_cycle[7] ),
    .B(\count_cycle[8] ),
    .C(_08346_),
    .X(_08349_));
 sky130_fd_sc_hd__clkbuf_4 _14712_ (.A(_03304_),
    .X(_08350_));
 sky130_fd_sc_hd__a21o_1 _14713_ (.A1(\count_cycle[7] ),
    .A2(_08346_),
    .B1(\count_cycle[8] ),
    .X(_08351_));
 sky130_fd_sc_hd__and3b_1 _14714_ (.A_N(_08349_),
    .B(_08350_),
    .C(_08351_),
    .X(_08352_));
 sky130_fd_sc_hd__clkbuf_1 _14715_ (.A(_08352_),
    .X(_01032_));
 sky130_fd_sc_hd__and4_2 _14716_ (.A(\count_cycle[7] ),
    .B(\count_cycle[8] ),
    .C(\count_cycle[9] ),
    .D(_08346_),
    .X(_08353_));
 sky130_fd_sc_hd__o21ai_1 _14717_ (.A1(\count_cycle[9] ),
    .A2(_08349_),
    .B1(_07877_),
    .Y(_08354_));
 sky130_fd_sc_hd__nor2_1 _14718_ (.A(_08353_),
    .B(_08354_),
    .Y(_01033_));
 sky130_fd_sc_hd__a21oi_1 _14719_ (.A1(\count_cycle[10] ),
    .A2(_08353_),
    .B1(_07826_),
    .Y(_08355_));
 sky130_fd_sc_hd__o21a_1 _14720_ (.A1(\count_cycle[10] ),
    .A2(_08353_),
    .B1(_08355_),
    .X(_01034_));
 sky130_fd_sc_hd__and3_1 _14721_ (.A(\count_cycle[10] ),
    .B(\count_cycle[11] ),
    .C(_08353_),
    .X(_08356_));
 sky130_fd_sc_hd__a21o_1 _14722_ (.A1(\count_cycle[10] ),
    .A2(_08353_),
    .B1(\count_cycle[11] ),
    .X(_08357_));
 sky130_fd_sc_hd__and3b_1 _14723_ (.A_N(_08356_),
    .B(_08350_),
    .C(_08357_),
    .X(_08358_));
 sky130_fd_sc_hd__clkbuf_1 _14724_ (.A(_08358_),
    .X(_01035_));
 sky130_fd_sc_hd__and4_2 _14725_ (.A(\count_cycle[10] ),
    .B(\count_cycle[11] ),
    .C(\count_cycle[12] ),
    .D(_08353_),
    .X(_08359_));
 sky130_fd_sc_hd__o21ai_1 _14726_ (.A1(\count_cycle[12] ),
    .A2(_08356_),
    .B1(_07877_),
    .Y(_08360_));
 sky130_fd_sc_hd__nor2_1 _14727_ (.A(_08359_),
    .B(_08360_),
    .Y(_01036_));
 sky130_fd_sc_hd__a21oi_1 _14728_ (.A1(\count_cycle[13] ),
    .A2(_08359_),
    .B1(_07826_),
    .Y(_08361_));
 sky130_fd_sc_hd__o21a_1 _14729_ (.A1(\count_cycle[13] ),
    .A2(_08359_),
    .B1(_08361_),
    .X(_01037_));
 sky130_fd_sc_hd__and3_1 _14730_ (.A(\count_cycle[13] ),
    .B(\count_cycle[14] ),
    .C(_08359_),
    .X(_08362_));
 sky130_fd_sc_hd__a21o_1 _14731_ (.A1(\count_cycle[13] ),
    .A2(_08359_),
    .B1(\count_cycle[14] ),
    .X(_08363_));
 sky130_fd_sc_hd__and3b_1 _14732_ (.A_N(_08362_),
    .B(_08350_),
    .C(_08363_),
    .X(_08364_));
 sky130_fd_sc_hd__clkbuf_1 _14733_ (.A(_08364_),
    .X(_01038_));
 sky130_fd_sc_hd__and4_2 _14734_ (.A(\count_cycle[13] ),
    .B(\count_cycle[14] ),
    .C(\count_cycle[15] ),
    .D(_08359_),
    .X(_08365_));
 sky130_fd_sc_hd__o21ai_1 _14735_ (.A1(\count_cycle[15] ),
    .A2(_08362_),
    .B1(_07877_),
    .Y(_08366_));
 sky130_fd_sc_hd__nor2_1 _14736_ (.A(_08365_),
    .B(_08366_),
    .Y(_01039_));
 sky130_fd_sc_hd__a21oi_1 _14737_ (.A1(\count_cycle[16] ),
    .A2(_08365_),
    .B1(_07826_),
    .Y(_08367_));
 sky130_fd_sc_hd__o21a_1 _14738_ (.A1(\count_cycle[16] ),
    .A2(_08365_),
    .B1(_08367_),
    .X(_01040_));
 sky130_fd_sc_hd__and3_1 _14739_ (.A(\count_cycle[16] ),
    .B(\count_cycle[17] ),
    .C(_08365_),
    .X(_08368_));
 sky130_fd_sc_hd__a21o_1 _14740_ (.A1(\count_cycle[16] ),
    .A2(_08365_),
    .B1(\count_cycle[17] ),
    .X(_01712_));
 sky130_fd_sc_hd__and3b_1 _14741_ (.A_N(_08368_),
    .B(_08350_),
    .C(_01712_),
    .X(_01713_));
 sky130_fd_sc_hd__clkbuf_1 _14742_ (.A(_01713_),
    .X(_01041_));
 sky130_fd_sc_hd__buf_4 _14743_ (.A(_03239_),
    .X(_01714_));
 sky130_fd_sc_hd__and4_2 _14744_ (.A(\count_cycle[16] ),
    .B(\count_cycle[17] ),
    .C(\count_cycle[18] ),
    .D(_08365_),
    .X(_01715_));
 sky130_fd_sc_hd__nor2_1 _14745_ (.A(_01714_),
    .B(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__o21a_1 _14746_ (.A1(\count_cycle[18] ),
    .A2(_08368_),
    .B1(_01716_),
    .X(_01042_));
 sky130_fd_sc_hd__clkbuf_4 _14747_ (.A(_03239_),
    .X(_01717_));
 sky130_fd_sc_hd__a21oi_1 _14748_ (.A1(\count_cycle[19] ),
    .A2(_01715_),
    .B1(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__o21a_1 _14749_ (.A1(\count_cycle[19] ),
    .A2(_01715_),
    .B1(_01718_),
    .X(_01043_));
 sky130_fd_sc_hd__and3_1 _14750_ (.A(\count_cycle[19] ),
    .B(\count_cycle[20] ),
    .C(_01715_),
    .X(_01719_));
 sky130_fd_sc_hd__a21o_1 _14751_ (.A1(\count_cycle[19] ),
    .A2(_01715_),
    .B1(\count_cycle[20] ),
    .X(_01720_));
 sky130_fd_sc_hd__and3b_1 _14752_ (.A_N(_01719_),
    .B(_08350_),
    .C(_01720_),
    .X(_01721_));
 sky130_fd_sc_hd__clkbuf_1 _14753_ (.A(_01721_),
    .X(_01044_));
 sky130_fd_sc_hd__and4_2 _14754_ (.A(\count_cycle[19] ),
    .B(\count_cycle[20] ),
    .C(\count_cycle[21] ),
    .D(_01715_),
    .X(_01722_));
 sky130_fd_sc_hd__clkbuf_4 _14755_ (.A(_06053_),
    .X(_01723_));
 sky130_fd_sc_hd__o21ai_1 _14756_ (.A1(\count_cycle[21] ),
    .A2(_01719_),
    .B1(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__nor2_1 _14757_ (.A(_01722_),
    .B(_01724_),
    .Y(_01045_));
 sky130_fd_sc_hd__a21oi_1 _14758_ (.A1(\count_cycle[22] ),
    .A2(_01722_),
    .B1(_01717_),
    .Y(_01725_));
 sky130_fd_sc_hd__o21a_1 _14759_ (.A1(\count_cycle[22] ),
    .A2(_01722_),
    .B1(_01725_),
    .X(_01046_));
 sky130_fd_sc_hd__and3_1 _14760_ (.A(\count_cycle[22] ),
    .B(\count_cycle[23] ),
    .C(_01722_),
    .X(_01726_));
 sky130_fd_sc_hd__a21o_1 _14761_ (.A1(\count_cycle[22] ),
    .A2(_01722_),
    .B1(\count_cycle[23] ),
    .X(_01727_));
 sky130_fd_sc_hd__and3b_1 _14762_ (.A_N(_01726_),
    .B(_08350_),
    .C(_01727_),
    .X(_01728_));
 sky130_fd_sc_hd__clkbuf_1 _14763_ (.A(_01728_),
    .X(_01047_));
 sky130_fd_sc_hd__and4_2 _14764_ (.A(\count_cycle[22] ),
    .B(\count_cycle[23] ),
    .C(\count_cycle[24] ),
    .D(_01722_),
    .X(_01729_));
 sky130_fd_sc_hd__o21ai_1 _14765_ (.A1(\count_cycle[24] ),
    .A2(_01726_),
    .B1(_01723_),
    .Y(_01730_));
 sky130_fd_sc_hd__nor2_1 _14766_ (.A(_01729_),
    .B(_01730_),
    .Y(_01048_));
 sky130_fd_sc_hd__a21oi_1 _14767_ (.A1(\count_cycle[25] ),
    .A2(_01729_),
    .B1(_01717_),
    .Y(_01731_));
 sky130_fd_sc_hd__o21a_1 _14768_ (.A1(\count_cycle[25] ),
    .A2(_01729_),
    .B1(_01731_),
    .X(_01049_));
 sky130_fd_sc_hd__and3_1 _14769_ (.A(\count_cycle[25] ),
    .B(\count_cycle[26] ),
    .C(_01729_),
    .X(_01732_));
 sky130_fd_sc_hd__a21o_1 _14770_ (.A1(\count_cycle[25] ),
    .A2(_01729_),
    .B1(\count_cycle[26] ),
    .X(_01733_));
 sky130_fd_sc_hd__and3b_1 _14771_ (.A_N(_01732_),
    .B(_08350_),
    .C(_01733_),
    .X(_01734_));
 sky130_fd_sc_hd__clkbuf_1 _14772_ (.A(_01734_),
    .X(_01050_));
 sky130_fd_sc_hd__and4_1 _14773_ (.A(\count_cycle[25] ),
    .B(\count_cycle[26] ),
    .C(\count_cycle[27] ),
    .D(_01729_),
    .X(_01735_));
 sky130_fd_sc_hd__clkbuf_2 _14774_ (.A(_01735_),
    .X(_01736_));
 sky130_fd_sc_hd__o21ai_1 _14775_ (.A1(\count_cycle[27] ),
    .A2(_01732_),
    .B1(_01723_),
    .Y(_01737_));
 sky130_fd_sc_hd__nor2_1 _14776_ (.A(_01736_),
    .B(_01737_),
    .Y(_01051_));
 sky130_fd_sc_hd__a21oi_1 _14777_ (.A1(\count_cycle[28] ),
    .A2(_01736_),
    .B1(_01717_),
    .Y(_01738_));
 sky130_fd_sc_hd__o21a_1 _14778_ (.A1(\count_cycle[28] ),
    .A2(_01736_),
    .B1(_01738_),
    .X(_01052_));
 sky130_fd_sc_hd__a21oi_1 _14779_ (.A1(\count_cycle[28] ),
    .A2(_01736_),
    .B1(\count_cycle[29] ),
    .Y(_01739_));
 sky130_fd_sc_hd__a31o_1 _14780_ (.A1(\count_cycle[28] ),
    .A2(\count_cycle[29] ),
    .A3(_01736_),
    .B1(_03240_),
    .X(_01740_));
 sky130_fd_sc_hd__nor2_1 _14781_ (.A(_01739_),
    .B(_01740_),
    .Y(_01053_));
 sky130_fd_sc_hd__and4_2 _14782_ (.A(\count_cycle[28] ),
    .B(\count_cycle[29] ),
    .C(\count_cycle[30] ),
    .D(_01736_),
    .X(_01741_));
 sky130_fd_sc_hd__a31o_1 _14783_ (.A1(\count_cycle[28] ),
    .A2(\count_cycle[29] ),
    .A3(_01736_),
    .B1(\count_cycle[30] ),
    .X(_01742_));
 sky130_fd_sc_hd__and3b_1 _14784_ (.A_N(_01741_),
    .B(_08350_),
    .C(_01742_),
    .X(_01743_));
 sky130_fd_sc_hd__clkbuf_1 _14785_ (.A(_01743_),
    .X(_01054_));
 sky130_fd_sc_hd__a21oi_1 _14786_ (.A1(\count_cycle[31] ),
    .A2(_01741_),
    .B1(_01717_),
    .Y(_01744_));
 sky130_fd_sc_hd__o21a_1 _14787_ (.A1(\count_cycle[31] ),
    .A2(_01741_),
    .B1(_01744_),
    .X(_01055_));
 sky130_fd_sc_hd__and3_1 _14788_ (.A(\count_cycle[32] ),
    .B(\count_cycle[31] ),
    .C(_01741_),
    .X(_01745_));
 sky130_fd_sc_hd__a21o_1 _14789_ (.A1(\count_cycle[31] ),
    .A2(_01741_),
    .B1(\count_cycle[32] ),
    .X(_01746_));
 sky130_fd_sc_hd__and3b_1 _14790_ (.A_N(_01745_),
    .B(_08350_),
    .C(_01746_),
    .X(_01747_));
 sky130_fd_sc_hd__clkbuf_1 _14791_ (.A(_01747_),
    .X(_01056_));
 sky130_fd_sc_hd__and4_2 _14792_ (.A(\count_cycle[32] ),
    .B(\count_cycle[33] ),
    .C(\count_cycle[31] ),
    .D(_01741_),
    .X(_01748_));
 sky130_fd_sc_hd__or2_1 _14793_ (.A(\count_cycle[33] ),
    .B(_01745_),
    .X(_01749_));
 sky130_fd_sc_hd__and3b_1 _14794_ (.A_N(_01748_),
    .B(_08350_),
    .C(_01749_),
    .X(_01750_));
 sky130_fd_sc_hd__clkbuf_1 _14795_ (.A(_01750_),
    .X(_01057_));
 sky130_fd_sc_hd__a21oi_1 _14796_ (.A1(\count_cycle[34] ),
    .A2(_01748_),
    .B1(_01717_),
    .Y(_01751_));
 sky130_fd_sc_hd__o21a_1 _14797_ (.A1(\count_cycle[34] ),
    .A2(_01748_),
    .B1(_01751_),
    .X(_01058_));
 sky130_fd_sc_hd__and3_1 _14798_ (.A(\count_cycle[34] ),
    .B(\count_cycle[35] ),
    .C(_01748_),
    .X(_01752_));
 sky130_fd_sc_hd__clkbuf_4 _14799_ (.A(_03304_),
    .X(_01753_));
 sky130_fd_sc_hd__a21o_1 _14800_ (.A1(\count_cycle[34] ),
    .A2(_01748_),
    .B1(\count_cycle[35] ),
    .X(_01754_));
 sky130_fd_sc_hd__and3b_1 _14801_ (.A_N(_01752_),
    .B(_01753_),
    .C(_01754_),
    .X(_01755_));
 sky130_fd_sc_hd__clkbuf_1 _14802_ (.A(_01755_),
    .X(_01059_));
 sky130_fd_sc_hd__and4_2 _14803_ (.A(\count_cycle[34] ),
    .B(\count_cycle[35] ),
    .C(\count_cycle[36] ),
    .D(_01748_),
    .X(_01756_));
 sky130_fd_sc_hd__o21ai_1 _14804_ (.A1(\count_cycle[36] ),
    .A2(_01752_),
    .B1(_01723_),
    .Y(_01757_));
 sky130_fd_sc_hd__nor2_1 _14805_ (.A(_01756_),
    .B(_01757_),
    .Y(_01060_));
 sky130_fd_sc_hd__a21oi_1 _14806_ (.A1(\count_cycle[37] ),
    .A2(_01756_),
    .B1(_01717_),
    .Y(_01758_));
 sky130_fd_sc_hd__o21a_1 _14807_ (.A1(\count_cycle[37] ),
    .A2(_01756_),
    .B1(_01758_),
    .X(_01061_));
 sky130_fd_sc_hd__and3_1 _14808_ (.A(\count_cycle[37] ),
    .B(\count_cycle[38] ),
    .C(_01756_),
    .X(_01759_));
 sky130_fd_sc_hd__a21o_1 _14809_ (.A1(\count_cycle[37] ),
    .A2(_01756_),
    .B1(\count_cycle[38] ),
    .X(_01760_));
 sky130_fd_sc_hd__and3b_1 _14810_ (.A_N(_01759_),
    .B(_01753_),
    .C(_01760_),
    .X(_01761_));
 sky130_fd_sc_hd__clkbuf_1 _14811_ (.A(_01761_),
    .X(_01062_));
 sky130_fd_sc_hd__and4_2 _14812_ (.A(\count_cycle[37] ),
    .B(\count_cycle[38] ),
    .C(\count_cycle[39] ),
    .D(_01756_),
    .X(_01762_));
 sky130_fd_sc_hd__o21ai_1 _14813_ (.A1(\count_cycle[39] ),
    .A2(_01759_),
    .B1(_01723_),
    .Y(_01763_));
 sky130_fd_sc_hd__nor2_1 _14814_ (.A(_01762_),
    .B(_01763_),
    .Y(_01063_));
 sky130_fd_sc_hd__a21oi_1 _14815_ (.A1(\count_cycle[40] ),
    .A2(_01762_),
    .B1(_01717_),
    .Y(_01764_));
 sky130_fd_sc_hd__o21a_1 _14816_ (.A1(\count_cycle[40] ),
    .A2(_01762_),
    .B1(_01764_),
    .X(_01064_));
 sky130_fd_sc_hd__and3_1 _14817_ (.A(\count_cycle[40] ),
    .B(\count_cycle[41] ),
    .C(_01762_),
    .X(_01765_));
 sky130_fd_sc_hd__a21o_1 _14818_ (.A1(\count_cycle[40] ),
    .A2(_01762_),
    .B1(\count_cycle[41] ),
    .X(_01766_));
 sky130_fd_sc_hd__and3b_1 _14819_ (.A_N(_01765_),
    .B(_01753_),
    .C(_01766_),
    .X(_01767_));
 sky130_fd_sc_hd__clkbuf_1 _14820_ (.A(_01767_),
    .X(_01065_));
 sky130_fd_sc_hd__and4_2 _14821_ (.A(\count_cycle[40] ),
    .B(\count_cycle[41] ),
    .C(\count_cycle[42] ),
    .D(_01762_),
    .X(_01768_));
 sky130_fd_sc_hd__o21ai_1 _14822_ (.A1(\count_cycle[42] ),
    .A2(_01765_),
    .B1(_01723_),
    .Y(_01769_));
 sky130_fd_sc_hd__nor2_1 _14823_ (.A(_01768_),
    .B(_01769_),
    .Y(_01066_));
 sky130_fd_sc_hd__a21oi_1 _14824_ (.A1(\count_cycle[43] ),
    .A2(_01768_),
    .B1(_01717_),
    .Y(_01770_));
 sky130_fd_sc_hd__o21a_1 _14825_ (.A1(\count_cycle[43] ),
    .A2(_01768_),
    .B1(_01770_),
    .X(_01067_));
 sky130_fd_sc_hd__and3_1 _14826_ (.A(\count_cycle[43] ),
    .B(\count_cycle[44] ),
    .C(_01768_),
    .X(_01771_));
 sky130_fd_sc_hd__a21o_1 _14827_ (.A1(\count_cycle[43] ),
    .A2(_01768_),
    .B1(\count_cycle[44] ),
    .X(_01772_));
 sky130_fd_sc_hd__and3b_1 _14828_ (.A_N(_01771_),
    .B(_01753_),
    .C(_01772_),
    .X(_01773_));
 sky130_fd_sc_hd__clkbuf_1 _14829_ (.A(_01773_),
    .X(_01068_));
 sky130_fd_sc_hd__and4_2 _14830_ (.A(\count_cycle[43] ),
    .B(\count_cycle[44] ),
    .C(\count_cycle[45] ),
    .D(_01768_),
    .X(_01774_));
 sky130_fd_sc_hd__o21ai_1 _14831_ (.A1(\count_cycle[45] ),
    .A2(_01771_),
    .B1(_01723_),
    .Y(_01775_));
 sky130_fd_sc_hd__nor2_1 _14832_ (.A(_01774_),
    .B(_01775_),
    .Y(_01069_));
 sky130_fd_sc_hd__a21oi_1 _14833_ (.A1(\count_cycle[46] ),
    .A2(_01774_),
    .B1(_01717_),
    .Y(_01776_));
 sky130_fd_sc_hd__o21a_1 _14834_ (.A1(\count_cycle[46] ),
    .A2(_01774_),
    .B1(_01776_),
    .X(_01070_));
 sky130_fd_sc_hd__and3_1 _14835_ (.A(\count_cycle[46] ),
    .B(\count_cycle[47] ),
    .C(_01774_),
    .X(_01777_));
 sky130_fd_sc_hd__a21o_1 _14836_ (.A1(\count_cycle[46] ),
    .A2(_01774_),
    .B1(\count_cycle[47] ),
    .X(_01778_));
 sky130_fd_sc_hd__and3b_1 _14837_ (.A_N(_01777_),
    .B(_01753_),
    .C(_01778_),
    .X(_01779_));
 sky130_fd_sc_hd__clkbuf_1 _14838_ (.A(_01779_),
    .X(_01071_));
 sky130_fd_sc_hd__and4_2 _14839_ (.A(\count_cycle[46] ),
    .B(\count_cycle[47] ),
    .C(\count_cycle[48] ),
    .D(_01774_),
    .X(_01780_));
 sky130_fd_sc_hd__o21ai_1 _14840_ (.A1(\count_cycle[48] ),
    .A2(_01777_),
    .B1(_01723_),
    .Y(_01781_));
 sky130_fd_sc_hd__nor2_1 _14841_ (.A(_01780_),
    .B(_01781_),
    .Y(_01072_));
 sky130_fd_sc_hd__a21oi_1 _14842_ (.A1(\count_cycle[49] ),
    .A2(_01780_),
    .B1(_01714_),
    .Y(_01782_));
 sky130_fd_sc_hd__o21a_1 _14843_ (.A1(\count_cycle[49] ),
    .A2(_01780_),
    .B1(_01782_),
    .X(_01073_));
 sky130_fd_sc_hd__and3_1 _14844_ (.A(\count_cycle[49] ),
    .B(\count_cycle[50] ),
    .C(_01780_),
    .X(_01783_));
 sky130_fd_sc_hd__a21o_1 _14845_ (.A1(\count_cycle[49] ),
    .A2(_01780_),
    .B1(\count_cycle[50] ),
    .X(_01784_));
 sky130_fd_sc_hd__and3b_1 _14846_ (.A_N(_01783_),
    .B(_01753_),
    .C(_01784_),
    .X(_01785_));
 sky130_fd_sc_hd__clkbuf_1 _14847_ (.A(_01785_),
    .X(_01074_));
 sky130_fd_sc_hd__and4_2 _14848_ (.A(\count_cycle[49] ),
    .B(\count_cycle[50] ),
    .C(\count_cycle[51] ),
    .D(_01780_),
    .X(_01786_));
 sky130_fd_sc_hd__o21ai_1 _14849_ (.A1(\count_cycle[51] ),
    .A2(_01783_),
    .B1(_01723_),
    .Y(_01787_));
 sky130_fd_sc_hd__nor2_1 _14850_ (.A(_01786_),
    .B(_01787_),
    .Y(_01075_));
 sky130_fd_sc_hd__a21oi_1 _14851_ (.A1(\count_cycle[52] ),
    .A2(_01786_),
    .B1(_01714_),
    .Y(_01788_));
 sky130_fd_sc_hd__o21a_1 _14852_ (.A1(\count_cycle[52] ),
    .A2(_01786_),
    .B1(_01788_),
    .X(_01076_));
 sky130_fd_sc_hd__and3_1 _14853_ (.A(\count_cycle[52] ),
    .B(\count_cycle[53] ),
    .C(_01786_),
    .X(_01789_));
 sky130_fd_sc_hd__a21o_1 _14854_ (.A1(\count_cycle[52] ),
    .A2(_01786_),
    .B1(\count_cycle[53] ),
    .X(_01790_));
 sky130_fd_sc_hd__and3b_1 _14855_ (.A_N(_01789_),
    .B(_01753_),
    .C(_01790_),
    .X(_01791_));
 sky130_fd_sc_hd__clkbuf_1 _14856_ (.A(_01791_),
    .X(_01077_));
 sky130_fd_sc_hd__and4_1 _14857_ (.A(\count_cycle[52] ),
    .B(\count_cycle[53] ),
    .C(\count_cycle[54] ),
    .D(_01786_),
    .X(_01792_));
 sky130_fd_sc_hd__o21ai_1 _14858_ (.A1(\count_cycle[54] ),
    .A2(_01789_),
    .B1(_01723_),
    .Y(_01793_));
 sky130_fd_sc_hd__nor2_1 _14859_ (.A(_01792_),
    .B(_01793_),
    .Y(_01078_));
 sky130_fd_sc_hd__a21oi_1 _14860_ (.A1(\count_cycle[55] ),
    .A2(_01792_),
    .B1(_01714_),
    .Y(_01794_));
 sky130_fd_sc_hd__o21a_1 _14861_ (.A1(\count_cycle[55] ),
    .A2(_01792_),
    .B1(_01794_),
    .X(_01079_));
 sky130_fd_sc_hd__and3_1 _14862_ (.A(\count_cycle[55] ),
    .B(\count_cycle[56] ),
    .C(_01792_),
    .X(_01795_));
 sky130_fd_sc_hd__a21o_1 _14863_ (.A1(\count_cycle[55] ),
    .A2(_01792_),
    .B1(\count_cycle[56] ),
    .X(_01796_));
 sky130_fd_sc_hd__and3b_1 _14864_ (.A_N(_01795_),
    .B(_01753_),
    .C(_01796_),
    .X(_01797_));
 sky130_fd_sc_hd__clkbuf_1 _14865_ (.A(_01797_),
    .X(_01080_));
 sky130_fd_sc_hd__and2_1 _14866_ (.A(\count_cycle[57] ),
    .B(_01795_),
    .X(_01798_));
 sky130_fd_sc_hd__o21ai_1 _14867_ (.A1(\count_cycle[57] ),
    .A2(_01795_),
    .B1(_07675_),
    .Y(_01799_));
 sky130_fd_sc_hd__nor2_1 _14868_ (.A(_01798_),
    .B(_01799_),
    .Y(_01081_));
 sky130_fd_sc_hd__a21oi_1 _14869_ (.A1(\count_cycle[58] ),
    .A2(_01798_),
    .B1(_01714_),
    .Y(_01800_));
 sky130_fd_sc_hd__o21a_1 _14870_ (.A1(\count_cycle[58] ),
    .A2(_01798_),
    .B1(_01800_),
    .X(_01082_));
 sky130_fd_sc_hd__and3_1 _14871_ (.A(\count_cycle[58] ),
    .B(\count_cycle[59] ),
    .C(_01798_),
    .X(_01801_));
 sky130_fd_sc_hd__a31o_1 _14872_ (.A1(\count_cycle[57] ),
    .A2(\count_cycle[58] ),
    .A3(_01795_),
    .B1(\count_cycle[59] ),
    .X(_01802_));
 sky130_fd_sc_hd__and3b_1 _14873_ (.A_N(_01801_),
    .B(_01753_),
    .C(_01802_),
    .X(_01803_));
 sky130_fd_sc_hd__clkbuf_1 _14874_ (.A(_01803_),
    .X(_01083_));
 sky130_fd_sc_hd__and2_1 _14875_ (.A(\count_cycle[60] ),
    .B(_01801_),
    .X(_01804_));
 sky130_fd_sc_hd__o21ai_1 _14876_ (.A1(\count_cycle[60] ),
    .A2(_01801_),
    .B1(_07675_),
    .Y(_01805_));
 sky130_fd_sc_hd__nor2_1 _14877_ (.A(_01804_),
    .B(_01805_),
    .Y(_01084_));
 sky130_fd_sc_hd__a31o_1 _14878_ (.A1(\count_cycle[60] ),
    .A2(\count_cycle[61] ),
    .A3(_01801_),
    .B1(_03240_),
    .X(_01806_));
 sky130_fd_sc_hd__o21ba_1 _14879_ (.A1(\count_cycle[61] ),
    .A2(_01804_),
    .B1_N(_01806_),
    .X(_01085_));
 sky130_fd_sc_hd__and3_1 _14880_ (.A(\count_cycle[61] ),
    .B(\count_cycle[62] ),
    .C(_01804_),
    .X(_01807_));
 sky130_fd_sc_hd__a31o_1 _14881_ (.A1(\count_cycle[60] ),
    .A2(\count_cycle[61] ),
    .A3(_01801_),
    .B1(\count_cycle[62] ),
    .X(_01808_));
 sky130_fd_sc_hd__and3b_1 _14882_ (.A_N(_01807_),
    .B(_01753_),
    .C(_01808_),
    .X(_01809_));
 sky130_fd_sc_hd__clkbuf_1 _14883_ (.A(_01809_),
    .X(_01086_));
 sky130_fd_sc_hd__a21oi_1 _14884_ (.A1(\count_cycle[63] ),
    .A2(_01807_),
    .B1(_01714_),
    .Y(_01810_));
 sky130_fd_sc_hd__o21a_1 _14885_ (.A1(\count_cycle[63] ),
    .A2(_01807_),
    .B1(_01810_),
    .X(_01087_));
 sky130_fd_sc_hd__nor2_1 _14886_ (.A(instr_sra),
    .B(instr_srai),
    .Y(_01811_));
 sky130_fd_sc_hd__o21a_1 _14887_ (.A1(_03400_),
    .A2(_01811_),
    .B1(_07224_),
    .X(_01812_));
 sky130_fd_sc_hd__xor2_1 _14888_ (.A(_05205_),
    .B(\decoded_imm[31] ),
    .X(_01813_));
 sky130_fd_sc_hd__nor3_1 _14889_ (.A(_07633_),
    .B(_07636_),
    .C(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__o21a_1 _14890_ (.A1(_07633_),
    .A2(_07636_),
    .B1(_01813_),
    .X(_01815_));
 sky130_fd_sc_hd__nor3_1 _14891_ (.A(_03631_),
    .B(_01814_),
    .C(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__a22o_1 _14892_ (.A1(_05174_),
    .A2(_07279_),
    .B1(_07274_),
    .B2(_05076_),
    .X(_01817_));
 sky130_fd_sc_hd__o2bb2a_1 _14893_ (.A1_N(\reg_pc[31] ),
    .A2_N(_07282_),
    .B1(_05200_),
    .B2(_03387_),
    .X(_01818_));
 sky130_fd_sc_hd__o2bb2a_1 _14894_ (.A1_N(_01817_),
    .A2_N(_07277_),
    .B1(_07284_),
    .B2(_01818_),
    .X(_01819_));
 sky130_fd_sc_hd__nand2_1 _14895_ (.A(_01812_),
    .B(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__o22a_1 _14896_ (.A1(_05205_),
    .A2(_01812_),
    .B1(_01816_),
    .B2(_01820_),
    .X(_01088_));
 sky130_fd_sc_hd__nor2_2 _14897_ (.A(_03196_),
    .B(net299),
    .Y(_01821_));
 sky130_fd_sc_hd__or2_2 _14898_ (.A(net224),
    .B(net257),
    .X(_01822_));
 sky130_fd_sc_hd__nand2_2 _14899_ (.A(_01821_),
    .B(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__clkbuf_4 _14900_ (.A(_01823_),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _14901_ (.A0(net214),
    .A1(net183),
    .S(_01824_),
    .X(_01825_));
 sky130_fd_sc_hd__clkbuf_1 _14902_ (.A(_01825_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _14903_ (.A0(net217),
    .A1(net186),
    .S(_01824_),
    .X(_01826_));
 sky130_fd_sc_hd__clkbuf_1 _14904_ (.A(_01826_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _14905_ (.A0(net218),
    .A1(net187),
    .S(_01824_),
    .X(_01827_));
 sky130_fd_sc_hd__clkbuf_1 _14906_ (.A(_01827_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _14907_ (.A0(net219),
    .A1(net188),
    .S(_01824_),
    .X(_01828_));
 sky130_fd_sc_hd__clkbuf_1 _14908_ (.A(_01828_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _14909_ (.A0(net220),
    .A1(net189),
    .S(_01824_),
    .X(_01829_));
 sky130_fd_sc_hd__clkbuf_1 _14910_ (.A(_01829_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _14911_ (.A0(net221),
    .A1(net190),
    .S(_01824_),
    .X(_01830_));
 sky130_fd_sc_hd__clkbuf_1 _14912_ (.A(_01830_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _14913_ (.A0(net222),
    .A1(net191),
    .S(_01824_),
    .X(_01831_));
 sky130_fd_sc_hd__clkbuf_1 _14914_ (.A(_01831_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _14915_ (.A0(net223),
    .A1(net192),
    .S(_01824_),
    .X(_01832_));
 sky130_fd_sc_hd__clkbuf_1 _14916_ (.A(_01832_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _14917_ (.A0(net194),
    .A1(net163),
    .S(_01824_),
    .X(_01833_));
 sky130_fd_sc_hd__clkbuf_1 _14918_ (.A(_01833_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _14919_ (.A0(net195),
    .A1(net164),
    .S(_01824_),
    .X(_01834_));
 sky130_fd_sc_hd__clkbuf_1 _14920_ (.A(_01834_),
    .X(_01098_));
 sky130_fd_sc_hd__clkbuf_4 _14921_ (.A(_01823_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _14922_ (.A0(net196),
    .A1(net165),
    .S(_01835_),
    .X(_01836_));
 sky130_fd_sc_hd__clkbuf_1 _14923_ (.A(_01836_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _14924_ (.A0(net197),
    .A1(net166),
    .S(_01835_),
    .X(_01837_));
 sky130_fd_sc_hd__clkbuf_1 _14925_ (.A(_01837_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _14926_ (.A0(net198),
    .A1(net167),
    .S(_01835_),
    .X(_01838_));
 sky130_fd_sc_hd__clkbuf_1 _14927_ (.A(_01838_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _14928_ (.A0(net199),
    .A1(net168),
    .S(_01835_),
    .X(_01839_));
 sky130_fd_sc_hd__clkbuf_1 _14929_ (.A(_01839_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _14930_ (.A0(net200),
    .A1(net169),
    .S(_01835_),
    .X(_01840_));
 sky130_fd_sc_hd__clkbuf_1 _14931_ (.A(_01840_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _14932_ (.A0(net201),
    .A1(net170),
    .S(_01835_),
    .X(_01841_));
 sky130_fd_sc_hd__clkbuf_1 _14933_ (.A(_01841_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _14934_ (.A0(net202),
    .A1(net171),
    .S(_01835_),
    .X(_01842_));
 sky130_fd_sc_hd__clkbuf_1 _14935_ (.A(_01842_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _14936_ (.A0(net203),
    .A1(net172),
    .S(_01835_),
    .X(_01843_));
 sky130_fd_sc_hd__clkbuf_1 _14937_ (.A(_01843_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _14938_ (.A0(net204),
    .A1(net173),
    .S(_01835_),
    .X(_01844_));
 sky130_fd_sc_hd__clkbuf_1 _14939_ (.A(_01844_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _14940_ (.A0(net205),
    .A1(net174),
    .S(_01835_),
    .X(_01845_));
 sky130_fd_sc_hd__clkbuf_1 _14941_ (.A(_01845_),
    .X(_01108_));
 sky130_fd_sc_hd__clkbuf_4 _14942_ (.A(_01823_),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_1 _14943_ (.A0(net206),
    .A1(net175),
    .S(_01846_),
    .X(_01847_));
 sky130_fd_sc_hd__clkbuf_1 _14944_ (.A(_01847_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _14945_ (.A0(net207),
    .A1(net176),
    .S(_01846_),
    .X(_01848_));
 sky130_fd_sc_hd__clkbuf_1 _14946_ (.A(_01848_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _14947_ (.A0(net208),
    .A1(net177),
    .S(_01846_),
    .X(_01849_));
 sky130_fd_sc_hd__clkbuf_1 _14948_ (.A(_01849_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _14949_ (.A0(net209),
    .A1(net178),
    .S(_01846_),
    .X(_01850_));
 sky130_fd_sc_hd__clkbuf_1 _14950_ (.A(_01850_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _14951_ (.A0(net210),
    .A1(net179),
    .S(_01846_),
    .X(_01851_));
 sky130_fd_sc_hd__clkbuf_1 _14952_ (.A(_01851_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _14953_ (.A0(net211),
    .A1(net180),
    .S(_01846_),
    .X(_01852_));
 sky130_fd_sc_hd__clkbuf_1 _14954_ (.A(_01852_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _14955_ (.A0(net212),
    .A1(net181),
    .S(_01846_),
    .X(_01853_));
 sky130_fd_sc_hd__clkbuf_1 _14956_ (.A(_01853_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _14957_ (.A0(net213),
    .A1(net182),
    .S(_01846_),
    .X(_01854_));
 sky130_fd_sc_hd__clkbuf_1 _14958_ (.A(_01854_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _14959_ (.A0(net215),
    .A1(net184),
    .S(_01846_),
    .X(_01855_));
 sky130_fd_sc_hd__clkbuf_1 _14960_ (.A(_01855_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _14961_ (.A0(net216),
    .A1(net185),
    .S(_01846_),
    .X(_01856_));
 sky130_fd_sc_hd__clkbuf_1 _14962_ (.A(_01856_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _14963_ (.A0(irq_delay),
    .A1(irq_active),
    .S(_07755_),
    .X(_01857_));
 sky130_fd_sc_hd__and2_1 _14964_ (.A(_07737_),
    .B(_01857_),
    .X(_01858_));
 sky130_fd_sc_hd__clkbuf_1 _14965_ (.A(_01858_),
    .X(_01119_));
 sky130_fd_sc_hd__nand2_1 _14966_ (.A(_06186_),
    .B(_03298_),
    .Y(_01859_));
 sky130_fd_sc_hd__a21o_1 _14967_ (.A1(_07679_),
    .A2(_01859_),
    .B1(_07680_),
    .X(_01860_));
 sky130_fd_sc_hd__o2bb2a_1 _14968_ (.A1_N(irq_active),
    .A2_N(_01860_),
    .B1(_01859_),
    .B2(_04150_),
    .X(_01861_));
 sky130_fd_sc_hd__nor2_1 _14969_ (.A(_08335_),
    .B(_01861_),
    .Y(_01120_));
 sky130_fd_sc_hd__nand2_1 _14970_ (.A(_03301_),
    .B(_04448_),
    .Y(_01862_));
 sky130_fd_sc_hd__clkbuf_4 _14971_ (.A(_01862_),
    .X(_01863_));
 sky130_fd_sc_hd__clkbuf_4 _14972_ (.A(_01863_),
    .X(_01864_));
 sky130_fd_sc_hd__clkbuf_4 _14973_ (.A(_01862_),
    .X(_01865_));
 sky130_fd_sc_hd__nor2_1 _14974_ (.A(_07208_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__a211o_1 _14975_ (.A1(\irq_mask[0] ),
    .A2(_01864_),
    .B1(_01866_),
    .C1(_08335_),
    .X(_01121_));
 sky130_fd_sc_hd__nor2_1 _14976_ (.A(_04101_),
    .B(_01865_),
    .Y(_01867_));
 sky130_fd_sc_hd__a211o_1 _14977_ (.A1(\irq_mask[1] ),
    .A2(_01864_),
    .B1(_01867_),
    .C1(_08335_),
    .X(_01122_));
 sky130_fd_sc_hd__nor2_1 _14978_ (.A(_04142_),
    .B(_01865_),
    .Y(_01868_));
 sky130_fd_sc_hd__a211o_1 _14979_ (.A1(\irq_mask[2] ),
    .A2(_01864_),
    .B1(_01868_),
    .C1(_08335_),
    .X(_01123_));
 sky130_fd_sc_hd__clkbuf_4 _14980_ (.A(_01862_),
    .X(_01869_));
 sky130_fd_sc_hd__nor2_1 _14981_ (.A(_04185_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__a211o_1 _14982_ (.A1(\irq_mask[3] ),
    .A2(_01864_),
    .B1(_01870_),
    .C1(_08335_),
    .X(_01124_));
 sky130_fd_sc_hd__nor2_1 _14983_ (.A(_04240_),
    .B(_01869_),
    .Y(_01871_));
 sky130_fd_sc_hd__a211o_1 _14984_ (.A1(\irq_mask[4] ),
    .A2(_01864_),
    .B1(_01871_),
    .C1(_08335_),
    .X(_01125_));
 sky130_fd_sc_hd__or3_4 _14985_ (.A(_04227_),
    .B(_04298_),
    .C(_04306_),
    .X(_01872_));
 sky130_fd_sc_hd__nor2_1 _14986_ (.A(_01872_),
    .B(_01869_),
    .Y(_01873_));
 sky130_fd_sc_hd__a211o_1 _14987_ (.A1(\irq_mask[5] ),
    .A2(_01864_),
    .B1(_01873_),
    .C1(_08335_),
    .X(_01126_));
 sky130_fd_sc_hd__nor2_1 _14988_ (.A(_04335_),
    .B(_01869_),
    .Y(_01874_));
 sky130_fd_sc_hd__a211o_1 _14989_ (.A1(\irq_mask[6] ),
    .A2(_01864_),
    .B1(_01874_),
    .C1(_08335_),
    .X(_01127_));
 sky130_fd_sc_hd__nor2_1 _14990_ (.A(_04382_),
    .B(_01869_),
    .Y(_01875_));
 sky130_fd_sc_hd__clkbuf_4 _14991_ (.A(_03240_),
    .X(_01876_));
 sky130_fd_sc_hd__a211o_1 _14992_ (.A1(\irq_mask[7] ),
    .A2(_01864_),
    .B1(_01875_),
    .C1(_01876_),
    .X(_01128_));
 sky130_fd_sc_hd__nor2_1 _14993_ (.A(_04414_),
    .B(_01869_),
    .Y(_01877_));
 sky130_fd_sc_hd__a211o_1 _14994_ (.A1(\irq_mask[8] ),
    .A2(_01864_),
    .B1(_01877_),
    .C1(_01876_),
    .X(_01129_));
 sky130_fd_sc_hd__a21o_1 _14995_ (.A1(\irq_mask[9] ),
    .A2(_01863_),
    .B1(_01714_),
    .X(_01878_));
 sky130_fd_sc_hd__a31o_1 _14996_ (.A1(_03303_),
    .A2(_04022_),
    .A3(_04447_),
    .B1(_01878_),
    .X(_01130_));
 sky130_fd_sc_hd__nor2_1 _14997_ (.A(_04493_),
    .B(_01869_),
    .Y(_01879_));
 sky130_fd_sc_hd__a211o_1 _14998_ (.A1(\irq_mask[10] ),
    .A2(_01864_),
    .B1(_01879_),
    .C1(_01876_),
    .X(_01131_));
 sky130_fd_sc_hd__clkbuf_4 _14999_ (.A(_01862_),
    .X(_01880_));
 sky130_fd_sc_hd__or3_4 _15000_ (.A(_04227_),
    .B(_04517_),
    .C(_04525_),
    .X(_01881_));
 sky130_fd_sc_hd__nor2_1 _15001_ (.A(_01881_),
    .B(_01869_),
    .Y(_01882_));
 sky130_fd_sc_hd__a211o_1 _15002_ (.A1(\irq_mask[11] ),
    .A2(_01880_),
    .B1(_01882_),
    .C1(_01876_),
    .X(_01132_));
 sky130_fd_sc_hd__nor2_1 _15003_ (.A(_04561_),
    .B(_01869_),
    .Y(_01883_));
 sky130_fd_sc_hd__a211o_1 _15004_ (.A1(\irq_mask[12] ),
    .A2(_01880_),
    .B1(_01883_),
    .C1(_01876_),
    .X(_01133_));
 sky130_fd_sc_hd__nor2_1 _15005_ (.A(_04592_),
    .B(_01869_),
    .Y(_01884_));
 sky130_fd_sc_hd__a211o_1 _15006_ (.A1(\irq_mask[13] ),
    .A2(_01880_),
    .B1(_01884_),
    .C1(_01876_),
    .X(_01134_));
 sky130_fd_sc_hd__clkbuf_4 _15007_ (.A(_01862_),
    .X(_01885_));
 sky130_fd_sc_hd__nor2_1 _15008_ (.A(_04631_),
    .B(_01885_),
    .Y(_01886_));
 sky130_fd_sc_hd__a211o_1 _15009_ (.A1(\irq_mask[14] ),
    .A2(_01880_),
    .B1(_01886_),
    .C1(_01876_),
    .X(_01135_));
 sky130_fd_sc_hd__nor2_1 _15010_ (.A(_04659_),
    .B(_01885_),
    .Y(_01887_));
 sky130_fd_sc_hd__a211o_1 _15011_ (.A1(\irq_mask[15] ),
    .A2(_01880_),
    .B1(_01887_),
    .C1(_01876_),
    .X(_01136_));
 sky130_fd_sc_hd__nor2_1 _15012_ (.A(_04702_),
    .B(_01885_),
    .Y(_01888_));
 sky130_fd_sc_hd__a211o_1 _15013_ (.A1(\irq_mask[16] ),
    .A2(_01880_),
    .B1(_01888_),
    .C1(_01876_),
    .X(_01137_));
 sky130_fd_sc_hd__nor2_1 _15014_ (.A(_04737_),
    .B(_01885_),
    .Y(_01889_));
 sky130_fd_sc_hd__a211o_1 _15015_ (.A1(\irq_mask[17] ),
    .A2(_01880_),
    .B1(_01889_),
    .C1(_01876_),
    .X(_01138_));
 sky130_fd_sc_hd__nor2_1 _15016_ (.A(_04776_),
    .B(_01885_),
    .Y(_01890_));
 sky130_fd_sc_hd__clkbuf_4 _15017_ (.A(_03240_),
    .X(_01891_));
 sky130_fd_sc_hd__a211o_1 _15018_ (.A1(\irq_mask[18] ),
    .A2(_01880_),
    .B1(_01890_),
    .C1(_01891_),
    .X(_01139_));
 sky130_fd_sc_hd__nor2_1 _15019_ (.A(_04805_),
    .B(_01885_),
    .Y(_01892_));
 sky130_fd_sc_hd__a211o_1 _15020_ (.A1(\irq_mask[19] ),
    .A2(_01880_),
    .B1(_01892_),
    .C1(_01891_),
    .X(_01140_));
 sky130_fd_sc_hd__a21o_1 _15021_ (.A1(\irq_mask[20] ),
    .A2(_01863_),
    .B1(_01714_),
    .X(_01893_));
 sky130_fd_sc_hd__a31o_1 _15022_ (.A1(_03303_),
    .A2(_04022_),
    .A3(_04842_),
    .B1(_01893_),
    .X(_01141_));
 sky130_fd_sc_hd__a21o_1 _15023_ (.A1(\irq_mask[21] ),
    .A2(_01863_),
    .B1(_01714_),
    .X(_01894_));
 sky130_fd_sc_hd__a31o_1 _15024_ (.A1(_03303_),
    .A2(_04022_),
    .A3(_04871_),
    .B1(_01894_),
    .X(_01142_));
 sky130_fd_sc_hd__nor2_1 _15025_ (.A(_04908_),
    .B(_01885_),
    .Y(_01895_));
 sky130_fd_sc_hd__a211o_1 _15026_ (.A1(\irq_mask[22] ),
    .A2(_01880_),
    .B1(_01895_),
    .C1(_01891_),
    .X(_01143_));
 sky130_fd_sc_hd__nor2_1 _15027_ (.A(_04940_),
    .B(_01885_),
    .Y(_01896_));
 sky130_fd_sc_hd__a211o_1 _15028_ (.A1(\irq_mask[23] ),
    .A2(_01865_),
    .B1(_01896_),
    .C1(_01891_),
    .X(_01144_));
 sky130_fd_sc_hd__a21o_1 _15029_ (.A1(\irq_mask[24] ),
    .A2(_01863_),
    .B1(_01714_),
    .X(_01897_));
 sky130_fd_sc_hd__a31o_1 _15030_ (.A1(_03303_),
    .A2(_04022_),
    .A3(_04979_),
    .B1(_01897_),
    .X(_01145_));
 sky130_fd_sc_hd__a21o_1 _15031_ (.A1(\irq_mask[25] ),
    .A2(_01863_),
    .B1(_03240_),
    .X(_01898_));
 sky130_fd_sc_hd__a31o_1 _15032_ (.A1(_03303_),
    .A2(_04022_),
    .A3(_05009_),
    .B1(_01898_),
    .X(_01146_));
 sky130_fd_sc_hd__nor2_1 _15033_ (.A(_05037_),
    .B(_01885_),
    .Y(_01899_));
 sky130_fd_sc_hd__a211o_1 _15034_ (.A1(\irq_mask[26] ),
    .A2(_01865_),
    .B1(_01899_),
    .C1(_01891_),
    .X(_01147_));
 sky130_fd_sc_hd__nor2_1 _15035_ (.A(_05069_),
    .B(_01885_),
    .Y(_01900_));
 sky130_fd_sc_hd__a211o_1 _15036_ (.A1(\irq_mask[27] ),
    .A2(_01865_),
    .B1(_01900_),
    .C1(_01891_),
    .X(_01148_));
 sky130_fd_sc_hd__nor2_1 _15037_ (.A(_05106_),
    .B(_01863_),
    .Y(_01901_));
 sky130_fd_sc_hd__a211o_1 _15038_ (.A1(\irq_mask[28] ),
    .A2(_01865_),
    .B1(_01901_),
    .C1(_01891_),
    .X(_01149_));
 sky130_fd_sc_hd__nor2_1 _15039_ (.A(_05138_),
    .B(_01863_),
    .Y(_01902_));
 sky130_fd_sc_hd__a211o_1 _15040_ (.A1(\irq_mask[29] ),
    .A2(_01865_),
    .B1(_01902_),
    .C1(_01891_),
    .X(_01150_));
 sky130_fd_sc_hd__nor2_1 _15041_ (.A(_05169_),
    .B(_01863_),
    .Y(_01903_));
 sky130_fd_sc_hd__a211o_1 _15042_ (.A1(\irq_mask[30] ),
    .A2(_01865_),
    .B1(_01903_),
    .C1(_01891_),
    .X(_01151_));
 sky130_fd_sc_hd__nor2_1 _15043_ (.A(_05200_),
    .B(_01863_),
    .Y(_01904_));
 sky130_fd_sc_hd__a211o_1 _15044_ (.A1(\irq_mask[31] ),
    .A2(_01865_),
    .B1(_01904_),
    .C1(_01891_),
    .X(_01152_));
 sky130_fd_sc_hd__buf_4 _15045_ (.A(_03272_),
    .X(_01905_));
 sky130_fd_sc_hd__buf_4 _15046_ (.A(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__buf_8 _15047_ (.A(_03664_),
    .X(_01907_));
 sky130_fd_sc_hd__buf_6 _15048_ (.A(_03670_),
    .X(_01908_));
 sky130_fd_sc_hd__buf_6 _15049_ (.A(_03671_),
    .X(_01909_));
 sky130_fd_sc_hd__mux4_1 _15050_ (.A0(\cpuregs.regs[12][0] ),
    .A1(\cpuregs.regs[13][0] ),
    .A2(\cpuregs.regs[14][0] ),
    .A3(\cpuregs.regs[15][0] ),
    .S0(_01908_),
    .S1(_01909_),
    .X(_01910_));
 sky130_fd_sc_hd__mux4_1 _15051_ (.A0(\cpuregs.regs[8][0] ),
    .A1(\cpuregs.regs[9][0] ),
    .A2(\cpuregs.regs[10][0] ),
    .A3(\cpuregs.regs[11][0] ),
    .S0(_03658_),
    .S1(_03659_),
    .X(_01911_));
 sky130_fd_sc_hd__or2_1 _15052_ (.A(_03666_),
    .B(_01911_),
    .X(_01912_));
 sky130_fd_sc_hd__o211a_1 _15053_ (.A1(_01907_),
    .A2(_01910_),
    .B1(_01912_),
    .C1(_03654_),
    .X(_01913_));
 sky130_fd_sc_hd__mux4_1 _15054_ (.A0(\cpuregs.regs[4][0] ),
    .A1(\cpuregs.regs[5][0] ),
    .A2(\cpuregs.regs[6][0] ),
    .A3(\cpuregs.regs[7][0] ),
    .S0(_03658_),
    .S1(_03659_),
    .X(_01914_));
 sky130_fd_sc_hd__mux4_1 _15055_ (.A0(\cpuregs.regs[0][0] ),
    .A1(\cpuregs.regs[1][0] ),
    .A2(\cpuregs.regs[2][0] ),
    .A3(\cpuregs.regs[3][0] ),
    .S0(_03658_),
    .S1(_03659_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _15056_ (.A0(_01914_),
    .A1(_01915_),
    .S(_03664_),
    .X(_01916_));
 sky130_fd_sc_hd__a21o_1 _15057_ (.A1(_03657_),
    .A2(_01916_),
    .B1(_03692_),
    .X(_01917_));
 sky130_fd_sc_hd__buf_8 _15058_ (.A(_03670_),
    .X(_01918_));
 sky130_fd_sc_hd__buf_6 _15059_ (.A(_03671_),
    .X(_01919_));
 sky130_fd_sc_hd__mux4_1 _15060_ (.A0(\cpuregs.regs[28][0] ),
    .A1(\cpuregs.regs[29][0] ),
    .A2(\cpuregs.regs[30][0] ),
    .A3(\cpuregs.regs[31][0] ),
    .S0(_01918_),
    .S1(_01919_),
    .X(_01920_));
 sky130_fd_sc_hd__mux4_1 _15061_ (.A0(\cpuregs.regs[24][0] ),
    .A1(\cpuregs.regs[25][0] ),
    .A2(\cpuregs.regs[26][0] ),
    .A3(\cpuregs.regs[27][0] ),
    .S0(_03670_),
    .S1(_03671_),
    .X(_01921_));
 sky130_fd_sc_hd__or2_1 _15062_ (.A(_03666_),
    .B(_01921_),
    .X(_01922_));
 sky130_fd_sc_hd__o211a_1 _15063_ (.A1(_01907_),
    .A2(_01920_),
    .B1(_01922_),
    .C1(_03654_),
    .X(_01923_));
 sky130_fd_sc_hd__mux4_1 _15064_ (.A0(\cpuregs.regs[20][0] ),
    .A1(\cpuregs.regs[21][0] ),
    .A2(\cpuregs.regs[22][0] ),
    .A3(\cpuregs.regs[23][0] ),
    .S0(_03670_),
    .S1(_03671_),
    .X(_01924_));
 sky130_fd_sc_hd__mux4_1 _15065_ (.A0(\cpuregs.regs[16][0] ),
    .A1(\cpuregs.regs[17][0] ),
    .A2(\cpuregs.regs[18][0] ),
    .A3(\cpuregs.regs[19][0] ),
    .S0(_03670_),
    .S1(_03671_),
    .X(_01925_));
 sky130_fd_sc_hd__mux2_1 _15066_ (.A0(_01924_),
    .A1(_01925_),
    .S(_03664_),
    .X(_01926_));
 sky130_fd_sc_hd__a21o_1 _15067_ (.A1(_03657_),
    .A2(_01926_),
    .B1(_03675_),
    .X(_01927_));
 sky130_fd_sc_hd__o22a_1 _15068_ (.A1(_01913_),
    .A2(_01917_),
    .B1(_01923_),
    .B2(_01927_),
    .X(_01928_));
 sky130_fd_sc_hd__nand2_2 _15069_ (.A(_03679_),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__nor2_1 _15070_ (.A(_03388_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__inv_2 _15071_ (.A(is_slli_srli_srai),
    .Y(_01931_));
 sky130_fd_sc_hd__a21o_2 _15072_ (.A1(_01931_),
    .A2(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B1(_03387_),
    .X(_01932_));
 sky130_fd_sc_hd__buf_4 _15073_ (.A(_01932_),
    .X(_01933_));
 sky130_fd_sc_hd__nand2_4 _15074_ (.A(_03277_),
    .B(_03301_),
    .Y(_01934_));
 sky130_fd_sc_hd__a221o_1 _15075_ (.A1(is_slli_srli_srai),
    .A2(\cpuregs.raddr2[0] ),
    .B1(\decoded_imm[0] ),
    .B2(_01933_),
    .C1(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__o22a_1 _15076_ (.A1(_05324_),
    .A2(_01906_),
    .B1(_01930_),
    .B2(_01935_),
    .X(_01153_));
 sky130_fd_sc_hd__buf_6 _15077_ (.A(_03669_),
    .X(_01936_));
 sky130_fd_sc_hd__clkbuf_8 _15078_ (.A(_03646_),
    .X(_01937_));
 sky130_fd_sc_hd__mux4_1 _15079_ (.A0(\cpuregs.regs[8][1] ),
    .A1(\cpuregs.regs[9][1] ),
    .A2(\cpuregs.regs[10][1] ),
    .A3(\cpuregs.regs[11][1] ),
    .S0(_01936_),
    .S1(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__mux4_1 _15080_ (.A0(\cpuregs.regs[12][1] ),
    .A1(\cpuregs.regs[13][1] ),
    .A2(\cpuregs.regs[14][1] ),
    .A3(\cpuregs.regs[15][1] ),
    .S0(_03669_),
    .S1(_03646_),
    .X(_01939_));
 sky130_fd_sc_hd__or2_1 _15081_ (.A(_03713_),
    .B(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__o211a_1 _15082_ (.A1(_03709_),
    .A2(_01938_),
    .B1(_01940_),
    .C1(_00067_),
    .X(_01941_));
 sky130_fd_sc_hd__mux4_1 _15083_ (.A0(\cpuregs.regs[4][1] ),
    .A1(\cpuregs.regs[5][1] ),
    .A2(\cpuregs.regs[6][1] ),
    .A3(\cpuregs.regs[7][1] ),
    .S0(_03669_),
    .S1(_03646_),
    .X(_01942_));
 sky130_fd_sc_hd__mux4_1 _15084_ (.A0(\cpuregs.regs[0][1] ),
    .A1(\cpuregs.regs[1][1] ),
    .A2(\cpuregs.regs[2][1] ),
    .A3(\cpuregs.regs[3][1] ),
    .S0(_03669_),
    .S1(_03646_),
    .X(_01943_));
 sky130_fd_sc_hd__mux2_1 _15085_ (.A0(_01942_),
    .A1(_01943_),
    .S(_03713_),
    .X(_01944_));
 sky130_fd_sc_hd__a21o_1 _15086_ (.A1(_03656_),
    .A2(_01944_),
    .B1(_00068_),
    .X(_01945_));
 sky130_fd_sc_hd__mux4_1 _15087_ (.A0(\cpuregs.regs[28][1] ),
    .A1(\cpuregs.regs[29][1] ),
    .A2(\cpuregs.regs[30][1] ),
    .A3(\cpuregs.regs[31][1] ),
    .S0(_01936_),
    .S1(_03647_),
    .X(_01946_));
 sky130_fd_sc_hd__mux4_1 _15088_ (.A0(\cpuregs.regs[24][1] ),
    .A1(\cpuregs.regs[25][1] ),
    .A2(\cpuregs.regs[26][1] ),
    .A3(\cpuregs.regs[27][1] ),
    .S0(_03669_),
    .S1(_03646_),
    .X(_01947_));
 sky130_fd_sc_hd__or2_1 _15089_ (.A(_03666_),
    .B(_01947_),
    .X(_01948_));
 sky130_fd_sc_hd__o211a_1 _15090_ (.A1(_03719_),
    .A2(_01946_),
    .B1(_01948_),
    .C1(_00067_),
    .X(_01949_));
 sky130_fd_sc_hd__mux4_1 _15091_ (.A0(\cpuregs.regs[20][1] ),
    .A1(\cpuregs.regs[21][1] ),
    .A2(\cpuregs.regs[22][1] ),
    .A3(\cpuregs.regs[23][1] ),
    .S0(_03669_),
    .S1(_03646_),
    .X(_01950_));
 sky130_fd_sc_hd__mux4_1 _15092_ (.A0(\cpuregs.regs[16][1] ),
    .A1(\cpuregs.regs[17][1] ),
    .A2(\cpuregs.regs[18][1] ),
    .A3(\cpuregs.regs[19][1] ),
    .S0(_03669_),
    .S1(_03646_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _15093_ (.A0(_01950_),
    .A1(_01951_),
    .S(_03713_),
    .X(_01952_));
 sky130_fd_sc_hd__a21o_1 _15094_ (.A1(_03656_),
    .A2(_01952_),
    .B1(_03674_),
    .X(_01953_));
 sky130_fd_sc_hd__o22a_2 _15095_ (.A1(_01941_),
    .A2(_01945_),
    .B1(_01949_),
    .B2(_01953_),
    .X(_01954_));
 sky130_fd_sc_hd__nand2_2 _15096_ (.A(_03679_),
    .B(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__nor2_1 _15097_ (.A(_03388_),
    .B(_01955_),
    .Y(_01956_));
 sky130_fd_sc_hd__a221o_1 _15098_ (.A1(is_slli_srli_srai),
    .A2(\cpuregs.raddr2[1] ),
    .B1(\decoded_imm[1] ),
    .B2(_01933_),
    .C1(_01934_),
    .X(_01957_));
 sky130_fd_sc_hd__o22a_1 _15099_ (.A1(_05286_),
    .A2(_01906_),
    .B1(_01956_),
    .B2(_01957_),
    .X(_01154_));
 sky130_fd_sc_hd__and2_1 _15100_ (.A(_03396_),
    .B(_03679_),
    .X(_01958_));
 sky130_fd_sc_hd__buf_4 _15101_ (.A(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__buf_8 _15102_ (.A(_01959_),
    .X(_01960_));
 sky130_fd_sc_hd__a221o_1 _15103_ (.A1(is_slli_srli_srai),
    .A2(\cpuregs.raddr2[2] ),
    .B1(\decoded_imm[2] ),
    .B2(_01932_),
    .C1(_01934_),
    .X(_01961_));
 sky130_fd_sc_hd__a21o_1 _15104_ (.A1(_03677_),
    .A2(_01960_),
    .B1(_01961_),
    .X(_01962_));
 sky130_fd_sc_hd__o21a_1 _15105_ (.A1(_05413_),
    .A2(_01906_),
    .B1(_01962_),
    .X(_01155_));
 sky130_fd_sc_hd__buf_6 _15106_ (.A(_01934_),
    .X(_01963_));
 sky130_fd_sc_hd__a221o_1 _15107_ (.A1(is_slli_srli_srai),
    .A2(\cpuregs.raddr2[3] ),
    .B1(\decoded_imm[3] ),
    .B2(_01933_),
    .C1(_01934_),
    .X(_01964_));
 sky130_fd_sc_hd__a21oi_2 _15108_ (.A1(_03396_),
    .A2(_03703_),
    .B1(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__a21oi_1 _15109_ (.A1(_05288_),
    .A2(_01963_),
    .B1(_01965_),
    .Y(_01156_));
 sky130_fd_sc_hd__a221o_1 _15110_ (.A1(is_slli_srli_srai),
    .A2(\cpuregs.raddr2[4] ),
    .B1(\decoded_imm[4] ),
    .B2(_01932_),
    .C1(_01934_),
    .X(_01966_));
 sky130_fd_sc_hd__a21o_1 _15111_ (.A1(_03396_),
    .A2(_03726_),
    .B1(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__o21a_1 _15112_ (.A1(_05255_),
    .A2(_01906_),
    .B1(_01967_),
    .X(_01157_));
 sky130_fd_sc_hd__buf_8 _15113_ (.A(_03654_),
    .X(_01968_));
 sky130_fd_sc_hd__buf_8 _15114_ (.A(_01968_),
    .X(_01969_));
 sky130_fd_sc_hd__buf_8 _15115_ (.A(_01918_),
    .X(_01970_));
 sky130_fd_sc_hd__buf_8 _15116_ (.A(_01919_),
    .X(_01971_));
 sky130_fd_sc_hd__mux4_1 _15117_ (.A0(\cpuregs.regs[4][5] ),
    .A1(\cpuregs.regs[5][5] ),
    .A2(\cpuregs.regs[6][5] ),
    .A3(\cpuregs.regs[7][5] ),
    .S0(_01970_),
    .S1(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__clkbuf_16 _15118_ (.A(_01918_),
    .X(_01973_));
 sky130_fd_sc_hd__buf_8 _15119_ (.A(_01919_),
    .X(_01974_));
 sky130_fd_sc_hd__mux4_1 _15120_ (.A0(\cpuregs.regs[0][5] ),
    .A1(\cpuregs.regs[1][5] ),
    .A2(\cpuregs.regs[2][5] ),
    .A3(\cpuregs.regs[3][5] ),
    .S0(_01973_),
    .S1(_01974_),
    .X(_01975_));
 sky130_fd_sc_hd__buf_8 _15121_ (.A(_01918_),
    .X(_01976_));
 sky130_fd_sc_hd__buf_6 _15122_ (.A(_01919_),
    .X(_01977_));
 sky130_fd_sc_hd__mux4_1 _15123_ (.A0(\cpuregs.regs[20][5] ),
    .A1(\cpuregs.regs[21][5] ),
    .A2(\cpuregs.regs[22][5] ),
    .A3(\cpuregs.regs[23][5] ),
    .S0(_01976_),
    .S1(_01977_),
    .X(_01978_));
 sky130_fd_sc_hd__clkbuf_16 _15124_ (.A(_01918_),
    .X(_01979_));
 sky130_fd_sc_hd__buf_8 _15125_ (.A(_01919_),
    .X(_01980_));
 sky130_fd_sc_hd__mux4_1 _15126_ (.A0(\cpuregs.regs[16][5] ),
    .A1(\cpuregs.regs[17][5] ),
    .A2(\cpuregs.regs[18][5] ),
    .A3(\cpuregs.regs[19][5] ),
    .S0(_01979_),
    .S1(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__buf_8 _15127_ (.A(_01907_),
    .X(_01982_));
 sky130_fd_sc_hd__mux4_1 _15128_ (.A0(_01972_),
    .A1(_01975_),
    .A2(_01978_),
    .A3(_01981_),
    .S0(_01982_),
    .S1(_03639_),
    .X(_01983_));
 sky130_fd_sc_hd__buf_8 _15129_ (.A(_03719_),
    .X(_01984_));
 sky130_fd_sc_hd__buf_8 _15130_ (.A(_01936_),
    .X(_01985_));
 sky130_fd_sc_hd__buf_6 _15131_ (.A(_03647_),
    .X(_01986_));
 sky130_fd_sc_hd__mux4_1 _15132_ (.A0(\cpuregs.regs[28][5] ),
    .A1(\cpuregs.regs[29][5] ),
    .A2(\cpuregs.regs[30][5] ),
    .A3(\cpuregs.regs[31][5] ),
    .S0(_01985_),
    .S1(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__or2_1 _15133_ (.A(_01984_),
    .B(_01987_),
    .X(_01988_));
 sky130_fd_sc_hd__buf_4 _15134_ (.A(_03666_),
    .X(_01989_));
 sky130_fd_sc_hd__buf_8 _15135_ (.A(_01936_),
    .X(_01990_));
 sky130_fd_sc_hd__buf_6 _15136_ (.A(_03642_),
    .X(_01991_));
 sky130_fd_sc_hd__buf_8 _15137_ (.A(_01991_),
    .X(_01992_));
 sky130_fd_sc_hd__mux4_1 _15138_ (.A0(\cpuregs.regs[24][5] ),
    .A1(\cpuregs.regs[25][5] ),
    .A2(\cpuregs.regs[26][5] ),
    .A3(\cpuregs.regs[27][5] ),
    .S0(_01990_),
    .S1(_01992_),
    .X(_01993_));
 sky130_fd_sc_hd__o21a_1 _15139_ (.A1(_01989_),
    .A2(_01993_),
    .B1(_03692_),
    .X(_01994_));
 sky130_fd_sc_hd__buf_6 _15140_ (.A(_03669_),
    .X(_01995_));
 sky130_fd_sc_hd__buf_8 _15141_ (.A(_01995_),
    .X(_01996_));
 sky130_fd_sc_hd__buf_8 _15142_ (.A(_03647_),
    .X(_01997_));
 sky130_fd_sc_hd__mux4_1 _15143_ (.A0(\cpuregs.regs[12][5] ),
    .A1(\cpuregs.regs[13][5] ),
    .A2(\cpuregs.regs[14][5] ),
    .A3(\cpuregs.regs[15][5] ),
    .S0(_01996_),
    .S1(_01997_),
    .X(_01998_));
 sky130_fd_sc_hd__buf_8 _15144_ (.A(_01995_),
    .X(_01999_));
 sky130_fd_sc_hd__buf_8 _15145_ (.A(_03647_),
    .X(_02000_));
 sky130_fd_sc_hd__mux4_1 _15146_ (.A0(\cpuregs.regs[8][5] ),
    .A1(\cpuregs.regs[9][5] ),
    .A2(\cpuregs.regs[10][5] ),
    .A3(\cpuregs.regs[11][5] ),
    .S0(_01999_),
    .S1(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__buf_8 _15147_ (.A(_03653_),
    .X(_02002_));
 sky130_fd_sc_hd__mux2_1 _15148_ (.A0(_01998_),
    .A1(_02001_),
    .S(_02002_),
    .X(_02003_));
 sky130_fd_sc_hd__buf_6 _15149_ (.A(_03675_),
    .X(_02004_));
 sky130_fd_sc_hd__clkbuf_8 _15150_ (.A(_03656_),
    .X(_02005_));
 sky130_fd_sc_hd__clkbuf_8 _15151_ (.A(_02005_),
    .X(_02006_));
 sky130_fd_sc_hd__a221o_1 _15152_ (.A1(_01988_),
    .A2(_01994_),
    .B1(_02003_),
    .B2(_02004_),
    .C1(_02006_),
    .X(_02007_));
 sky130_fd_sc_hd__o211a_1 _15153_ (.A1(_01969_),
    .A2(_01983_),
    .B1(_02007_),
    .C1(_01960_),
    .X(_02008_));
 sky130_fd_sc_hd__buf_4 _15154_ (.A(_01933_),
    .X(_02009_));
 sky130_fd_sc_hd__a21o_1 _15155_ (.A1(\decoded_imm[5] ),
    .A2(_02009_),
    .B1(_01963_),
    .X(_02010_));
 sky130_fd_sc_hd__o22a_1 _15156_ (.A1(net126),
    .A2(_01906_),
    .B1(_02008_),
    .B2(_02010_),
    .X(_01158_));
 sky130_fd_sc_hd__mux4_1 _15157_ (.A0(\cpuregs.regs[8][6] ),
    .A1(\cpuregs.regs[9][6] ),
    .A2(\cpuregs.regs[10][6] ),
    .A3(\cpuregs.regs[11][6] ),
    .S0(_01970_),
    .S1(_01971_),
    .X(_02011_));
 sky130_fd_sc_hd__buf_6 _15158_ (.A(_03653_),
    .X(_02012_));
 sky130_fd_sc_hd__buf_8 _15159_ (.A(_01936_),
    .X(_02013_));
 sky130_fd_sc_hd__clkbuf_8 _15160_ (.A(_03643_),
    .X(_02014_));
 sky130_fd_sc_hd__mux4_1 _15161_ (.A0(\cpuregs.regs[12][6] ),
    .A1(\cpuregs.regs[13][6] ),
    .A2(\cpuregs.regs[14][6] ),
    .A3(\cpuregs.regs[15][6] ),
    .S0(_02013_),
    .S1(_02014_),
    .X(_02015_));
 sky130_fd_sc_hd__or2_1 _15162_ (.A(_02012_),
    .B(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__buf_6 _15163_ (.A(_03674_),
    .X(_02017_));
 sky130_fd_sc_hd__clkbuf_8 _15164_ (.A(_02017_),
    .X(_02018_));
 sky130_fd_sc_hd__o211a_1 _15165_ (.A1(_01989_),
    .A2(_02011_),
    .B1(_02016_),
    .C1(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__buf_6 _15166_ (.A(_03639_),
    .X(_02020_));
 sky130_fd_sc_hd__mux4_1 _15167_ (.A0(\cpuregs.regs[28][6] ),
    .A1(\cpuregs.regs[29][6] ),
    .A2(\cpuregs.regs[30][6] ),
    .A3(\cpuregs.regs[31][6] ),
    .S0(_01990_),
    .S1(_01992_),
    .X(_02021_));
 sky130_fd_sc_hd__buf_6 _15168_ (.A(_01936_),
    .X(_02022_));
 sky130_fd_sc_hd__clkbuf_8 _15169_ (.A(_03647_),
    .X(_02023_));
 sky130_fd_sc_hd__mux4_1 _15170_ (.A0(\cpuregs.regs[24][6] ),
    .A1(\cpuregs.regs[25][6] ),
    .A2(\cpuregs.regs[26][6] ),
    .A3(\cpuregs.regs[27][6] ),
    .S0(_02022_),
    .S1(_02023_),
    .X(_02024_));
 sky130_fd_sc_hd__mux2_1 _15171_ (.A0(_02021_),
    .A1(_02024_),
    .S(_01984_),
    .X(_02025_));
 sky130_fd_sc_hd__a21o_1 _15172_ (.A1(_02020_),
    .A2(_02025_),
    .B1(_02006_),
    .X(_02026_));
 sky130_fd_sc_hd__buf_8 _15173_ (.A(_01959_),
    .X(_02027_));
 sky130_fd_sc_hd__mux4_1 _15174_ (.A0(\cpuregs.regs[4][6] ),
    .A1(\cpuregs.regs[5][6] ),
    .A2(\cpuregs.regs[6][6] ),
    .A3(\cpuregs.regs[7][6] ),
    .S0(_02013_),
    .S1(_02014_),
    .X(_02028_));
 sky130_fd_sc_hd__or2_1 _15175_ (.A(_02012_),
    .B(_02028_),
    .X(_02029_));
 sky130_fd_sc_hd__buf_6 _15176_ (.A(_03649_),
    .X(_02030_));
 sky130_fd_sc_hd__buf_6 _15177_ (.A(_03684_),
    .X(_02031_));
 sky130_fd_sc_hd__mux4_1 _15178_ (.A0(\cpuregs.regs[0][6] ),
    .A1(\cpuregs.regs[1][6] ),
    .A2(\cpuregs.regs[2][6] ),
    .A3(\cpuregs.regs[3][6] ),
    .S0(_02030_),
    .S1(_02031_),
    .X(_02032_));
 sky130_fd_sc_hd__o21a_1 _15179_ (.A1(_01989_),
    .A2(_02032_),
    .B1(_02017_),
    .X(_02033_));
 sky130_fd_sc_hd__mux4_1 _15180_ (.A0(\cpuregs.regs[20][6] ),
    .A1(\cpuregs.regs[21][6] ),
    .A2(\cpuregs.regs[22][6] ),
    .A3(\cpuregs.regs[23][6] ),
    .S0(_02022_),
    .S1(_02023_),
    .X(_02034_));
 sky130_fd_sc_hd__mux4_1 _15181_ (.A0(\cpuregs.regs[16][6] ),
    .A1(\cpuregs.regs[17][6] ),
    .A2(\cpuregs.regs[18][6] ),
    .A3(\cpuregs.regs[19][6] ),
    .S0(_01985_),
    .S1(_01986_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _15182_ (.A0(_02034_),
    .A1(_02035_),
    .S(_02002_),
    .X(_02036_));
 sky130_fd_sc_hd__clkbuf_8 _15183_ (.A(_03692_),
    .X(_02037_));
 sky130_fd_sc_hd__a221o_1 _15184_ (.A1(_02029_),
    .A2(_02033_),
    .B1(_02036_),
    .B2(_02037_),
    .C1(_01969_),
    .X(_02038_));
 sky130_fd_sc_hd__o211a_2 _15185_ (.A1(_02019_),
    .A2(_02026_),
    .B1(_02027_),
    .C1(_02038_),
    .X(_02039_));
 sky130_fd_sc_hd__a21o_1 _15186_ (.A1(\decoded_imm[6] ),
    .A2(_02009_),
    .B1(_01963_),
    .X(_02040_));
 sky130_fd_sc_hd__o22a_1 _15187_ (.A1(net127),
    .A2(_01906_),
    .B1(_02039_),
    .B2(_02040_),
    .X(_01159_));
 sky130_fd_sc_hd__mux4_1 _15188_ (.A0(\cpuregs.regs[4][7] ),
    .A1(\cpuregs.regs[5][7] ),
    .A2(\cpuregs.regs[6][7] ),
    .A3(\cpuregs.regs[7][7] ),
    .S0(_03670_),
    .S1(_03671_),
    .X(_02041_));
 sky130_fd_sc_hd__mux4_1 _15189_ (.A0(\cpuregs.regs[0][7] ),
    .A1(\cpuregs.regs[1][7] ),
    .A2(\cpuregs.regs[2][7] ),
    .A3(\cpuregs.regs[3][7] ),
    .S0(_03670_),
    .S1(_03671_),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_1 _15190_ (.A0(_02041_),
    .A1(_02042_),
    .S(_03664_),
    .X(_02043_));
 sky130_fd_sc_hd__mux4_1 _15191_ (.A0(\cpuregs.regs[12][7] ),
    .A1(\cpuregs.regs[13][7] ),
    .A2(\cpuregs.regs[14][7] ),
    .A3(\cpuregs.regs[15][7] ),
    .S0(_01936_),
    .S1(_03647_),
    .X(_02044_));
 sky130_fd_sc_hd__o21a_1 _15192_ (.A1(_03719_),
    .A2(_02044_),
    .B1(_00067_),
    .X(_02045_));
 sky130_fd_sc_hd__buf_6 _15193_ (.A(_03669_),
    .X(_02046_));
 sky130_fd_sc_hd__clkbuf_8 _15194_ (.A(_03646_),
    .X(_02047_));
 sky130_fd_sc_hd__mux4_1 _15195_ (.A0(\cpuregs.regs[8][7] ),
    .A1(\cpuregs.regs[9][7] ),
    .A2(\cpuregs.regs[10][7] ),
    .A3(\cpuregs.regs[11][7] ),
    .S0(_02046_),
    .S1(_02047_),
    .X(_02048_));
 sky130_fd_sc_hd__or2_1 _15196_ (.A(_03709_),
    .B(_02048_),
    .X(_02049_));
 sky130_fd_sc_hd__a221o_2 _15197_ (.A1(_02005_),
    .A2(_02043_),
    .B1(_02045_),
    .B2(_02049_),
    .C1(_03639_),
    .X(_02050_));
 sky130_fd_sc_hd__mux4_1 _15198_ (.A0(\cpuregs.regs[20][7] ),
    .A1(\cpuregs.regs[21][7] ),
    .A2(\cpuregs.regs[22][7] ),
    .A3(\cpuregs.regs[23][7] ),
    .S0(_03649_),
    .S1(_03643_),
    .X(_02051_));
 sky130_fd_sc_hd__mux4_1 _15199_ (.A0(\cpuregs.regs[16][7] ),
    .A1(\cpuregs.regs[17][7] ),
    .A2(\cpuregs.regs[18][7] ),
    .A3(\cpuregs.regs[19][7] ),
    .S0(_03645_),
    .S1(_01991_),
    .X(_02052_));
 sky130_fd_sc_hd__mux2_1 _15200_ (.A0(_02051_),
    .A1(_02052_),
    .S(_03719_),
    .X(_02053_));
 sky130_fd_sc_hd__mux4_1 _15201_ (.A0(\cpuregs.regs[24][7] ),
    .A1(\cpuregs.regs[25][7] ),
    .A2(\cpuregs.regs[26][7] ),
    .A3(\cpuregs.regs[27][7] ),
    .S0(_03661_),
    .S1(_03662_),
    .X(_02054_));
 sky130_fd_sc_hd__mux4_1 _15202_ (.A0(\cpuregs.regs[28][7] ),
    .A1(\cpuregs.regs[29][7] ),
    .A2(\cpuregs.regs[30][7] ),
    .A3(\cpuregs.regs[31][7] ),
    .S0(_03640_),
    .S1(_03642_),
    .X(_02055_));
 sky130_fd_sc_hd__mux2_1 _15203_ (.A0(_02054_),
    .A1(_02055_),
    .S(_03666_),
    .X(_02056_));
 sky130_fd_sc_hd__a21o_1 _15204_ (.A1(_03654_),
    .A2(_02056_),
    .B1(_03675_),
    .X(_02057_));
 sky130_fd_sc_hd__a21o_1 _15205_ (.A1(_02005_),
    .A2(_02053_),
    .B1(_02057_),
    .X(_02058_));
 sky130_fd_sc_hd__a32o_1 _15206_ (.A1(_01959_),
    .A2(_02050_),
    .A3(_02058_),
    .B1(_01933_),
    .B2(\decoded_imm[7] ),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _15207_ (.A0(net128),
    .A1(_02059_),
    .S(_01905_),
    .X(_02060_));
 sky130_fd_sc_hd__clkbuf_1 _15208_ (.A(_02060_),
    .X(_01160_));
 sky130_fd_sc_hd__mux4_1 _15209_ (.A0(\cpuregs.regs[20][8] ),
    .A1(\cpuregs.regs[21][8] ),
    .A2(\cpuregs.regs[22][8] ),
    .A3(\cpuregs.regs[23][8] ),
    .S0(_01970_),
    .S1(_01971_),
    .X(_02061_));
 sky130_fd_sc_hd__mux4_1 _15210_ (.A0(\cpuregs.regs[16][8] ),
    .A1(\cpuregs.regs[17][8] ),
    .A2(\cpuregs.regs[18][8] ),
    .A3(\cpuregs.regs[19][8] ),
    .S0(_01973_),
    .S1(_01974_),
    .X(_02062_));
 sky130_fd_sc_hd__mux4_1 _15211_ (.A0(\cpuregs.regs[4][8] ),
    .A1(\cpuregs.regs[5][8] ),
    .A2(\cpuregs.regs[6][8] ),
    .A3(\cpuregs.regs[7][8] ),
    .S0(_01976_),
    .S1(_01977_),
    .X(_02063_));
 sky130_fd_sc_hd__mux4_1 _15212_ (.A0(\cpuregs.regs[0][8] ),
    .A1(\cpuregs.regs[1][8] ),
    .A2(\cpuregs.regs[2][8] ),
    .A3(\cpuregs.regs[3][8] ),
    .S0(_01979_),
    .S1(_01980_),
    .X(_02064_));
 sky130_fd_sc_hd__mux4_1 _15213_ (.A0(_02061_),
    .A1(_02062_),
    .A2(_02063_),
    .A3(_02064_),
    .S0(_01982_),
    .S1(_02004_),
    .X(_02065_));
 sky130_fd_sc_hd__buf_6 _15214_ (.A(_03709_),
    .X(_02066_));
 sky130_fd_sc_hd__mux4_2 _15215_ (.A0(\cpuregs.regs[8][8] ),
    .A1(\cpuregs.regs[9][8] ),
    .A2(\cpuregs.regs[10][8] ),
    .A3(\cpuregs.regs[11][8] ),
    .S0(_01985_),
    .S1(_01986_),
    .X(_02067_));
 sky130_fd_sc_hd__or2_1 _15216_ (.A(_02066_),
    .B(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__buf_8 _15217_ (.A(_01936_),
    .X(_02069_));
 sky130_fd_sc_hd__buf_8 _15218_ (.A(_01991_),
    .X(_02070_));
 sky130_fd_sc_hd__mux4_1 _15219_ (.A0(\cpuregs.regs[12][8] ),
    .A1(\cpuregs.regs[13][8] ),
    .A2(\cpuregs.regs[14][8] ),
    .A3(\cpuregs.regs[15][8] ),
    .S0(_02069_),
    .S1(_02070_),
    .X(_02071_));
 sky130_fd_sc_hd__o21a_1 _15220_ (.A1(_02012_),
    .A2(_02071_),
    .B1(_02017_),
    .X(_02072_));
 sky130_fd_sc_hd__mux4_1 _15221_ (.A0(\cpuregs.regs[24][8] ),
    .A1(\cpuregs.regs[25][8] ),
    .A2(\cpuregs.regs[26][8] ),
    .A3(\cpuregs.regs[27][8] ),
    .S0(_01996_),
    .S1(_01997_),
    .X(_02073_));
 sky130_fd_sc_hd__buf_8 _15222_ (.A(_01995_),
    .X(_02074_));
 sky130_fd_sc_hd__buf_6 _15223_ (.A(_01937_),
    .X(_02075_));
 sky130_fd_sc_hd__mux4_1 _15224_ (.A0(\cpuregs.regs[28][8] ),
    .A1(\cpuregs.regs[29][8] ),
    .A2(\cpuregs.regs[30][8] ),
    .A3(\cpuregs.regs[31][8] ),
    .S0(_02074_),
    .S1(_02075_),
    .X(_02076_));
 sky130_fd_sc_hd__mux2_1 _15225_ (.A0(_02073_),
    .A1(_02076_),
    .S(_03687_),
    .X(_02077_));
 sky130_fd_sc_hd__a221o_1 _15226_ (.A1(_02068_),
    .A2(_02072_),
    .B1(_02077_),
    .B2(_02037_),
    .C1(_02006_),
    .X(_02078_));
 sky130_fd_sc_hd__o211a_4 _15227_ (.A1(_01969_),
    .A2(_02065_),
    .B1(_02078_),
    .C1(_01960_),
    .X(_02079_));
 sky130_fd_sc_hd__a21o_1 _15228_ (.A1(\decoded_imm[8] ),
    .A2(_02009_),
    .B1(_01963_),
    .X(_02080_));
 sky130_fd_sc_hd__o22a_1 _15229_ (.A1(net129),
    .A2(_01906_),
    .B1(_02079_),
    .B2(_02080_),
    .X(_01161_));
 sky130_fd_sc_hd__buf_2 _15230_ (.A(_01905_),
    .X(_02081_));
 sky130_fd_sc_hd__mux4_1 _15231_ (.A0(\cpuregs.regs[12][9] ),
    .A1(\cpuregs.regs[13][9] ),
    .A2(\cpuregs.regs[14][9] ),
    .A3(\cpuregs.regs[15][9] ),
    .S0(_01970_),
    .S1(_01971_),
    .X(_02082_));
 sky130_fd_sc_hd__mux4_1 _15232_ (.A0(\cpuregs.regs[8][9] ),
    .A1(\cpuregs.regs[9][9] ),
    .A2(\cpuregs.regs[10][9] ),
    .A3(\cpuregs.regs[11][9] ),
    .S0(_01973_),
    .S1(_01974_),
    .X(_02083_));
 sky130_fd_sc_hd__mux4_1 _15233_ (.A0(\cpuregs.regs[4][9] ),
    .A1(\cpuregs.regs[5][9] ),
    .A2(\cpuregs.regs[6][9] ),
    .A3(\cpuregs.regs[7][9] ),
    .S0(_01976_),
    .S1(_01977_),
    .X(_02084_));
 sky130_fd_sc_hd__buf_12 _15234_ (.A(_01918_),
    .X(_02085_));
 sky130_fd_sc_hd__buf_8 _15235_ (.A(_01919_),
    .X(_02086_));
 sky130_fd_sc_hd__mux4_1 _15236_ (.A0(\cpuregs.regs[0][9] ),
    .A1(\cpuregs.regs[1][9] ),
    .A2(\cpuregs.regs[2][9] ),
    .A3(\cpuregs.regs[3][9] ),
    .S0(_02085_),
    .S1(_02086_),
    .X(_02087_));
 sky130_fd_sc_hd__clkbuf_8 _15237_ (.A(_02005_),
    .X(_02088_));
 sky130_fd_sc_hd__mux4_1 _15238_ (.A0(_02082_),
    .A1(_02083_),
    .A2(_02084_),
    .A3(_02087_),
    .S0(_01982_),
    .S1(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__mux4_1 _15239_ (.A0(\cpuregs.regs[28][9] ),
    .A1(\cpuregs.regs[29][9] ),
    .A2(\cpuregs.regs[30][9] ),
    .A3(\cpuregs.regs[31][9] ),
    .S0(_01985_),
    .S1(_01986_),
    .X(_02090_));
 sky130_fd_sc_hd__or2_1 _15240_ (.A(_01984_),
    .B(_02090_),
    .X(_02091_));
 sky130_fd_sc_hd__mux4_1 _15241_ (.A0(\cpuregs.regs[24][9] ),
    .A1(\cpuregs.regs[25][9] ),
    .A2(\cpuregs.regs[26][9] ),
    .A3(\cpuregs.regs[27][9] ),
    .S0(_02069_),
    .S1(_02070_),
    .X(_02092_));
 sky130_fd_sc_hd__o21a_1 _15242_ (.A1(_01989_),
    .A2(_02092_),
    .B1(_03654_),
    .X(_02093_));
 sky130_fd_sc_hd__mux4_1 _15243_ (.A0(\cpuregs.regs[16][9] ),
    .A1(\cpuregs.regs[17][9] ),
    .A2(\cpuregs.regs[18][9] ),
    .A3(\cpuregs.regs[19][9] ),
    .S0(_01999_),
    .S1(_02000_),
    .X(_02094_));
 sky130_fd_sc_hd__mux4_1 _15244_ (.A0(\cpuregs.regs[20][9] ),
    .A1(\cpuregs.regs[21][9] ),
    .A2(\cpuregs.regs[22][9] ),
    .A3(\cpuregs.regs[23][9] ),
    .S0(_02074_),
    .S1(_02075_),
    .X(_02095_));
 sky130_fd_sc_hd__mux2_1 _15245_ (.A0(_02094_),
    .A1(_02095_),
    .S(_03687_),
    .X(_02096_));
 sky130_fd_sc_hd__a221o_1 _15246_ (.A1(_02091_),
    .A2(_02093_),
    .B1(_02096_),
    .B2(_02088_),
    .C1(_02018_),
    .X(_02097_));
 sky130_fd_sc_hd__o211a_4 _15247_ (.A1(_02020_),
    .A2(_02089_),
    .B1(_02097_),
    .C1(_01960_),
    .X(_02098_));
 sky130_fd_sc_hd__a21o_1 _15248_ (.A1(\decoded_imm[9] ),
    .A2(_02009_),
    .B1(_01963_),
    .X(_02099_));
 sky130_fd_sc_hd__o22a_1 _15249_ (.A1(net130),
    .A2(_02081_),
    .B1(_02098_),
    .B2(_02099_),
    .X(_01162_));
 sky130_fd_sc_hd__mux4_1 _15250_ (.A0(\cpuregs.regs[12][10] ),
    .A1(\cpuregs.regs[13][10] ),
    .A2(\cpuregs.regs[14][10] ),
    .A3(\cpuregs.regs[15][10] ),
    .S0(_01970_),
    .S1(_01971_),
    .X(_02100_));
 sky130_fd_sc_hd__mux4_1 _15251_ (.A0(\cpuregs.regs[8][10] ),
    .A1(\cpuregs.regs[9][10] ),
    .A2(\cpuregs.regs[10][10] ),
    .A3(\cpuregs.regs[11][10] ),
    .S0(_02013_),
    .S1(_02014_),
    .X(_02101_));
 sky130_fd_sc_hd__or2_1 _15252_ (.A(_01989_),
    .B(_02101_),
    .X(_02102_));
 sky130_fd_sc_hd__o211a_1 _15253_ (.A1(_01982_),
    .A2(_02100_),
    .B1(_02102_),
    .C1(_02018_),
    .X(_02103_));
 sky130_fd_sc_hd__mux4_1 _15254_ (.A0(\cpuregs.regs[24][10] ),
    .A1(\cpuregs.regs[25][10] ),
    .A2(\cpuregs.regs[26][10] ),
    .A3(\cpuregs.regs[27][10] ),
    .S0(_01990_),
    .S1(_01992_),
    .X(_02104_));
 sky130_fd_sc_hd__mux4_1 _15255_ (.A0(\cpuregs.regs[28][10] ),
    .A1(\cpuregs.regs[29][10] ),
    .A2(\cpuregs.regs[30][10] ),
    .A3(\cpuregs.regs[31][10] ),
    .S0(_02022_),
    .S1(_02023_),
    .X(_02105_));
 sky130_fd_sc_hd__mux2_1 _15256_ (.A0(_02104_),
    .A1(_02105_),
    .S(_03687_),
    .X(_02106_));
 sky130_fd_sc_hd__a21o_1 _15257_ (.A1(_02020_),
    .A2(_02106_),
    .B1(_02006_),
    .X(_02107_));
 sky130_fd_sc_hd__mux4_1 _15258_ (.A0(\cpuregs.regs[0][10] ),
    .A1(\cpuregs.regs[1][10] ),
    .A2(\cpuregs.regs[2][10] ),
    .A3(\cpuregs.regs[3][10] ),
    .S0(_01990_),
    .S1(_01992_),
    .X(_02108_));
 sky130_fd_sc_hd__or2_1 _15259_ (.A(_02066_),
    .B(_02108_),
    .X(_02109_));
 sky130_fd_sc_hd__clkbuf_8 _15260_ (.A(_03664_),
    .X(_02110_));
 sky130_fd_sc_hd__clkbuf_8 _15261_ (.A(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__mux4_1 _15262_ (.A0(\cpuregs.regs[4][10] ),
    .A1(\cpuregs.regs[5][10] ),
    .A2(\cpuregs.regs[6][10] ),
    .A3(\cpuregs.regs[7][10] ),
    .S0(_02013_),
    .S1(_02014_),
    .X(_02112_));
 sky130_fd_sc_hd__o21a_1 _15263_ (.A1(_02111_),
    .A2(_02112_),
    .B1(_02017_),
    .X(_02113_));
 sky130_fd_sc_hd__mux4_1 _15264_ (.A0(\cpuregs.regs[20][10] ),
    .A1(\cpuregs.regs[21][10] ),
    .A2(\cpuregs.regs[22][10] ),
    .A3(\cpuregs.regs[23][10] ),
    .S0(_02022_),
    .S1(_02023_),
    .X(_02114_));
 sky130_fd_sc_hd__mux4_1 _15265_ (.A0(\cpuregs.regs[16][10] ),
    .A1(\cpuregs.regs[17][10] ),
    .A2(\cpuregs.regs[18][10] ),
    .A3(\cpuregs.regs[19][10] ),
    .S0(_01985_),
    .S1(_01986_),
    .X(_02115_));
 sky130_fd_sc_hd__mux2_1 _15266_ (.A0(_02114_),
    .A1(_02115_),
    .S(_02002_),
    .X(_02116_));
 sky130_fd_sc_hd__a221o_1 _15267_ (.A1(_02109_),
    .A2(_02113_),
    .B1(_02116_),
    .B2(_02037_),
    .C1(_01969_),
    .X(_02117_));
 sky130_fd_sc_hd__o211a_4 _15268_ (.A1(_02103_),
    .A2(_02107_),
    .B1(_02027_),
    .C1(_02117_),
    .X(_02118_));
 sky130_fd_sc_hd__a21o_1 _15269_ (.A1(\decoded_imm[10] ),
    .A2(_02009_),
    .B1(_01963_),
    .X(_02119_));
 sky130_fd_sc_hd__o22a_1 _15270_ (.A1(net100),
    .A2(_02081_),
    .B1(_02118_),
    .B2(_02119_),
    .X(_01163_));
 sky130_fd_sc_hd__mux4_1 _15271_ (.A0(\cpuregs.regs[12][11] ),
    .A1(\cpuregs.regs[13][11] ),
    .A2(\cpuregs.regs[14][11] ),
    .A3(\cpuregs.regs[15][11] ),
    .S0(_01970_),
    .S1(_01971_),
    .X(_02120_));
 sky130_fd_sc_hd__mux4_1 _15272_ (.A0(\cpuregs.regs[8][11] ),
    .A1(\cpuregs.regs[9][11] ),
    .A2(\cpuregs.regs[10][11] ),
    .A3(\cpuregs.regs[11][11] ),
    .S0(_01973_),
    .S1(_01974_),
    .X(_02121_));
 sky130_fd_sc_hd__mux4_1 _15273_ (.A0(\cpuregs.regs[4][11] ),
    .A1(\cpuregs.regs[5][11] ),
    .A2(\cpuregs.regs[6][11] ),
    .A3(\cpuregs.regs[7][11] ),
    .S0(_01976_),
    .S1(_01977_),
    .X(_02122_));
 sky130_fd_sc_hd__mux4_1 _15274_ (.A0(\cpuregs.regs[0][11] ),
    .A1(\cpuregs.regs[1][11] ),
    .A2(\cpuregs.regs[2][11] ),
    .A3(\cpuregs.regs[3][11] ),
    .S0(_02085_),
    .S1(_02086_),
    .X(_02123_));
 sky130_fd_sc_hd__mux4_1 _15275_ (.A0(_02120_),
    .A1(_02121_),
    .A2(_02122_),
    .A3(_02123_),
    .S0(_01982_),
    .S1(_02088_),
    .X(_02124_));
 sky130_fd_sc_hd__mux4_1 _15276_ (.A0(\cpuregs.regs[16][11] ),
    .A1(\cpuregs.regs[17][11] ),
    .A2(\cpuregs.regs[18][11] ),
    .A3(\cpuregs.regs[19][11] ),
    .S0(_01985_),
    .S1(_01986_),
    .X(_02125_));
 sky130_fd_sc_hd__or2_1 _15277_ (.A(_02066_),
    .B(_02125_),
    .X(_02126_));
 sky130_fd_sc_hd__mux4_1 _15278_ (.A0(\cpuregs.regs[20][11] ),
    .A1(\cpuregs.regs[21][11] ),
    .A2(\cpuregs.regs[22][11] ),
    .A3(\cpuregs.regs[23][11] ),
    .S0(_02069_),
    .S1(_02070_),
    .X(_02127_));
 sky130_fd_sc_hd__o21a_1 _15279_ (.A1(_02012_),
    .A2(_02127_),
    .B1(_02005_),
    .X(_02128_));
 sky130_fd_sc_hd__mux4_1 _15280_ (.A0(\cpuregs.regs[28][11] ),
    .A1(\cpuregs.regs[29][11] ),
    .A2(\cpuregs.regs[30][11] ),
    .A3(\cpuregs.regs[31][11] ),
    .S0(_01999_),
    .S1(_02000_),
    .X(_02129_));
 sky130_fd_sc_hd__mux4_1 _15281_ (.A0(\cpuregs.regs[24][11] ),
    .A1(\cpuregs.regs[25][11] ),
    .A2(\cpuregs.regs[26][11] ),
    .A3(\cpuregs.regs[27][11] ),
    .S0(_02074_),
    .S1(_02075_),
    .X(_02130_));
 sky130_fd_sc_hd__mux2_1 _15282_ (.A0(_02129_),
    .A1(_02130_),
    .S(_02002_),
    .X(_02131_));
 sky130_fd_sc_hd__a221o_1 _15283_ (.A1(_02126_),
    .A2(_02128_),
    .B1(_02131_),
    .B2(_03683_),
    .C1(_02018_),
    .X(_02132_));
 sky130_fd_sc_hd__o211a_2 _15284_ (.A1(_02020_),
    .A2(_02124_),
    .B1(_02132_),
    .C1(_01960_),
    .X(_02133_));
 sky130_fd_sc_hd__a21o_1 _15285_ (.A1(\decoded_imm[11] ),
    .A2(_02009_),
    .B1(_01963_),
    .X(_02134_));
 sky130_fd_sc_hd__o22a_1 _15286_ (.A1(net101),
    .A2(_02081_),
    .B1(_02133_),
    .B2(_02134_),
    .X(_01164_));
 sky130_fd_sc_hd__mux4_1 _15287_ (.A0(\cpuregs.regs[4][12] ),
    .A1(\cpuregs.regs[5][12] ),
    .A2(\cpuregs.regs[6][12] ),
    .A3(\cpuregs.regs[7][12] ),
    .S0(_01970_),
    .S1(_01971_),
    .X(_02135_));
 sky130_fd_sc_hd__mux4_1 _15288_ (.A0(\cpuregs.regs[0][12] ),
    .A1(\cpuregs.regs[1][12] ),
    .A2(\cpuregs.regs[2][12] ),
    .A3(\cpuregs.regs[3][12] ),
    .S0(_01973_),
    .S1(_01974_),
    .X(_02136_));
 sky130_fd_sc_hd__mux4_1 _15289_ (.A0(\cpuregs.regs[12][12] ),
    .A1(\cpuregs.regs[13][12] ),
    .A2(\cpuregs.regs[14][12] ),
    .A3(\cpuregs.regs[15][12] ),
    .S0(_01976_),
    .S1(_01977_),
    .X(_02137_));
 sky130_fd_sc_hd__mux4_1 _15290_ (.A0(\cpuregs.regs[8][12] ),
    .A1(\cpuregs.regs[9][12] ),
    .A2(\cpuregs.regs[10][12] ),
    .A3(\cpuregs.regs[11][12] ),
    .S0(_02085_),
    .S1(_02086_),
    .X(_02138_));
 sky130_fd_sc_hd__mux4_1 _15291_ (.A0(_02135_),
    .A1(_02136_),
    .A2(_02137_),
    .A3(_02138_),
    .S0(_01982_),
    .S1(_03683_),
    .X(_02139_));
 sky130_fd_sc_hd__mux4_1 _15292_ (.A0(\cpuregs.regs[28][12] ),
    .A1(\cpuregs.regs[29][12] ),
    .A2(\cpuregs.regs[30][12] ),
    .A3(\cpuregs.regs[31][12] ),
    .S0(_01985_),
    .S1(_01986_),
    .X(_02140_));
 sky130_fd_sc_hd__or2_1 _15293_ (.A(_01984_),
    .B(_02140_),
    .X(_02141_));
 sky130_fd_sc_hd__mux4_1 _15294_ (.A0(\cpuregs.regs[24][12] ),
    .A1(\cpuregs.regs[25][12] ),
    .A2(\cpuregs.regs[26][12] ),
    .A3(\cpuregs.regs[27][12] ),
    .S0(_02069_),
    .S1(_02070_),
    .X(_02142_));
 sky130_fd_sc_hd__o21a_1 _15295_ (.A1(_02066_),
    .A2(_02142_),
    .B1(_03654_),
    .X(_02143_));
 sky130_fd_sc_hd__mux4_1 _15296_ (.A0(\cpuregs.regs[20][12] ),
    .A1(\cpuregs.regs[21][12] ),
    .A2(\cpuregs.regs[22][12] ),
    .A3(\cpuregs.regs[23][12] ),
    .S0(_01999_),
    .S1(_02000_),
    .X(_02144_));
 sky130_fd_sc_hd__mux4_1 _15297_ (.A0(\cpuregs.regs[16][12] ),
    .A1(\cpuregs.regs[17][12] ),
    .A2(\cpuregs.regs[18][12] ),
    .A3(\cpuregs.regs[19][12] ),
    .S0(_02074_),
    .S1(_02075_),
    .X(_02145_));
 sky130_fd_sc_hd__mux2_1 _15298_ (.A0(_02144_),
    .A1(_02145_),
    .S(_02002_),
    .X(_02146_));
 sky130_fd_sc_hd__a221o_1 _15299_ (.A1(_02141_),
    .A2(_02143_),
    .B1(_02146_),
    .B2(_02088_),
    .C1(_02018_),
    .X(_02147_));
 sky130_fd_sc_hd__o211a_4 _15300_ (.A1(_02020_),
    .A2(_02139_),
    .B1(_02147_),
    .C1(_01960_),
    .X(_02148_));
 sky130_fd_sc_hd__a21o_1 _15301_ (.A1(\decoded_imm[12] ),
    .A2(_02009_),
    .B1(_01963_),
    .X(_02149_));
 sky130_fd_sc_hd__o22a_1 _15302_ (.A1(net102),
    .A2(_02081_),
    .B1(_02148_),
    .B2(_02149_),
    .X(_01165_));
 sky130_fd_sc_hd__mux4_1 _15303_ (.A0(\cpuregs.regs[12][13] ),
    .A1(\cpuregs.regs[13][13] ),
    .A2(\cpuregs.regs[14][13] ),
    .A3(\cpuregs.regs[15][13] ),
    .S0(_01970_),
    .S1(_01971_),
    .X(_02150_));
 sky130_fd_sc_hd__mux4_1 _15304_ (.A0(\cpuregs.regs[8][13] ),
    .A1(\cpuregs.regs[9][13] ),
    .A2(\cpuregs.regs[10][13] ),
    .A3(\cpuregs.regs[11][13] ),
    .S0(_02013_),
    .S1(_02014_),
    .X(_02151_));
 sky130_fd_sc_hd__or2_1 _15305_ (.A(_01989_),
    .B(_02151_),
    .X(_02152_));
 sky130_fd_sc_hd__o211a_1 _15306_ (.A1(_01982_),
    .A2(_02150_),
    .B1(_02152_),
    .C1(_02018_),
    .X(_02153_));
 sky130_fd_sc_hd__mux4_1 _15307_ (.A0(\cpuregs.regs[28][13] ),
    .A1(\cpuregs.regs[29][13] ),
    .A2(\cpuregs.regs[30][13] ),
    .A3(\cpuregs.regs[31][13] ),
    .S0(_01990_),
    .S1(_01992_),
    .X(_02154_));
 sky130_fd_sc_hd__mux4_1 _15308_ (.A0(\cpuregs.regs[24][13] ),
    .A1(\cpuregs.regs[25][13] ),
    .A2(\cpuregs.regs[26][13] ),
    .A3(\cpuregs.regs[27][13] ),
    .S0(_02022_),
    .S1(_02023_),
    .X(_02155_));
 sky130_fd_sc_hd__mux2_1 _15309_ (.A0(_02154_),
    .A1(_02155_),
    .S(_01984_),
    .X(_02156_));
 sky130_fd_sc_hd__a21o_1 _15310_ (.A1(_02037_),
    .A2(_02156_),
    .B1(_02006_),
    .X(_02157_));
 sky130_fd_sc_hd__mux4_1 _15311_ (.A0(\cpuregs.regs[20][13] ),
    .A1(\cpuregs.regs[21][13] ),
    .A2(\cpuregs.regs[22][13] ),
    .A3(\cpuregs.regs[23][13] ),
    .S0(_01990_),
    .S1(_01992_),
    .X(_02158_));
 sky130_fd_sc_hd__or2_1 _15312_ (.A(_02012_),
    .B(_02158_),
    .X(_02159_));
 sky130_fd_sc_hd__mux4_1 _15313_ (.A0(\cpuregs.regs[16][13] ),
    .A1(\cpuregs.regs[17][13] ),
    .A2(\cpuregs.regs[18][13] ),
    .A3(\cpuregs.regs[19][13] ),
    .S0(_02013_),
    .S1(_02014_),
    .X(_02160_));
 sky130_fd_sc_hd__o21a_1 _15314_ (.A1(_01989_),
    .A2(_02160_),
    .B1(_03639_),
    .X(_02161_));
 sky130_fd_sc_hd__mux4_1 _15315_ (.A0(\cpuregs.regs[4][13] ),
    .A1(\cpuregs.regs[5][13] ),
    .A2(\cpuregs.regs[6][13] ),
    .A3(\cpuregs.regs[7][13] ),
    .S0(_02022_),
    .S1(_02023_),
    .X(_02162_));
 sky130_fd_sc_hd__mux4_1 _15316_ (.A0(\cpuregs.regs[0][13] ),
    .A1(\cpuregs.regs[1][13] ),
    .A2(\cpuregs.regs[2][13] ),
    .A3(\cpuregs.regs[3][13] ),
    .S0(_01985_),
    .S1(_01986_),
    .X(_02163_));
 sky130_fd_sc_hd__mux2_1 _15317_ (.A0(_02162_),
    .A1(_02163_),
    .S(_02002_),
    .X(_02164_));
 sky130_fd_sc_hd__a221o_1 _15318_ (.A1(_02159_),
    .A2(_02161_),
    .B1(_02164_),
    .B2(_02004_),
    .C1(_01969_),
    .X(_02165_));
 sky130_fd_sc_hd__o211a_4 _15319_ (.A1(_02153_),
    .A2(_02157_),
    .B1(_02027_),
    .C1(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__a21o_1 _15320_ (.A1(\decoded_imm[13] ),
    .A2(_02009_),
    .B1(_01963_),
    .X(_02167_));
 sky130_fd_sc_hd__o22a_1 _15321_ (.A1(net103),
    .A2(_02081_),
    .B1(_02166_),
    .B2(_02167_),
    .X(_01166_));
 sky130_fd_sc_hd__mux4_1 _15322_ (.A0(\cpuregs.regs[4][14] ),
    .A1(\cpuregs.regs[5][14] ),
    .A2(\cpuregs.regs[6][14] ),
    .A3(\cpuregs.regs[7][14] ),
    .S0(_01979_),
    .S1(_01980_),
    .X(_02168_));
 sky130_fd_sc_hd__mux4_1 _15323_ (.A0(\cpuregs.regs[0][14] ),
    .A1(\cpuregs.regs[1][14] ),
    .A2(\cpuregs.regs[2][14] ),
    .A3(\cpuregs.regs[3][14] ),
    .S0(_01973_),
    .S1(_01974_),
    .X(_02169_));
 sky130_fd_sc_hd__mux4_1 _15324_ (.A0(\cpuregs.regs[20][14] ),
    .A1(\cpuregs.regs[21][14] ),
    .A2(\cpuregs.regs[22][14] ),
    .A3(\cpuregs.regs[23][14] ),
    .S0(_01976_),
    .S1(_01977_),
    .X(_02170_));
 sky130_fd_sc_hd__mux4_1 _15325_ (.A0(\cpuregs.regs[16][14] ),
    .A1(\cpuregs.regs[17][14] ),
    .A2(\cpuregs.regs[18][14] ),
    .A3(\cpuregs.regs[19][14] ),
    .S0(_02085_),
    .S1(_02086_),
    .X(_02171_));
 sky130_fd_sc_hd__mux4_1 _15326_ (.A0(_02168_),
    .A1(_02169_),
    .A2(_02170_),
    .A3(_02171_),
    .S0(_01982_),
    .S1(_03639_),
    .X(_02172_));
 sky130_fd_sc_hd__mux4_1 _15327_ (.A0(\cpuregs.regs[8][14] ),
    .A1(\cpuregs.regs[9][14] ),
    .A2(\cpuregs.regs[10][14] ),
    .A3(\cpuregs.regs[11][14] ),
    .S0(_01996_),
    .S1(_01997_),
    .X(_02173_));
 sky130_fd_sc_hd__or2_1 _15328_ (.A(_02066_),
    .B(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__mux4_1 _15329_ (.A0(\cpuregs.regs[12][14] ),
    .A1(\cpuregs.regs[13][14] ),
    .A2(\cpuregs.regs[14][14] ),
    .A3(\cpuregs.regs[15][14] ),
    .S0(_02069_),
    .S1(_02070_),
    .X(_02175_));
 sky130_fd_sc_hd__o21a_1 _15330_ (.A1(_02012_),
    .A2(_02175_),
    .B1(_02017_),
    .X(_02176_));
 sky130_fd_sc_hd__mux4_1 _15331_ (.A0(\cpuregs.regs[28][14] ),
    .A1(\cpuregs.regs[29][14] ),
    .A2(\cpuregs.regs[30][14] ),
    .A3(\cpuregs.regs[31][14] ),
    .S0(_01999_),
    .S1(_02000_),
    .X(_02177_));
 sky130_fd_sc_hd__mux4_1 _15332_ (.A0(\cpuregs.regs[24][14] ),
    .A1(\cpuregs.regs[25][14] ),
    .A2(\cpuregs.regs[26][14] ),
    .A3(\cpuregs.regs[27][14] ),
    .S0(_02074_),
    .S1(_02075_),
    .X(_02178_));
 sky130_fd_sc_hd__mux2_1 _15333_ (.A0(_02177_),
    .A1(_02178_),
    .S(_02002_),
    .X(_02179_));
 sky130_fd_sc_hd__a221o_1 _15334_ (.A1(_02174_),
    .A2(_02176_),
    .B1(_02179_),
    .B2(_02037_),
    .C1(_02006_),
    .X(_02180_));
 sky130_fd_sc_hd__o211a_4 _15335_ (.A1(_01969_),
    .A2(_02172_),
    .B1(_02180_),
    .C1(_01960_),
    .X(_02181_));
 sky130_fd_sc_hd__a21o_1 _15336_ (.A1(\decoded_imm[14] ),
    .A2(_02009_),
    .B1(_01963_),
    .X(_02182_));
 sky130_fd_sc_hd__o22a_1 _15337_ (.A1(net104),
    .A2(_02081_),
    .B1(_02181_),
    .B2(_02182_),
    .X(_01167_));
 sky130_fd_sc_hd__mux4_1 _15338_ (.A0(\cpuregs.regs[12][15] ),
    .A1(\cpuregs.regs[13][15] ),
    .A2(\cpuregs.regs[14][15] ),
    .A3(\cpuregs.regs[15][15] ),
    .S0(_01979_),
    .S1(_01980_),
    .X(_02183_));
 sky130_fd_sc_hd__mux4_1 _15339_ (.A0(\cpuregs.regs[8][15] ),
    .A1(\cpuregs.regs[9][15] ),
    .A2(\cpuregs.regs[10][15] ),
    .A3(\cpuregs.regs[11][15] ),
    .S0(_02030_),
    .S1(_02031_),
    .X(_02184_));
 sky130_fd_sc_hd__mux4_1 _15340_ (.A0(\cpuregs.regs[4][15] ),
    .A1(\cpuregs.regs[5][15] ),
    .A2(\cpuregs.regs[6][15] ),
    .A3(\cpuregs.regs[7][15] ),
    .S0(_01976_),
    .S1(_01977_),
    .X(_02185_));
 sky130_fd_sc_hd__mux4_1 _15341_ (.A0(\cpuregs.regs[0][15] ),
    .A1(\cpuregs.regs[1][15] ),
    .A2(\cpuregs.regs[2][15] ),
    .A3(\cpuregs.regs[3][15] ),
    .S0(_02085_),
    .S1(_02086_),
    .X(_02186_));
 sky130_fd_sc_hd__mux4_1 _15342_ (.A0(_02183_),
    .A1(_02184_),
    .A2(_02185_),
    .A3(_02186_),
    .S0(_02111_),
    .S1(_02088_),
    .X(_02187_));
 sky130_fd_sc_hd__mux4_1 _15343_ (.A0(\cpuregs.regs[16][15] ),
    .A1(\cpuregs.regs[17][15] ),
    .A2(\cpuregs.regs[18][15] ),
    .A3(\cpuregs.regs[19][15] ),
    .S0(_01996_),
    .S1(_01997_),
    .X(_02188_));
 sky130_fd_sc_hd__or2_1 _15344_ (.A(_02066_),
    .B(_02188_),
    .X(_02189_));
 sky130_fd_sc_hd__mux4_1 _15345_ (.A0(\cpuregs.regs[20][15] ),
    .A1(\cpuregs.regs[21][15] ),
    .A2(\cpuregs.regs[22][15] ),
    .A3(\cpuregs.regs[23][15] ),
    .S0(_02069_),
    .S1(_02070_),
    .X(_02190_));
 sky130_fd_sc_hd__o21a_1 _15346_ (.A1(_02012_),
    .A2(_02190_),
    .B1(_02005_),
    .X(_02191_));
 sky130_fd_sc_hd__mux4_1 _15347_ (.A0(\cpuregs.regs[28][15] ),
    .A1(\cpuregs.regs[29][15] ),
    .A2(\cpuregs.regs[30][15] ),
    .A3(\cpuregs.regs[31][15] ),
    .S0(_01999_),
    .S1(_02000_),
    .X(_02192_));
 sky130_fd_sc_hd__mux4_1 _15348_ (.A0(\cpuregs.regs[24][15] ),
    .A1(\cpuregs.regs[25][15] ),
    .A2(\cpuregs.regs[26][15] ),
    .A3(\cpuregs.regs[27][15] ),
    .S0(_02074_),
    .S1(_02075_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_1 _15349_ (.A0(_02192_),
    .A1(_02193_),
    .S(_02002_),
    .X(_02194_));
 sky130_fd_sc_hd__a221o_1 _15350_ (.A1(_02189_),
    .A2(_02191_),
    .B1(_02194_),
    .B2(_03683_),
    .C1(_02018_),
    .X(_02195_));
 sky130_fd_sc_hd__o211a_4 _15351_ (.A1(_02020_),
    .A2(_02187_),
    .B1(_02195_),
    .C1(_01960_),
    .X(_02196_));
 sky130_fd_sc_hd__clkbuf_4 _15352_ (.A(_01934_),
    .X(_02197_));
 sky130_fd_sc_hd__a21o_1 _15353_ (.A1(\decoded_imm[15] ),
    .A2(_02009_),
    .B1(_02197_),
    .X(_02198_));
 sky130_fd_sc_hd__o22a_1 _15354_ (.A1(net105),
    .A2(_02081_),
    .B1(_02196_),
    .B2(_02198_),
    .X(_01168_));
 sky130_fd_sc_hd__mux4_1 _15355_ (.A0(\cpuregs.regs[20][16] ),
    .A1(\cpuregs.regs[21][16] ),
    .A2(\cpuregs.regs[22][16] ),
    .A3(\cpuregs.regs[23][16] ),
    .S0(_01970_),
    .S1(_01971_),
    .X(_02199_));
 sky130_fd_sc_hd__mux4_1 _15356_ (.A0(\cpuregs.regs[16][16] ),
    .A1(\cpuregs.regs[17][16] ),
    .A2(\cpuregs.regs[18][16] ),
    .A3(\cpuregs.regs[19][16] ),
    .S0(_02013_),
    .S1(_02014_),
    .X(_02200_));
 sky130_fd_sc_hd__or2_1 _15357_ (.A(_01989_),
    .B(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__o211a_1 _15358_ (.A1(_01982_),
    .A2(_02199_),
    .B1(_02201_),
    .C1(_02006_),
    .X(_02202_));
 sky130_fd_sc_hd__mux4_1 _15359_ (.A0(\cpuregs.regs[28][16] ),
    .A1(\cpuregs.regs[29][16] ),
    .A2(\cpuregs.regs[30][16] ),
    .A3(\cpuregs.regs[31][16] ),
    .S0(_01990_),
    .S1(_01992_),
    .X(_02203_));
 sky130_fd_sc_hd__mux4_1 _15360_ (.A0(\cpuregs.regs[24][16] ),
    .A1(\cpuregs.regs[25][16] ),
    .A2(\cpuregs.regs[26][16] ),
    .A3(\cpuregs.regs[27][16] ),
    .S0(_02022_),
    .S1(_02023_),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_1 _15361_ (.A0(_02203_),
    .A1(_02204_),
    .S(_01984_),
    .X(_02205_));
 sky130_fd_sc_hd__a21o_1 _15362_ (.A1(_03683_),
    .A2(_02205_),
    .B1(_02018_),
    .X(_02206_));
 sky130_fd_sc_hd__mux4_1 _15363_ (.A0(\cpuregs.regs[8][16] ),
    .A1(\cpuregs.regs[9][16] ),
    .A2(\cpuregs.regs[10][16] ),
    .A3(\cpuregs.regs[11][16] ),
    .S0(_01990_),
    .S1(_01992_),
    .X(_02207_));
 sky130_fd_sc_hd__or2_1 _15364_ (.A(_02066_),
    .B(_02207_),
    .X(_02208_));
 sky130_fd_sc_hd__mux4_1 _15365_ (.A0(\cpuregs.regs[12][16] ),
    .A1(\cpuregs.regs[13][16] ),
    .A2(\cpuregs.regs[14][16] ),
    .A3(\cpuregs.regs[15][16] ),
    .S0(_02013_),
    .S1(_02014_),
    .X(_02209_));
 sky130_fd_sc_hd__o21a_1 _15366_ (.A1(_02012_),
    .A2(_02209_),
    .B1(_01968_),
    .X(_02210_));
 sky130_fd_sc_hd__mux4_1 _15367_ (.A0(\cpuregs.regs[4][16] ),
    .A1(\cpuregs.regs[5][16] ),
    .A2(\cpuregs.regs[6][16] ),
    .A3(\cpuregs.regs[7][16] ),
    .S0(_02022_),
    .S1(_02023_),
    .X(_02211_));
 sky130_fd_sc_hd__mux4_1 _15368_ (.A0(\cpuregs.regs[0][16] ),
    .A1(\cpuregs.regs[1][16] ),
    .A2(\cpuregs.regs[2][16] ),
    .A3(\cpuregs.regs[3][16] ),
    .S0(_01985_),
    .S1(_01986_),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_1 _15369_ (.A0(_02211_),
    .A1(_02212_),
    .S(_02002_),
    .X(_02213_));
 sky130_fd_sc_hd__a221o_1 _15370_ (.A1(_02208_),
    .A2(_02210_),
    .B1(_02213_),
    .B2(_02088_),
    .C1(_02020_),
    .X(_02214_));
 sky130_fd_sc_hd__o211a_4 _15371_ (.A1(_02202_),
    .A2(_02206_),
    .B1(_02027_),
    .C1(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__buf_4 _15372_ (.A(_01932_),
    .X(_02216_));
 sky130_fd_sc_hd__a21o_1 _15373_ (.A1(\decoded_imm[16] ),
    .A2(_02216_),
    .B1(_02197_),
    .X(_02217_));
 sky130_fd_sc_hd__o22a_1 _15374_ (.A1(net106),
    .A2(_02081_),
    .B1(_02215_),
    .B2(_02217_),
    .X(_01169_));
 sky130_fd_sc_hd__mux4_1 _15375_ (.A0(\cpuregs.regs[4][17] ),
    .A1(\cpuregs.regs[5][17] ),
    .A2(\cpuregs.regs[6][17] ),
    .A3(\cpuregs.regs[7][17] ),
    .S0(_01908_),
    .S1(_01909_),
    .X(_02218_));
 sky130_fd_sc_hd__mux4_1 _15376_ (.A0(\cpuregs.regs[0][17] ),
    .A1(\cpuregs.regs[1][17] ),
    .A2(\cpuregs.regs[2][17] ),
    .A3(\cpuregs.regs[3][17] ),
    .S0(_01908_),
    .S1(_01909_),
    .X(_02219_));
 sky130_fd_sc_hd__mux2_1 _15377_ (.A0(_02218_),
    .A1(_02219_),
    .S(_01907_),
    .X(_02220_));
 sky130_fd_sc_hd__buf_6 _15378_ (.A(_03658_),
    .X(_02221_));
 sky130_fd_sc_hd__clkbuf_8 _15379_ (.A(_03659_),
    .X(_02222_));
 sky130_fd_sc_hd__mux4_1 _15380_ (.A0(\cpuregs.regs[12][17] ),
    .A1(\cpuregs.regs[13][17] ),
    .A2(\cpuregs.regs[14][17] ),
    .A3(\cpuregs.regs[15][17] ),
    .S0(_02221_),
    .S1(_02222_),
    .X(_02223_));
 sky130_fd_sc_hd__mux4_1 _15381_ (.A0(\cpuregs.regs[8][17] ),
    .A1(\cpuregs.regs[9][17] ),
    .A2(\cpuregs.regs[10][17] ),
    .A3(\cpuregs.regs[11][17] ),
    .S0(_03641_),
    .S1(_03684_),
    .X(_02224_));
 sky130_fd_sc_hd__mux2_1 _15382_ (.A0(_02223_),
    .A1(_02224_),
    .S(_02110_),
    .X(_02225_));
 sky130_fd_sc_hd__mux4_1 _15383_ (.A0(\cpuregs.regs[20][17] ),
    .A1(\cpuregs.regs[21][17] ),
    .A2(\cpuregs.regs[22][17] ),
    .A3(\cpuregs.regs[23][17] ),
    .S0(_02221_),
    .S1(_02222_),
    .X(_02226_));
 sky130_fd_sc_hd__mux4_1 _15384_ (.A0(\cpuregs.regs[16][17] ),
    .A1(\cpuregs.regs[17][17] ),
    .A2(\cpuregs.regs[18][17] ),
    .A3(\cpuregs.regs[19][17] ),
    .S0(_02221_),
    .S1(_02222_),
    .X(_02227_));
 sky130_fd_sc_hd__mux2_1 _15385_ (.A0(_02226_),
    .A1(_02227_),
    .S(_02110_),
    .X(_02228_));
 sky130_fd_sc_hd__mux4_1 _15386_ (.A0(\cpuregs.regs[28][17] ),
    .A1(\cpuregs.regs[29][17] ),
    .A2(\cpuregs.regs[30][17] ),
    .A3(\cpuregs.regs[31][17] ),
    .S0(_01908_),
    .S1(_01909_),
    .X(_02229_));
 sky130_fd_sc_hd__mux4_1 _15387_ (.A0(\cpuregs.regs[24][17] ),
    .A1(\cpuregs.regs[25][17] ),
    .A2(\cpuregs.regs[26][17] ),
    .A3(\cpuregs.regs[27][17] ),
    .S0(_02221_),
    .S1(_02222_),
    .X(_02230_));
 sky130_fd_sc_hd__mux2_1 _15388_ (.A0(_02229_),
    .A1(_02230_),
    .S(_02110_),
    .X(_02231_));
 sky130_fd_sc_hd__mux4_2 _15389_ (.A0(_02220_),
    .A1(_02225_),
    .A2(_02228_),
    .A3(_02231_),
    .S0(_01968_),
    .S1(_02037_),
    .X(_02232_));
 sky130_fd_sc_hd__a221o_2 _15390_ (.A1(\decoded_imm[17] ),
    .A2(_02216_),
    .B1(_02027_),
    .B2(_02232_),
    .C1(_02197_),
    .X(_02233_));
 sky130_fd_sc_hd__o21a_1 _15391_ (.A1(net107),
    .A2(_01906_),
    .B1(_02233_),
    .X(_01170_));
 sky130_fd_sc_hd__mux4_1 _15392_ (.A0(\cpuregs.regs[20][18] ),
    .A1(\cpuregs.regs[21][18] ),
    .A2(\cpuregs.regs[22][18] ),
    .A3(\cpuregs.regs[23][18] ),
    .S0(_01995_),
    .S1(_01937_),
    .X(_02234_));
 sky130_fd_sc_hd__or2_1 _15393_ (.A(_03653_),
    .B(_02234_),
    .X(_02235_));
 sky130_fd_sc_hd__mux4_1 _15394_ (.A0(\cpuregs.regs[16][18] ),
    .A1(\cpuregs.regs[17][18] ),
    .A2(\cpuregs.regs[18][18] ),
    .A3(\cpuregs.regs[19][18] ),
    .S0(_01936_),
    .S1(_01937_),
    .X(_02236_));
 sky130_fd_sc_hd__o21a_1 _15395_ (.A1(_03709_),
    .A2(_02236_),
    .B1(_00068_),
    .X(_02237_));
 sky130_fd_sc_hd__mux4_1 _15396_ (.A0(\cpuregs.regs[4][18] ),
    .A1(\cpuregs.regs[5][18] ),
    .A2(\cpuregs.regs[6][18] ),
    .A3(\cpuregs.regs[7][18] ),
    .S0(_02046_),
    .S1(_02047_),
    .X(_02238_));
 sky130_fd_sc_hd__mux4_1 _15397_ (.A0(\cpuregs.regs[0][18] ),
    .A1(\cpuregs.regs[1][18] ),
    .A2(\cpuregs.regs[2][18] ),
    .A3(\cpuregs.regs[3][18] ),
    .S0(_02046_),
    .S1(_02047_),
    .X(_02239_));
 sky130_fd_sc_hd__mux2_1 _15398_ (.A0(_02238_),
    .A1(_02239_),
    .S(_03653_),
    .X(_02240_));
 sky130_fd_sc_hd__a221o_2 _15399_ (.A1(_02235_),
    .A2(_02237_),
    .B1(_02240_),
    .B2(_02017_),
    .C1(_01968_),
    .X(_02241_));
 sky130_fd_sc_hd__mux4_1 _15400_ (.A0(\cpuregs.regs[12][18] ),
    .A1(\cpuregs.regs[13][18] ),
    .A2(\cpuregs.regs[14][18] ),
    .A3(\cpuregs.regs[15][18] ),
    .S0(_03649_),
    .S1(_03643_),
    .X(_02242_));
 sky130_fd_sc_hd__mux4_1 _15401_ (.A0(\cpuregs.regs[8][18] ),
    .A1(\cpuregs.regs[9][18] ),
    .A2(\cpuregs.regs[10][18] ),
    .A3(\cpuregs.regs[11][18] ),
    .S0(_03645_),
    .S1(_01991_),
    .X(_02243_));
 sky130_fd_sc_hd__mux2_1 _15402_ (.A0(_02242_),
    .A1(_02243_),
    .S(_03719_),
    .X(_02244_));
 sky130_fd_sc_hd__mux4_1 _15403_ (.A0(\cpuregs.regs[28][18] ),
    .A1(\cpuregs.regs[29][18] ),
    .A2(\cpuregs.regs[30][18] ),
    .A3(\cpuregs.regs[31][18] ),
    .S0(_03661_),
    .S1(_03662_),
    .X(_02245_));
 sky130_fd_sc_hd__mux4_1 _15404_ (.A0(\cpuregs.regs[24][18] ),
    .A1(\cpuregs.regs[25][18] ),
    .A2(\cpuregs.regs[26][18] ),
    .A3(\cpuregs.regs[27][18] ),
    .S0(_03640_),
    .S1(_03642_),
    .X(_02246_));
 sky130_fd_sc_hd__mux2_1 _15405_ (.A0(_02245_),
    .A1(_02246_),
    .S(_03713_),
    .X(_02247_));
 sky130_fd_sc_hd__a21o_1 _15406_ (.A1(_03692_),
    .A2(_02247_),
    .B1(_03657_),
    .X(_02248_));
 sky130_fd_sc_hd__a21o_1 _15407_ (.A1(_02004_),
    .A2(_02244_),
    .B1(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__a32o_2 _15408_ (.A1(_01959_),
    .A2(_02241_),
    .A3(_02249_),
    .B1(_01933_),
    .B2(\decoded_imm[18] ),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _15409_ (.A0(net108),
    .A1(_02250_),
    .S(_01905_),
    .X(_02251_));
 sky130_fd_sc_hd__clkbuf_1 _15410_ (.A(_02251_),
    .X(_01171_));
 sky130_fd_sc_hd__mux4_1 _15411_ (.A0(\cpuregs.regs[4][19] ),
    .A1(\cpuregs.regs[5][19] ),
    .A2(\cpuregs.regs[6][19] ),
    .A3(\cpuregs.regs[7][19] ),
    .S0(_03670_),
    .S1(_03671_),
    .X(_02252_));
 sky130_fd_sc_hd__mux4_1 _15412_ (.A0(\cpuregs.regs[0][19] ),
    .A1(\cpuregs.regs[1][19] ),
    .A2(\cpuregs.regs[2][19] ),
    .A3(\cpuregs.regs[3][19] ),
    .S0(_03670_),
    .S1(_03671_),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _15413_ (.A0(_02252_),
    .A1(_02253_),
    .S(_03664_),
    .X(_02254_));
 sky130_fd_sc_hd__mux4_1 _15414_ (.A0(\cpuregs.regs[12][19] ),
    .A1(\cpuregs.regs[13][19] ),
    .A2(\cpuregs.regs[14][19] ),
    .A3(\cpuregs.regs[15][19] ),
    .S0(_01936_),
    .S1(_03647_),
    .X(_02255_));
 sky130_fd_sc_hd__o21a_1 _15415_ (.A1(_03719_),
    .A2(_02255_),
    .B1(_00067_),
    .X(_02256_));
 sky130_fd_sc_hd__mux4_1 _15416_ (.A0(\cpuregs.regs[8][19] ),
    .A1(\cpuregs.regs[9][19] ),
    .A2(\cpuregs.regs[10][19] ),
    .A3(\cpuregs.regs[11][19] ),
    .S0(_02046_),
    .S1(_02047_),
    .X(_02257_));
 sky130_fd_sc_hd__or2_1 _15417_ (.A(_03666_),
    .B(_02257_),
    .X(_02258_));
 sky130_fd_sc_hd__a221o_2 _15418_ (.A1(_02005_),
    .A2(_02254_),
    .B1(_02256_),
    .B2(_02258_),
    .C1(_03692_),
    .X(_02259_));
 sky130_fd_sc_hd__mux4_1 _15419_ (.A0(\cpuregs.regs[20][19] ),
    .A1(\cpuregs.regs[21][19] ),
    .A2(\cpuregs.regs[22][19] ),
    .A3(\cpuregs.regs[23][19] ),
    .S0(_03649_),
    .S1(_01991_),
    .X(_02260_));
 sky130_fd_sc_hd__mux4_1 _15420_ (.A0(\cpuregs.regs[16][19] ),
    .A1(\cpuregs.regs[17][19] ),
    .A2(\cpuregs.regs[18][19] ),
    .A3(\cpuregs.regs[19][19] ),
    .S0(_03645_),
    .S1(_01991_),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _15421_ (.A0(_02260_),
    .A1(_02261_),
    .S(_03653_),
    .X(_02262_));
 sky130_fd_sc_hd__mux4_1 _15422_ (.A0(\cpuregs.regs[28][19] ),
    .A1(\cpuregs.regs[29][19] ),
    .A2(\cpuregs.regs[30][19] ),
    .A3(\cpuregs.regs[31][19] ),
    .S0(_03661_),
    .S1(_03662_),
    .X(_02263_));
 sky130_fd_sc_hd__mux4_1 _15423_ (.A0(\cpuregs.regs[24][19] ),
    .A1(\cpuregs.regs[25][19] ),
    .A2(\cpuregs.regs[26][19] ),
    .A3(\cpuregs.regs[27][19] ),
    .S0(_03640_),
    .S1(_03642_),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _15424_ (.A0(_02263_),
    .A1(_02264_),
    .S(_03713_),
    .X(_02265_));
 sky130_fd_sc_hd__a21o_1 _15425_ (.A1(_03654_),
    .A2(_02265_),
    .B1(_03675_),
    .X(_02266_));
 sky130_fd_sc_hd__a21o_1 _15426_ (.A1(_02005_),
    .A2(_02262_),
    .B1(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__a32o_2 _15427_ (.A1(_01959_),
    .A2(_02259_),
    .A3(_02267_),
    .B1(_01933_),
    .B2(\decoded_imm[19] ),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _15428_ (.A0(net109),
    .A1(_02268_),
    .S(_01905_),
    .X(_02269_));
 sky130_fd_sc_hd__clkbuf_1 _15429_ (.A(_02269_),
    .X(_01172_));
 sky130_fd_sc_hd__mux4_1 _15430_ (.A0(\cpuregs.regs[12][20] ),
    .A1(\cpuregs.regs[13][20] ),
    .A2(\cpuregs.regs[14][20] ),
    .A3(\cpuregs.regs[15][20] ),
    .S0(_01979_),
    .S1(_01980_),
    .X(_02270_));
 sky130_fd_sc_hd__mux4_1 _15431_ (.A0(\cpuregs.regs[8][20] ),
    .A1(\cpuregs.regs[9][20] ),
    .A2(\cpuregs.regs[10][20] ),
    .A3(\cpuregs.regs[11][20] ),
    .S0(_02030_),
    .S1(_02031_),
    .X(_02271_));
 sky130_fd_sc_hd__mux4_1 _15432_ (.A0(\cpuregs.regs[4][20] ),
    .A1(\cpuregs.regs[5][20] ),
    .A2(\cpuregs.regs[6][20] ),
    .A3(\cpuregs.regs[7][20] ),
    .S0(_01976_),
    .S1(_01977_),
    .X(_02272_));
 sky130_fd_sc_hd__mux4_1 _15433_ (.A0(\cpuregs.regs[0][20] ),
    .A1(\cpuregs.regs[1][20] ),
    .A2(\cpuregs.regs[2][20] ),
    .A3(\cpuregs.regs[3][20] ),
    .S0(_02085_),
    .S1(_02086_),
    .X(_02273_));
 sky130_fd_sc_hd__mux4_1 _15434_ (.A0(_02270_),
    .A1(_02271_),
    .A2(_02272_),
    .A3(_02273_),
    .S0(_02111_),
    .S1(_02088_),
    .X(_02274_));
 sky130_fd_sc_hd__mux4_1 _15435_ (.A0(\cpuregs.regs[20][20] ),
    .A1(\cpuregs.regs[21][20] ),
    .A2(\cpuregs.regs[22][20] ),
    .A3(\cpuregs.regs[23][20] ),
    .S0(_01918_),
    .S1(_01919_),
    .X(_02275_));
 sky130_fd_sc_hd__mux4_1 _15436_ (.A0(\cpuregs.regs[16][20] ),
    .A1(\cpuregs.regs[17][20] ),
    .A2(\cpuregs.regs[18][20] ),
    .A3(\cpuregs.regs[19][20] ),
    .S0(_01918_),
    .S1(_01919_),
    .X(_02276_));
 sky130_fd_sc_hd__mux2_1 _15437_ (.A0(_02275_),
    .A1(_02276_),
    .S(_01907_),
    .X(_02277_));
 sky130_fd_sc_hd__mux4_1 _15438_ (.A0(\cpuregs.regs[28][20] ),
    .A1(\cpuregs.regs[29][20] ),
    .A2(\cpuregs.regs[30][20] ),
    .A3(\cpuregs.regs[31][20] ),
    .S0(_02030_),
    .S1(_02031_),
    .X(_02278_));
 sky130_fd_sc_hd__o21a_1 _15439_ (.A1(_02111_),
    .A2(_02278_),
    .B1(_01968_),
    .X(_02279_));
 sky130_fd_sc_hd__mux4_1 _15440_ (.A0(\cpuregs.regs[24][20] ),
    .A1(\cpuregs.regs[25][20] ),
    .A2(\cpuregs.regs[26][20] ),
    .A3(\cpuregs.regs[27][20] ),
    .S0(_01996_),
    .S1(_01997_),
    .X(_02280_));
 sky130_fd_sc_hd__or2_1 _15441_ (.A(_03687_),
    .B(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__a221o_1 _15442_ (.A1(_02088_),
    .A2(_02277_),
    .B1(_02279_),
    .B2(_02281_),
    .C1(_02018_),
    .X(_02282_));
 sky130_fd_sc_hd__o211a_2 _15443_ (.A1(_02020_),
    .A2(_02274_),
    .B1(_02282_),
    .C1(_01960_),
    .X(_02283_));
 sky130_fd_sc_hd__a21o_1 _15444_ (.A1(\decoded_imm[20] ),
    .A2(_02216_),
    .B1(_02197_),
    .X(_02284_));
 sky130_fd_sc_hd__o22a_1 _15445_ (.A1(net111),
    .A2(_02081_),
    .B1(_02283_),
    .B2(_02284_),
    .X(_01173_));
 sky130_fd_sc_hd__mux4_1 _15446_ (.A0(\cpuregs.regs[4][21] ),
    .A1(\cpuregs.regs[5][21] ),
    .A2(\cpuregs.regs[6][21] ),
    .A3(\cpuregs.regs[7][21] ),
    .S0(_01979_),
    .S1(_01980_),
    .X(_02285_));
 sky130_fd_sc_hd__mux4_1 _15447_ (.A0(\cpuregs.regs[0][21] ),
    .A1(\cpuregs.regs[1][21] ),
    .A2(\cpuregs.regs[2][21] ),
    .A3(\cpuregs.regs[3][21] ),
    .S0(_02030_),
    .S1(_02031_),
    .X(_02286_));
 sky130_fd_sc_hd__mux4_1 _15448_ (.A0(\cpuregs.regs[12][21] ),
    .A1(\cpuregs.regs[13][21] ),
    .A2(\cpuregs.regs[14][21] ),
    .A3(\cpuregs.regs[15][21] ),
    .S0(_01976_),
    .S1(_01977_),
    .X(_02287_));
 sky130_fd_sc_hd__mux4_1 _15449_ (.A0(\cpuregs.regs[8][21] ),
    .A1(\cpuregs.regs[9][21] ),
    .A2(\cpuregs.regs[10][21] ),
    .A3(\cpuregs.regs[11][21] ),
    .S0(_02085_),
    .S1(_02086_),
    .X(_02288_));
 sky130_fd_sc_hd__mux4_1 _15450_ (.A0(_02285_),
    .A1(_02286_),
    .A2(_02287_),
    .A3(_02288_),
    .S0(_02111_),
    .S1(_03683_),
    .X(_02289_));
 sky130_fd_sc_hd__mux4_1 _15451_ (.A0(\cpuregs.regs[16][21] ),
    .A1(\cpuregs.regs[17][21] ),
    .A2(\cpuregs.regs[18][21] ),
    .A3(\cpuregs.regs[19][21] ),
    .S0(_01996_),
    .S1(_01997_),
    .X(_02290_));
 sky130_fd_sc_hd__or2_1 _15452_ (.A(_02066_),
    .B(_02290_),
    .X(_02291_));
 sky130_fd_sc_hd__mux4_1 _15453_ (.A0(\cpuregs.regs[20][21] ),
    .A1(\cpuregs.regs[21][21] ),
    .A2(\cpuregs.regs[22][21] ),
    .A3(\cpuregs.regs[23][21] ),
    .S0(_02069_),
    .S1(_02070_),
    .X(_02292_));
 sky130_fd_sc_hd__o21a_1 _15454_ (.A1(_02012_),
    .A2(_02292_),
    .B1(_02005_),
    .X(_02293_));
 sky130_fd_sc_hd__mux4_1 _15455_ (.A0(\cpuregs.regs[28][21] ),
    .A1(\cpuregs.regs[29][21] ),
    .A2(\cpuregs.regs[30][21] ),
    .A3(\cpuregs.regs[31][21] ),
    .S0(_01999_),
    .S1(_02000_),
    .X(_02294_));
 sky130_fd_sc_hd__mux4_1 _15456_ (.A0(\cpuregs.regs[24][21] ),
    .A1(\cpuregs.regs[25][21] ),
    .A2(\cpuregs.regs[26][21] ),
    .A3(\cpuregs.regs[27][21] ),
    .S0(_02074_),
    .S1(_02075_),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _15457_ (.A0(_02294_),
    .A1(_02295_),
    .S(_01907_),
    .X(_02296_));
 sky130_fd_sc_hd__a221o_1 _15458_ (.A1(_02291_),
    .A2(_02293_),
    .B1(_02296_),
    .B2(_03683_),
    .C1(_02004_),
    .X(_02297_));
 sky130_fd_sc_hd__o211a_2 _15459_ (.A1(_02020_),
    .A2(_02289_),
    .B1(_02297_),
    .C1(_01960_),
    .X(_02298_));
 sky130_fd_sc_hd__a21o_1 _15460_ (.A1(\decoded_imm[21] ),
    .A2(_02216_),
    .B1(_02197_),
    .X(_02299_));
 sky130_fd_sc_hd__o22a_1 _15461_ (.A1(net112),
    .A2(_02081_),
    .B1(_02298_),
    .B2(_02299_),
    .X(_01174_));
 sky130_fd_sc_hd__mux4_1 _15462_ (.A0(\cpuregs.regs[20][22] ),
    .A1(\cpuregs.regs[21][22] ),
    .A2(\cpuregs.regs[22][22] ),
    .A3(\cpuregs.regs[23][22] ),
    .S0(_01979_),
    .S1(_01980_),
    .X(_02300_));
 sky130_fd_sc_hd__mux4_1 _15463_ (.A0(\cpuregs.regs[16][22] ),
    .A1(\cpuregs.regs[17][22] ),
    .A2(\cpuregs.regs[18][22] ),
    .A3(\cpuregs.regs[19][22] ),
    .S0(_02030_),
    .S1(_02031_),
    .X(_02301_));
 sky130_fd_sc_hd__mux4_1 _15464_ (.A0(\cpuregs.regs[4][22] ),
    .A1(\cpuregs.regs[5][22] ),
    .A2(\cpuregs.regs[6][22] ),
    .A3(\cpuregs.regs[7][22] ),
    .S0(_01973_),
    .S1(_01974_),
    .X(_02302_));
 sky130_fd_sc_hd__mux4_1 _15465_ (.A0(\cpuregs.regs[0][22] ),
    .A1(\cpuregs.regs[1][22] ),
    .A2(\cpuregs.regs[2][22] ),
    .A3(\cpuregs.regs[3][22] ),
    .S0(_02085_),
    .S1(_02086_),
    .X(_02303_));
 sky130_fd_sc_hd__mux4_1 _15466_ (.A0(_02300_),
    .A1(_02301_),
    .A2(_02302_),
    .A3(_02303_),
    .S0(_02111_),
    .S1(_02004_),
    .X(_02304_));
 sky130_fd_sc_hd__mux4_1 _15467_ (.A0(\cpuregs.regs[28][22] ),
    .A1(\cpuregs.regs[29][22] ),
    .A2(\cpuregs.regs[30][22] ),
    .A3(\cpuregs.regs[31][22] ),
    .S0(_01996_),
    .S1(_01997_),
    .X(_02305_));
 sky130_fd_sc_hd__or2_1 _15468_ (.A(_01984_),
    .B(_02305_),
    .X(_02306_));
 sky130_fd_sc_hd__mux4_1 _15469_ (.A0(\cpuregs.regs[24][22] ),
    .A1(\cpuregs.regs[25][22] ),
    .A2(\cpuregs.regs[26][22] ),
    .A3(\cpuregs.regs[27][22] ),
    .S0(_02069_),
    .S1(_02070_),
    .X(_02307_));
 sky130_fd_sc_hd__o21a_1 _15470_ (.A1(_02066_),
    .A2(_02307_),
    .B1(_03692_),
    .X(_02308_));
 sky130_fd_sc_hd__mux4_1 _15471_ (.A0(\cpuregs.regs[8][22] ),
    .A1(\cpuregs.regs[9][22] ),
    .A2(\cpuregs.regs[10][22] ),
    .A3(\cpuregs.regs[11][22] ),
    .S0(_01999_),
    .S1(_02000_),
    .X(_02309_));
 sky130_fd_sc_hd__mux4_1 _15472_ (.A0(\cpuregs.regs[12][22] ),
    .A1(\cpuregs.regs[13][22] ),
    .A2(\cpuregs.regs[14][22] ),
    .A3(\cpuregs.regs[15][22] ),
    .S0(_02074_),
    .S1(_02075_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _15473_ (.A0(_02309_),
    .A1(_02310_),
    .S(_03687_),
    .X(_02311_));
 sky130_fd_sc_hd__a221o_1 _15474_ (.A1(_02306_),
    .A2(_02308_),
    .B1(_02311_),
    .B2(_02004_),
    .C1(_02006_),
    .X(_02312_));
 sky130_fd_sc_hd__o211a_4 _15475_ (.A1(_01969_),
    .A2(_02304_),
    .B1(_02312_),
    .C1(_02027_),
    .X(_02313_));
 sky130_fd_sc_hd__a21o_1 _15476_ (.A1(\decoded_imm[22] ),
    .A2(_02216_),
    .B1(_02197_),
    .X(_02314_));
 sky130_fd_sc_hd__o22a_1 _15477_ (.A1(net113),
    .A2(_01905_),
    .B1(_02313_),
    .B2(_02314_),
    .X(_01175_));
 sky130_fd_sc_hd__mux4_1 _15478_ (.A0(\cpuregs.regs[0][23] ),
    .A1(\cpuregs.regs[1][23] ),
    .A2(\cpuregs.regs[2][23] ),
    .A3(\cpuregs.regs[3][23] ),
    .S0(_01995_),
    .S1(_01937_),
    .X(_02315_));
 sky130_fd_sc_hd__or2_1 _15479_ (.A(_03709_),
    .B(_02315_),
    .X(_02316_));
 sky130_fd_sc_hd__mux4_1 _15480_ (.A0(\cpuregs.regs[4][23] ),
    .A1(\cpuregs.regs[5][23] ),
    .A2(\cpuregs.regs[6][23] ),
    .A3(\cpuregs.regs[7][23] ),
    .S0(_01995_),
    .S1(_01937_),
    .X(_02317_));
 sky130_fd_sc_hd__o21a_1 _15481_ (.A1(_03719_),
    .A2(_02317_),
    .B1(_03674_),
    .X(_02318_));
 sky130_fd_sc_hd__mux4_1 _15482_ (.A0(\cpuregs.regs[20][23] ),
    .A1(\cpuregs.regs[21][23] ),
    .A2(\cpuregs.regs[22][23] ),
    .A3(\cpuregs.regs[23][23] ),
    .S0(_02046_),
    .S1(_02047_),
    .X(_02319_));
 sky130_fd_sc_hd__mux4_1 _15483_ (.A0(\cpuregs.regs[16][23] ),
    .A1(\cpuregs.regs[17][23] ),
    .A2(\cpuregs.regs[18][23] ),
    .A3(\cpuregs.regs[19][23] ),
    .S0(_02046_),
    .S1(_02047_),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _15484_ (.A0(_02319_),
    .A1(_02320_),
    .S(_03653_),
    .X(_02321_));
 sky130_fd_sc_hd__a221o_1 _15485_ (.A1(_02316_),
    .A2(_02318_),
    .B1(_02321_),
    .B2(_03692_),
    .C1(_01968_),
    .X(_02322_));
 sky130_fd_sc_hd__mux4_1 _15486_ (.A0(\cpuregs.regs[28][23] ),
    .A1(\cpuregs.regs[29][23] ),
    .A2(\cpuregs.regs[30][23] ),
    .A3(\cpuregs.regs[31][23] ),
    .S0(_03645_),
    .S1(_01991_),
    .X(_02323_));
 sky130_fd_sc_hd__mux4_1 _15487_ (.A0(\cpuregs.regs[24][23] ),
    .A1(\cpuregs.regs[25][23] ),
    .A2(\cpuregs.regs[26][23] ),
    .A3(\cpuregs.regs[27][23] ),
    .S0(_03645_),
    .S1(_01991_),
    .X(_02324_));
 sky130_fd_sc_hd__mux2_1 _15488_ (.A0(_02323_),
    .A1(_02324_),
    .S(_03653_),
    .X(_02325_));
 sky130_fd_sc_hd__mux4_1 _15489_ (.A0(\cpuregs.regs[12][23] ),
    .A1(\cpuregs.regs[13][23] ),
    .A2(\cpuregs.regs[14][23] ),
    .A3(\cpuregs.regs[15][23] ),
    .S0(_03661_),
    .S1(_03662_),
    .X(_02326_));
 sky130_fd_sc_hd__mux4_1 _15490_ (.A0(\cpuregs.regs[8][23] ),
    .A1(\cpuregs.regs[9][23] ),
    .A2(\cpuregs.regs[10][23] ),
    .A3(\cpuregs.regs[11][23] ),
    .S0(_03640_),
    .S1(_03642_),
    .X(_02327_));
 sky130_fd_sc_hd__mux2_1 _15491_ (.A0(_02326_),
    .A1(_02327_),
    .S(_03713_),
    .X(_02328_));
 sky130_fd_sc_hd__a21o_1 _15492_ (.A1(_03675_),
    .A2(_02328_),
    .B1(_03657_),
    .X(_02329_));
 sky130_fd_sc_hd__a21o_1 _15493_ (.A1(_03639_),
    .A2(_02325_),
    .B1(_02329_),
    .X(_02330_));
 sky130_fd_sc_hd__a32o_4 _15494_ (.A1(_01959_),
    .A2(_02322_),
    .A3(_02330_),
    .B1(_01933_),
    .B2(\decoded_imm[23] ),
    .X(_02331_));
 sky130_fd_sc_hd__mux2_1 _15495_ (.A0(net114),
    .A1(_02331_),
    .S(_03272_),
    .X(_02332_));
 sky130_fd_sc_hd__clkbuf_1 _15496_ (.A(_02332_),
    .X(_01176_));
 sky130_fd_sc_hd__mux4_1 _15497_ (.A0(\cpuregs.regs[12][24] ),
    .A1(\cpuregs.regs[13][24] ),
    .A2(\cpuregs.regs[14][24] ),
    .A3(\cpuregs.regs[15][24] ),
    .S0(_01970_),
    .S1(_01971_),
    .X(_02333_));
 sky130_fd_sc_hd__mux4_1 _15498_ (.A0(\cpuregs.regs[8][24] ),
    .A1(\cpuregs.regs[9][24] ),
    .A2(\cpuregs.regs[10][24] ),
    .A3(\cpuregs.regs[11][24] ),
    .S0(_02013_),
    .S1(_02014_),
    .X(_02334_));
 sky130_fd_sc_hd__or2_1 _15499_ (.A(_01989_),
    .B(_02334_),
    .X(_02335_));
 sky130_fd_sc_hd__o211a_1 _15500_ (.A1(_01982_),
    .A2(_02333_),
    .B1(_02335_),
    .C1(_02018_),
    .X(_02336_));
 sky130_fd_sc_hd__mux4_1 _15501_ (.A0(\cpuregs.regs[28][24] ),
    .A1(\cpuregs.regs[29][24] ),
    .A2(\cpuregs.regs[30][24] ),
    .A3(\cpuregs.regs[31][24] ),
    .S0(_01990_),
    .S1(_01992_),
    .X(_02337_));
 sky130_fd_sc_hd__mux4_1 _15502_ (.A0(\cpuregs.regs[24][24] ),
    .A1(\cpuregs.regs[25][24] ),
    .A2(\cpuregs.regs[26][24] ),
    .A3(\cpuregs.regs[27][24] ),
    .S0(_02022_),
    .S1(_02023_),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _15503_ (.A0(_02337_),
    .A1(_02338_),
    .S(_01984_),
    .X(_02339_));
 sky130_fd_sc_hd__a21o_1 _15504_ (.A1(_02037_),
    .A2(_02339_),
    .B1(_02006_),
    .X(_02340_));
 sky130_fd_sc_hd__mux4_1 _15505_ (.A0(\cpuregs.regs[4][24] ),
    .A1(\cpuregs.regs[5][24] ),
    .A2(\cpuregs.regs[6][24] ),
    .A3(\cpuregs.regs[7][24] ),
    .S0(_01990_),
    .S1(_01992_),
    .X(_02341_));
 sky130_fd_sc_hd__or2_1 _15506_ (.A(_01984_),
    .B(_02341_),
    .X(_02342_));
 sky130_fd_sc_hd__mux4_1 _15507_ (.A0(\cpuregs.regs[0][24] ),
    .A1(\cpuregs.regs[1][24] ),
    .A2(\cpuregs.regs[2][24] ),
    .A3(\cpuregs.regs[3][24] ),
    .S0(_02013_),
    .S1(_02014_),
    .X(_02343_));
 sky130_fd_sc_hd__o21a_1 _15508_ (.A1(_01989_),
    .A2(_02343_),
    .B1(_02017_),
    .X(_02344_));
 sky130_fd_sc_hd__mux4_1 _15509_ (.A0(\cpuregs.regs[20][24] ),
    .A1(\cpuregs.regs[21][24] ),
    .A2(\cpuregs.regs[22][24] ),
    .A3(\cpuregs.regs[23][24] ),
    .S0(_02022_),
    .S1(_02023_),
    .X(_02345_));
 sky130_fd_sc_hd__mux4_1 _15510_ (.A0(\cpuregs.regs[16][24] ),
    .A1(\cpuregs.regs[17][24] ),
    .A2(\cpuregs.regs[18][24] ),
    .A3(\cpuregs.regs[19][24] ),
    .S0(_01985_),
    .S1(_01986_),
    .X(_02346_));
 sky130_fd_sc_hd__mux2_1 _15511_ (.A0(_02345_),
    .A1(_02346_),
    .S(_02002_),
    .X(_02347_));
 sky130_fd_sc_hd__a221o_1 _15512_ (.A1(_02342_),
    .A2(_02344_),
    .B1(_02347_),
    .B2(_02037_),
    .C1(_01969_),
    .X(_02348_));
 sky130_fd_sc_hd__o211a_2 _15513_ (.A1(_02336_),
    .A2(_02340_),
    .B1(_02027_),
    .C1(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__a21o_1 _15514_ (.A1(\decoded_imm[24] ),
    .A2(_02216_),
    .B1(_02197_),
    .X(_02350_));
 sky130_fd_sc_hd__o22a_1 _15515_ (.A1(net115),
    .A2(_01905_),
    .B1(_02349_),
    .B2(_02350_),
    .X(_01177_));
 sky130_fd_sc_hd__mux4_1 _15516_ (.A0(\cpuregs.regs[4][25] ),
    .A1(\cpuregs.regs[5][25] ),
    .A2(\cpuregs.regs[6][25] ),
    .A3(\cpuregs.regs[7][25] ),
    .S0(_01979_),
    .S1(_01980_),
    .X(_02351_));
 sky130_fd_sc_hd__mux4_1 _15517_ (.A0(\cpuregs.regs[0][25] ),
    .A1(\cpuregs.regs[1][25] ),
    .A2(\cpuregs.regs[2][25] ),
    .A3(\cpuregs.regs[3][25] ),
    .S0(_02030_),
    .S1(_02031_),
    .X(_02352_));
 sky130_fd_sc_hd__mux4_1 _15518_ (.A0(\cpuregs.regs[20][25] ),
    .A1(\cpuregs.regs[21][25] ),
    .A2(\cpuregs.regs[22][25] ),
    .A3(\cpuregs.regs[23][25] ),
    .S0(_01973_),
    .S1(_01974_),
    .X(_02353_));
 sky130_fd_sc_hd__mux4_1 _15519_ (.A0(\cpuregs.regs[16][25] ),
    .A1(\cpuregs.regs[17][25] ),
    .A2(\cpuregs.regs[18][25] ),
    .A3(\cpuregs.regs[19][25] ),
    .S0(_02085_),
    .S1(_02086_),
    .X(_02354_));
 sky130_fd_sc_hd__mux4_1 _15520_ (.A0(_02351_),
    .A1(_02352_),
    .A2(_02353_),
    .A3(_02354_),
    .S0(_02111_),
    .S1(_03639_),
    .X(_02355_));
 sky130_fd_sc_hd__mux4_1 _15521_ (.A0(\cpuregs.regs[8][25] ),
    .A1(\cpuregs.regs[9][25] ),
    .A2(\cpuregs.regs[10][25] ),
    .A3(\cpuregs.regs[11][25] ),
    .S0(_01996_),
    .S1(_01997_),
    .X(_02356_));
 sky130_fd_sc_hd__or2_1 _15522_ (.A(_03687_),
    .B(_02356_),
    .X(_02357_));
 sky130_fd_sc_hd__mux4_1 _15523_ (.A0(\cpuregs.regs[12][25] ),
    .A1(\cpuregs.regs[13][25] ),
    .A2(\cpuregs.regs[14][25] ),
    .A3(\cpuregs.regs[15][25] ),
    .S0(_02069_),
    .S1(_02070_),
    .X(_02358_));
 sky130_fd_sc_hd__o21a_1 _15524_ (.A1(_02012_),
    .A2(_02358_),
    .B1(_02017_),
    .X(_02359_));
 sky130_fd_sc_hd__mux4_1 _15525_ (.A0(\cpuregs.regs[28][25] ),
    .A1(\cpuregs.regs[29][25] ),
    .A2(\cpuregs.regs[30][25] ),
    .A3(\cpuregs.regs[31][25] ),
    .S0(_01999_),
    .S1(_02000_),
    .X(_02360_));
 sky130_fd_sc_hd__mux4_1 _15526_ (.A0(\cpuregs.regs[24][25] ),
    .A1(\cpuregs.regs[25][25] ),
    .A2(\cpuregs.regs[26][25] ),
    .A3(\cpuregs.regs[27][25] ),
    .S0(_02074_),
    .S1(_02075_),
    .X(_02361_));
 sky130_fd_sc_hd__mux2_1 _15527_ (.A0(_02360_),
    .A1(_02361_),
    .S(_01907_),
    .X(_02362_));
 sky130_fd_sc_hd__a221o_1 _15528_ (.A1(_02357_),
    .A2(_02359_),
    .B1(_02362_),
    .B2(_02037_),
    .C1(_02006_),
    .X(_02363_));
 sky130_fd_sc_hd__o211a_2 _15529_ (.A1(_01969_),
    .A2(_02355_),
    .B1(_02363_),
    .C1(_02027_),
    .X(_02364_));
 sky130_fd_sc_hd__a21o_1 _15530_ (.A1(\decoded_imm[25] ),
    .A2(_02216_),
    .B1(_02197_),
    .X(_02365_));
 sky130_fd_sc_hd__o22a_1 _15531_ (.A1(net116),
    .A2(_01905_),
    .B1(_02364_),
    .B2(_02365_),
    .X(_01178_));
 sky130_fd_sc_hd__mux4_1 _15532_ (.A0(\cpuregs.regs[16][26] ),
    .A1(\cpuregs.regs[17][26] ),
    .A2(\cpuregs.regs[18][26] ),
    .A3(\cpuregs.regs[19][26] ),
    .S0(_01995_),
    .S1(_01937_),
    .X(_02366_));
 sky130_fd_sc_hd__or2_1 _15533_ (.A(_03709_),
    .B(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__mux4_1 _15534_ (.A0(\cpuregs.regs[20][26] ),
    .A1(\cpuregs.regs[21][26] ),
    .A2(\cpuregs.regs[22][26] ),
    .A3(\cpuregs.regs[23][26] ),
    .S0(_01995_),
    .S1(_01937_),
    .X(_02368_));
 sky130_fd_sc_hd__o21a_1 _15535_ (.A1(_03719_),
    .A2(_02368_),
    .B1(_00068_),
    .X(_02369_));
 sky130_fd_sc_hd__mux4_1 _15536_ (.A0(\cpuregs.regs[4][26] ),
    .A1(\cpuregs.regs[5][26] ),
    .A2(\cpuregs.regs[6][26] ),
    .A3(\cpuregs.regs[7][26] ),
    .S0(_02046_),
    .S1(_02047_),
    .X(_02370_));
 sky130_fd_sc_hd__mux4_1 _15537_ (.A0(\cpuregs.regs[0][26] ),
    .A1(\cpuregs.regs[1][26] ),
    .A2(\cpuregs.regs[2][26] ),
    .A3(\cpuregs.regs[3][26] ),
    .S0(_02046_),
    .S1(_02047_),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _15538_ (.A0(_02370_),
    .A1(_02371_),
    .S(_03653_),
    .X(_02372_));
 sky130_fd_sc_hd__a221o_1 _15539_ (.A1(_02367_),
    .A2(_02369_),
    .B1(_02372_),
    .B2(_02017_),
    .C1(_01968_),
    .X(_02373_));
 sky130_fd_sc_hd__mux4_1 _15540_ (.A0(\cpuregs.regs[24][26] ),
    .A1(\cpuregs.regs[25][26] ),
    .A2(\cpuregs.regs[26][26] ),
    .A3(\cpuregs.regs[27][26] ),
    .S0(_03645_),
    .S1(_01991_),
    .X(_02374_));
 sky130_fd_sc_hd__mux4_1 _15541_ (.A0(\cpuregs.regs[28][26] ),
    .A1(\cpuregs.regs[29][26] ),
    .A2(\cpuregs.regs[30][26] ),
    .A3(\cpuregs.regs[31][26] ),
    .S0(_03645_),
    .S1(_03647_),
    .X(_02375_));
 sky130_fd_sc_hd__mux2_1 _15542_ (.A0(_02374_),
    .A1(_02375_),
    .S(_03709_),
    .X(_02376_));
 sky130_fd_sc_hd__mux4_1 _15543_ (.A0(\cpuregs.regs[12][26] ),
    .A1(\cpuregs.regs[13][26] ),
    .A2(\cpuregs.regs[14][26] ),
    .A3(\cpuregs.regs[15][26] ),
    .S0(_03661_),
    .S1(_03642_),
    .X(_02377_));
 sky130_fd_sc_hd__mux4_1 _15544_ (.A0(\cpuregs.regs[8][26] ),
    .A1(\cpuregs.regs[9][26] ),
    .A2(\cpuregs.regs[10][26] ),
    .A3(\cpuregs.regs[11][26] ),
    .S0(_03640_),
    .S1(_03642_),
    .X(_02378_));
 sky130_fd_sc_hd__mux2_1 _15545_ (.A0(_02377_),
    .A1(_02378_),
    .S(_03713_),
    .X(_02379_));
 sky130_fd_sc_hd__a21o_1 _15546_ (.A1(_03675_),
    .A2(_02379_),
    .B1(_03657_),
    .X(_02380_));
 sky130_fd_sc_hd__a21o_1 _15547_ (.A1(_03639_),
    .A2(_02376_),
    .B1(_02380_),
    .X(_02381_));
 sky130_fd_sc_hd__a32o_2 _15548_ (.A1(_01959_),
    .A2(_02373_),
    .A3(_02381_),
    .B1(_01933_),
    .B2(\decoded_imm[26] ),
    .X(_02382_));
 sky130_fd_sc_hd__mux2_1 _15549_ (.A0(net117),
    .A1(_02382_),
    .S(_03272_),
    .X(_02383_));
 sky130_fd_sc_hd__clkbuf_1 _15550_ (.A(_02383_),
    .X(_01179_));
 sky130_fd_sc_hd__mux4_1 _15551_ (.A0(\cpuregs.regs[20][27] ),
    .A1(\cpuregs.regs[21][27] ),
    .A2(\cpuregs.regs[22][27] ),
    .A3(\cpuregs.regs[23][27] ),
    .S0(_01979_),
    .S1(_01980_),
    .X(_02384_));
 sky130_fd_sc_hd__mux4_1 _15552_ (.A0(\cpuregs.regs[16][27] ),
    .A1(\cpuregs.regs[17][27] ),
    .A2(\cpuregs.regs[18][27] ),
    .A3(\cpuregs.regs[19][27] ),
    .S0(_02030_),
    .S1(_02031_),
    .X(_02385_));
 sky130_fd_sc_hd__mux4_1 _15553_ (.A0(\cpuregs.regs[4][27] ),
    .A1(\cpuregs.regs[5][27] ),
    .A2(\cpuregs.regs[6][27] ),
    .A3(\cpuregs.regs[7][27] ),
    .S0(_01973_),
    .S1(_01974_),
    .X(_02386_));
 sky130_fd_sc_hd__mux4_1 _15554_ (.A0(\cpuregs.regs[0][27] ),
    .A1(\cpuregs.regs[1][27] ),
    .A2(\cpuregs.regs[2][27] ),
    .A3(\cpuregs.regs[3][27] ),
    .S0(_02085_),
    .S1(_02086_),
    .X(_02387_));
 sky130_fd_sc_hd__mux4_1 _15555_ (.A0(_02384_),
    .A1(_02385_),
    .A2(_02386_),
    .A3(_02387_),
    .S0(_02111_),
    .S1(_02004_),
    .X(_02388_));
 sky130_fd_sc_hd__mux4_1 _15556_ (.A0(\cpuregs.regs[28][27] ),
    .A1(\cpuregs.regs[29][27] ),
    .A2(\cpuregs.regs[30][27] ),
    .A3(\cpuregs.regs[31][27] ),
    .S0(_01996_),
    .S1(_01997_),
    .X(_02389_));
 sky130_fd_sc_hd__or2_1 _15557_ (.A(_01984_),
    .B(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__mux4_1 _15558_ (.A0(\cpuregs.regs[24][27] ),
    .A1(\cpuregs.regs[25][27] ),
    .A2(\cpuregs.regs[26][27] ),
    .A3(\cpuregs.regs[27][27] ),
    .S0(_02069_),
    .S1(_02070_),
    .X(_02391_));
 sky130_fd_sc_hd__o21a_1 _15559_ (.A1(_02066_),
    .A2(_02391_),
    .B1(_03692_),
    .X(_02392_));
 sky130_fd_sc_hd__mux4_1 _15560_ (.A0(\cpuregs.regs[12][27] ),
    .A1(\cpuregs.regs[13][27] ),
    .A2(\cpuregs.regs[14][27] ),
    .A3(\cpuregs.regs[15][27] ),
    .S0(_01999_),
    .S1(_02000_),
    .X(_02393_));
 sky130_fd_sc_hd__mux4_1 _15561_ (.A0(\cpuregs.regs[8][27] ),
    .A1(\cpuregs.regs[9][27] ),
    .A2(\cpuregs.regs[10][27] ),
    .A3(\cpuregs.regs[11][27] ),
    .S0(_02074_),
    .S1(_02075_),
    .X(_02394_));
 sky130_fd_sc_hd__mux2_1 _15562_ (.A0(_02393_),
    .A1(_02394_),
    .S(_01907_),
    .X(_02395_));
 sky130_fd_sc_hd__a221o_1 _15563_ (.A1(_02390_),
    .A2(_02392_),
    .B1(_02395_),
    .B2(_02004_),
    .C1(_02088_),
    .X(_02396_));
 sky130_fd_sc_hd__o211a_2 _15564_ (.A1(_01969_),
    .A2(_02388_),
    .B1(_02396_),
    .C1(_02027_),
    .X(_02397_));
 sky130_fd_sc_hd__a21o_1 _15565_ (.A1(\decoded_imm[27] ),
    .A2(_02216_),
    .B1(_02197_),
    .X(_02398_));
 sky130_fd_sc_hd__o22a_1 _15566_ (.A1(net118),
    .A2(_01905_),
    .B1(_02397_),
    .B2(_02398_),
    .X(_01180_));
 sky130_fd_sc_hd__mux4_1 _15567_ (.A0(\cpuregs.regs[12][28] ),
    .A1(\cpuregs.regs[13][28] ),
    .A2(\cpuregs.regs[14][28] ),
    .A3(\cpuregs.regs[15][28] ),
    .S0(_01979_),
    .S1(_01980_),
    .X(_02399_));
 sky130_fd_sc_hd__mux4_1 _15568_ (.A0(\cpuregs.regs[8][28] ),
    .A1(\cpuregs.regs[9][28] ),
    .A2(\cpuregs.regs[10][28] ),
    .A3(\cpuregs.regs[11][28] ),
    .S0(_02030_),
    .S1(_02031_),
    .X(_02400_));
 sky130_fd_sc_hd__mux4_1 _15569_ (.A0(\cpuregs.regs[4][28] ),
    .A1(\cpuregs.regs[5][28] ),
    .A2(\cpuregs.regs[6][28] ),
    .A3(\cpuregs.regs[7][28] ),
    .S0(_01973_),
    .S1(_01974_),
    .X(_02401_));
 sky130_fd_sc_hd__mux4_1 _15570_ (.A0(\cpuregs.regs[0][28] ),
    .A1(\cpuregs.regs[1][28] ),
    .A2(\cpuregs.regs[2][28] ),
    .A3(\cpuregs.regs[3][28] ),
    .S0(_01976_),
    .S1(_01977_),
    .X(_02402_));
 sky130_fd_sc_hd__mux4_1 _15571_ (.A0(_02399_),
    .A1(_02400_),
    .A2(_02401_),
    .A3(_02402_),
    .S0(_02111_),
    .S1(_02005_),
    .X(_02403_));
 sky130_fd_sc_hd__mux4_1 _15572_ (.A0(\cpuregs.regs[16][28] ),
    .A1(\cpuregs.regs[17][28] ),
    .A2(\cpuregs.regs[18][28] ),
    .A3(\cpuregs.regs[19][28] ),
    .S0(_01918_),
    .S1(_01919_),
    .X(_02404_));
 sky130_fd_sc_hd__mux4_1 _15573_ (.A0(\cpuregs.regs[20][28] ),
    .A1(\cpuregs.regs[21][28] ),
    .A2(\cpuregs.regs[22][28] ),
    .A3(\cpuregs.regs[23][28] ),
    .S0(_01918_),
    .S1(_01919_),
    .X(_02405_));
 sky130_fd_sc_hd__mux2_1 _15574_ (.A0(_02404_),
    .A1(_02405_),
    .S(_03687_),
    .X(_02406_));
 sky130_fd_sc_hd__mux4_1 _15575_ (.A0(\cpuregs.regs[28][28] ),
    .A1(\cpuregs.regs[29][28] ),
    .A2(\cpuregs.regs[30][28] ),
    .A3(\cpuregs.regs[31][28] ),
    .S0(_02030_),
    .S1(_02031_),
    .X(_02407_));
 sky130_fd_sc_hd__o21a_1 _15576_ (.A1(_02111_),
    .A2(_02407_),
    .B1(_01968_),
    .X(_02408_));
 sky130_fd_sc_hd__mux4_1 _15577_ (.A0(\cpuregs.regs[24][28] ),
    .A1(\cpuregs.regs[25][28] ),
    .A2(\cpuregs.regs[26][28] ),
    .A3(\cpuregs.regs[27][28] ),
    .S0(_01996_),
    .S1(_01997_),
    .X(_02409_));
 sky130_fd_sc_hd__or2_1 _15578_ (.A(_03687_),
    .B(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__a221o_1 _15579_ (.A1(_02088_),
    .A2(_02406_),
    .B1(_02408_),
    .B2(_02410_),
    .C1(_02004_),
    .X(_02411_));
 sky130_fd_sc_hd__o211a_2 _15580_ (.A1(_02020_),
    .A2(_02403_),
    .B1(_02411_),
    .C1(_02027_),
    .X(_02412_));
 sky130_fd_sc_hd__a21o_1 _15581_ (.A1(\decoded_imm[28] ),
    .A2(_02216_),
    .B1(_02197_),
    .X(_02413_));
 sky130_fd_sc_hd__o22a_1 _15582_ (.A1(net119),
    .A2(_01905_),
    .B1(_02412_),
    .B2(_02413_),
    .X(_01181_));
 sky130_fd_sc_hd__mux4_1 _15583_ (.A0(\cpuregs.regs[4][29] ),
    .A1(\cpuregs.regs[5][29] ),
    .A2(\cpuregs.regs[6][29] ),
    .A3(\cpuregs.regs[7][29] ),
    .S0(_01908_),
    .S1(_01909_),
    .X(_02414_));
 sky130_fd_sc_hd__mux4_1 _15584_ (.A0(\cpuregs.regs[0][29] ),
    .A1(\cpuregs.regs[1][29] ),
    .A2(\cpuregs.regs[2][29] ),
    .A3(\cpuregs.regs[3][29] ),
    .S0(_01908_),
    .S1(_01909_),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _15585_ (.A0(_02414_),
    .A1(_02415_),
    .S(_01907_),
    .X(_02416_));
 sky130_fd_sc_hd__mux4_1 _15586_ (.A0(\cpuregs.regs[12][29] ),
    .A1(\cpuregs.regs[13][29] ),
    .A2(\cpuregs.regs[14][29] ),
    .A3(\cpuregs.regs[15][29] ),
    .S0(_03641_),
    .S1(_03684_),
    .X(_02417_));
 sky130_fd_sc_hd__mux4_1 _15587_ (.A0(\cpuregs.regs[8][29] ),
    .A1(\cpuregs.regs[9][29] ),
    .A2(\cpuregs.regs[10][29] ),
    .A3(\cpuregs.regs[11][29] ),
    .S0(_03641_),
    .S1(_03684_),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _15588_ (.A0(_02417_),
    .A1(_02418_),
    .S(_02110_),
    .X(_02419_));
 sky130_fd_sc_hd__mux4_1 _15589_ (.A0(\cpuregs.regs[20][29] ),
    .A1(\cpuregs.regs[21][29] ),
    .A2(\cpuregs.regs[22][29] ),
    .A3(\cpuregs.regs[23][29] ),
    .S0(_02221_),
    .S1(_02222_),
    .X(_02420_));
 sky130_fd_sc_hd__mux4_1 _15590_ (.A0(\cpuregs.regs[16][29] ),
    .A1(\cpuregs.regs[17][29] ),
    .A2(\cpuregs.regs[18][29] ),
    .A3(\cpuregs.regs[19][29] ),
    .S0(_02221_),
    .S1(_02222_),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _15591_ (.A0(_02420_),
    .A1(_02421_),
    .S(_02110_),
    .X(_02422_));
 sky130_fd_sc_hd__mux4_1 _15592_ (.A0(\cpuregs.regs[28][29] ),
    .A1(\cpuregs.regs[29][29] ),
    .A2(\cpuregs.regs[30][29] ),
    .A3(\cpuregs.regs[31][29] ),
    .S0(_01908_),
    .S1(_01909_),
    .X(_02423_));
 sky130_fd_sc_hd__mux4_1 _15593_ (.A0(\cpuregs.regs[24][29] ),
    .A1(\cpuregs.regs[25][29] ),
    .A2(\cpuregs.regs[26][29] ),
    .A3(\cpuregs.regs[27][29] ),
    .S0(_02221_),
    .S1(_02222_),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _15594_ (.A0(_02423_),
    .A1(_02424_),
    .S(_02110_),
    .X(_02425_));
 sky130_fd_sc_hd__mux4_2 _15595_ (.A0(_02416_),
    .A1(_02419_),
    .A2(_02422_),
    .A3(_02425_),
    .S0(_01968_),
    .S1(_02037_),
    .X(_02426_));
 sky130_fd_sc_hd__a221o_2 _15596_ (.A1(\decoded_imm[29] ),
    .A2(_02216_),
    .B1(_01959_),
    .B2(_02426_),
    .C1(_01934_),
    .X(_02427_));
 sky130_fd_sc_hd__o21a_1 _15597_ (.A1(net120),
    .A2(_01906_),
    .B1(_02427_),
    .X(_01182_));
 sky130_fd_sc_hd__mux4_1 _15598_ (.A0(\cpuregs.regs[4][30] ),
    .A1(\cpuregs.regs[5][30] ),
    .A2(\cpuregs.regs[6][30] ),
    .A3(\cpuregs.regs[7][30] ),
    .S0(_01908_),
    .S1(_01909_),
    .X(_02428_));
 sky130_fd_sc_hd__mux4_1 _15599_ (.A0(\cpuregs.regs[0][30] ),
    .A1(\cpuregs.regs[1][30] ),
    .A2(\cpuregs.regs[2][30] ),
    .A3(\cpuregs.regs[3][30] ),
    .S0(_01908_),
    .S1(_01909_),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _15600_ (.A0(_02428_),
    .A1(_02429_),
    .S(_01907_),
    .X(_02430_));
 sky130_fd_sc_hd__mux4_1 _15601_ (.A0(\cpuregs.regs[12][30] ),
    .A1(\cpuregs.regs[13][30] ),
    .A2(\cpuregs.regs[14][30] ),
    .A3(\cpuregs.regs[15][30] ),
    .S0(_03641_),
    .S1(_03684_),
    .X(_02431_));
 sky130_fd_sc_hd__mux4_1 _15602_ (.A0(\cpuregs.regs[8][30] ),
    .A1(\cpuregs.regs[9][30] ),
    .A2(\cpuregs.regs[10][30] ),
    .A3(\cpuregs.regs[11][30] ),
    .S0(_03641_),
    .S1(_03684_),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _15603_ (.A0(_02431_),
    .A1(_02432_),
    .S(_02110_),
    .X(_02433_));
 sky130_fd_sc_hd__mux4_1 _15604_ (.A0(\cpuregs.regs[20][30] ),
    .A1(\cpuregs.regs[21][30] ),
    .A2(\cpuregs.regs[22][30] ),
    .A3(\cpuregs.regs[23][30] ),
    .S0(_02221_),
    .S1(_02222_),
    .X(_02434_));
 sky130_fd_sc_hd__mux4_1 _15605_ (.A0(\cpuregs.regs[16][30] ),
    .A1(\cpuregs.regs[17][30] ),
    .A2(\cpuregs.regs[18][30] ),
    .A3(\cpuregs.regs[19][30] ),
    .S0(_02221_),
    .S1(_02222_),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _15606_ (.A0(_02434_),
    .A1(_02435_),
    .S(_02110_),
    .X(_02436_));
 sky130_fd_sc_hd__mux4_1 _15607_ (.A0(\cpuregs.regs[28][30] ),
    .A1(\cpuregs.regs[29][30] ),
    .A2(\cpuregs.regs[30][30] ),
    .A3(\cpuregs.regs[31][30] ),
    .S0(_01908_),
    .S1(_01909_),
    .X(_02437_));
 sky130_fd_sc_hd__mux4_1 _15608_ (.A0(\cpuregs.regs[24][30] ),
    .A1(\cpuregs.regs[25][30] ),
    .A2(\cpuregs.regs[26][30] ),
    .A3(\cpuregs.regs[27][30] ),
    .S0(_02221_),
    .S1(_02222_),
    .X(_02438_));
 sky130_fd_sc_hd__mux2_1 _15609_ (.A0(_02437_),
    .A1(_02438_),
    .S(_02110_),
    .X(_02439_));
 sky130_fd_sc_hd__mux4_2 _15610_ (.A0(_02430_),
    .A1(_02433_),
    .A2(_02436_),
    .A3(_02439_),
    .S0(_01968_),
    .S1(_03639_),
    .X(_02440_));
 sky130_fd_sc_hd__a221o_4 _15611_ (.A1(\decoded_imm[30] ),
    .A2(_01933_),
    .B1(_01959_),
    .B2(_02440_),
    .C1(_01934_),
    .X(_02441_));
 sky130_fd_sc_hd__o21a_1 _15612_ (.A1(net122),
    .A2(_01906_),
    .B1(_02441_),
    .X(_01183_));
 sky130_fd_sc_hd__mux4_1 _15613_ (.A0(\cpuregs.regs[16][31] ),
    .A1(\cpuregs.regs[17][31] ),
    .A2(\cpuregs.regs[18][31] ),
    .A3(\cpuregs.regs[19][31] ),
    .S0(_01995_),
    .S1(_01937_),
    .X(_02442_));
 sky130_fd_sc_hd__or2_1 _15614_ (.A(_03709_),
    .B(_02442_),
    .X(_02443_));
 sky130_fd_sc_hd__mux4_1 _15615_ (.A0(\cpuregs.regs[20][31] ),
    .A1(\cpuregs.regs[21][31] ),
    .A2(\cpuregs.regs[22][31] ),
    .A3(\cpuregs.regs[23][31] ),
    .S0(_01995_),
    .S1(_01937_),
    .X(_02444_));
 sky130_fd_sc_hd__o21a_1 _15616_ (.A1(_03719_),
    .A2(_02444_),
    .B1(_00068_),
    .X(_02445_));
 sky130_fd_sc_hd__mux4_1 _15617_ (.A0(\cpuregs.regs[4][31] ),
    .A1(\cpuregs.regs[5][31] ),
    .A2(\cpuregs.regs[6][31] ),
    .A3(\cpuregs.regs[7][31] ),
    .S0(_02046_),
    .S1(_02047_),
    .X(_02446_));
 sky130_fd_sc_hd__mux4_1 _15618_ (.A0(\cpuregs.regs[0][31] ),
    .A1(\cpuregs.regs[1][31] ),
    .A2(\cpuregs.regs[2][31] ),
    .A3(\cpuregs.regs[3][31] ),
    .S0(_02046_),
    .S1(_02047_),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _15619_ (.A0(_02446_),
    .A1(_02447_),
    .S(_03653_),
    .X(_02448_));
 sky130_fd_sc_hd__a221o_2 _15620_ (.A1(_02443_),
    .A2(_02445_),
    .B1(_02448_),
    .B2(_03675_),
    .C1(_03654_),
    .X(_02449_));
 sky130_fd_sc_hd__mux4_1 _15621_ (.A0(\cpuregs.regs[8][31] ),
    .A1(\cpuregs.regs[9][31] ),
    .A2(\cpuregs.regs[10][31] ),
    .A3(\cpuregs.regs[11][31] ),
    .S0(_03645_),
    .S1(_01991_),
    .X(_02450_));
 sky130_fd_sc_hd__mux4_1 _15622_ (.A0(\cpuregs.regs[12][31] ),
    .A1(\cpuregs.regs[13][31] ),
    .A2(\cpuregs.regs[14][31] ),
    .A3(\cpuregs.regs[15][31] ),
    .S0(_03645_),
    .S1(_03647_),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _15623_ (.A0(_02450_),
    .A1(_02451_),
    .S(_03709_),
    .X(_02452_));
 sky130_fd_sc_hd__mux4_1 _15624_ (.A0(\cpuregs.regs[24][31] ),
    .A1(\cpuregs.regs[25][31] ),
    .A2(\cpuregs.regs[26][31] ),
    .A3(\cpuregs.regs[27][31] ),
    .S0(_03640_),
    .S1(_03642_),
    .X(_02453_));
 sky130_fd_sc_hd__mux4_1 _15625_ (.A0(\cpuregs.regs[28][31] ),
    .A1(\cpuregs.regs[29][31] ),
    .A2(\cpuregs.regs[30][31] ),
    .A3(\cpuregs.regs[31][31] ),
    .S0(_03640_),
    .S1(_03642_),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _15626_ (.A0(_02453_),
    .A1(_02454_),
    .S(_03666_),
    .X(_02455_));
 sky130_fd_sc_hd__a21o_1 _15627_ (.A1(_00068_),
    .A2(_02455_),
    .B1(_03657_),
    .X(_02456_));
 sky130_fd_sc_hd__a21o_1 _15628_ (.A1(_02017_),
    .A2(_02452_),
    .B1(_02456_),
    .X(_02457_));
 sky130_fd_sc_hd__a32o_2 _15629_ (.A1(_01959_),
    .A2(_02449_),
    .A3(_02457_),
    .B1(_01932_),
    .B2(\decoded_imm[31] ),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _15630_ (.A0(net123),
    .A1(_02458_),
    .S(_03272_),
    .X(_02459_));
 sky130_fd_sc_hd__clkbuf_1 _15631_ (.A(_02459_),
    .X(_01184_));
 sky130_fd_sc_hd__nor2_1 _15632_ (.A(_04271_),
    .B(instr_jalr),
    .Y(_02460_));
 sky130_fd_sc_hd__mux2_1 _15633_ (.A0(_02460_),
    .A1(mem_do_prefetch),
    .S(_03380_),
    .X(_02461_));
 sky130_fd_sc_hd__and3_1 _15634_ (.A(_07778_),
    .B(_03237_),
    .C(_02461_),
    .X(_02462_));
 sky130_fd_sc_hd__clkbuf_1 _15635_ (.A(_02462_),
    .X(_01185_));
 sky130_fd_sc_hd__nand2_1 _15636_ (.A(\cpu_state[2] ),
    .B(_03254_),
    .Y(_02463_));
 sky130_fd_sc_hd__o211a_1 _15637_ (.A1(_03298_),
    .A2(_03410_),
    .B1(_03400_),
    .C1(_03277_),
    .X(_02464_));
 sky130_fd_sc_hd__and3_1 _15638_ (.A(_02463_),
    .B(_03307_),
    .C(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__o21ba_1 _15639_ (.A1(decoder_trigger),
    .A2(do_waitirq),
    .B1_N(\irq_state[0] ),
    .X(_02466_));
 sky130_fd_sc_hd__o21a_1 _15640_ (.A1(_03379_),
    .A2(_07994_),
    .B1(_03364_),
    .X(_02467_));
 sky130_fd_sc_hd__a211oi_1 _15641_ (.A1(_07992_),
    .A2(_02466_),
    .B1(_02467_),
    .C1(_03410_),
    .Y(_02468_));
 sky130_fd_sc_hd__a22o_1 _15642_ (.A1(is_lb_lh_lw_lbu_lhu),
    .A2(_03270_),
    .B1(_03396_),
    .B2(is_sb_sh_sw),
    .X(_02469_));
 sky130_fd_sc_hd__a22o_1 _15643_ (.A1(mem_do_prefetch),
    .A2(_03410_),
    .B1(_02469_),
    .B2(_03301_),
    .X(_02470_));
 sky130_fd_sc_hd__or3b_1 _15644_ (.A(_02468_),
    .B(_02470_),
    .C_N(_02465_),
    .X(_02471_));
 sky130_fd_sc_hd__nor2_1 _15645_ (.A(_03239_),
    .B(_03310_),
    .Y(_02472_));
 sky130_fd_sc_hd__o211a_1 _15646_ (.A1(_03199_),
    .A2(_02465_),
    .B1(_02471_),
    .C1(_02472_),
    .X(_02473_));
 sky130_fd_sc_hd__a41o_1 _15647_ (.A1(_03309_),
    .A2(_03411_),
    .A3(_03630_),
    .A4(_07905_),
    .B1(_02473_),
    .X(_01186_));
 sky130_fd_sc_hd__a21o_1 _15648_ (.A1(_03218_),
    .A2(_02472_),
    .B1(_03291_),
    .X(_01187_));
 sky130_fd_sc_hd__or4b_1 _15649_ (.A(mem_do_wdata),
    .B(_03278_),
    .C(_04006_),
    .D_N(_07904_),
    .X(_02474_));
 sky130_fd_sc_hd__a2bb2o_1 _15650_ (.A1_N(\cpu_state[0] ),
    .A2_N(_02474_),
    .B1(_02472_),
    .B2(mem_do_wdata),
    .X(_01188_));
 sky130_fd_sc_hd__and2_1 _15651_ (.A(_03301_),
    .B(_04187_),
    .X(_02475_));
 sky130_fd_sc_hd__buf_2 _15652_ (.A(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__clkbuf_4 _15653_ (.A(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__nor2_1 _15654_ (.A(\timer[0] ),
    .B(_03427_),
    .Y(_02478_));
 sky130_fd_sc_hd__clkbuf_4 _15655_ (.A(_02475_),
    .X(_02479_));
 sky130_fd_sc_hd__nand2_1 _15656_ (.A(_07208_),
    .B(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__clkbuf_4 _15657_ (.A(_07778_),
    .X(_02481_));
 sky130_fd_sc_hd__o211a_1 _15658_ (.A1(_02477_),
    .A2(_02478_),
    .B1(_02480_),
    .C1(_02481_),
    .X(_01189_));
 sky130_fd_sc_hd__inv_2 _15659_ (.A(\timer[1] ),
    .Y(_02482_));
 sky130_fd_sc_hd__nand2_1 _15660_ (.A(_02482_),
    .B(_02478_),
    .Y(_02483_));
 sky130_fd_sc_hd__nand2_2 _15661_ (.A(_03301_),
    .B(_04024_),
    .Y(_02484_));
 sky130_fd_sc_hd__o21a_1 _15662_ (.A1(_02482_),
    .A2(_02478_),
    .B1(_02484_),
    .X(_02485_));
 sky130_fd_sc_hd__a221oi_1 _15663_ (.A1(_04101_),
    .A2(_02477_),
    .B1(_02483_),
    .B2(_02485_),
    .C1(_07775_),
    .Y(_01190_));
 sky130_fd_sc_hd__clkbuf_4 _15664_ (.A(_02484_),
    .X(_02486_));
 sky130_fd_sc_hd__nor2_1 _15665_ (.A(\timer[2] ),
    .B(_02483_),
    .Y(_02487_));
 sky130_fd_sc_hd__clkbuf_4 _15666_ (.A(_02475_),
    .X(_02488_));
 sky130_fd_sc_hd__a21o_1 _15667_ (.A1(\timer[2] ),
    .A2(_02483_),
    .B1(_02488_),
    .X(_02489_));
 sky130_fd_sc_hd__o221a_1 _15668_ (.A1(_07250_),
    .A2(_02486_),
    .B1(_02487_),
    .B2(_02489_),
    .C1(_06026_),
    .X(_01191_));
 sky130_fd_sc_hd__or3_1 _15669_ (.A(\timer[3] ),
    .B(\timer[2] ),
    .C(_02483_),
    .X(_02490_));
 sky130_fd_sc_hd__o21ai_1 _15670_ (.A1(\timer[2] ),
    .A2(_02483_),
    .B1(\timer[3] ),
    .Y(_02491_));
 sky130_fd_sc_hd__a31o_1 _15671_ (.A1(_02484_),
    .A2(_02490_),
    .A3(_02491_),
    .B1(_03240_),
    .X(_02492_));
 sky130_fd_sc_hd__a21oi_1 _15672_ (.A1(_04185_),
    .A2(_02477_),
    .B1(_02492_),
    .Y(_01192_));
 sky130_fd_sc_hd__or2_1 _15673_ (.A(\timer[4] ),
    .B(_02490_),
    .X(_02493_));
 sky130_fd_sc_hd__a21oi_1 _15674_ (.A1(\timer[4] ),
    .A2(_02490_),
    .B1(_02488_),
    .Y(_02494_));
 sky130_fd_sc_hd__a221oi_1 _15675_ (.A1(_04240_),
    .A2(_02477_),
    .B1(_02493_),
    .B2(_02494_),
    .C1(_07775_),
    .Y(_01193_));
 sky130_fd_sc_hd__or2_1 _15676_ (.A(\timer[5] ),
    .B(_02493_),
    .X(_02495_));
 sky130_fd_sc_hd__a21oi_1 _15677_ (.A1(\timer[5] ),
    .A2(_02493_),
    .B1(_02488_),
    .Y(_02496_));
 sky130_fd_sc_hd__a221oi_1 _15678_ (.A1(_01872_),
    .A2(_02479_),
    .B1(_02495_),
    .B2(_02496_),
    .C1(_07775_),
    .Y(_01194_));
 sky130_fd_sc_hd__xnor2_1 _15679_ (.A(\timer[6] ),
    .B(_02495_),
    .Y(_02497_));
 sky130_fd_sc_hd__nand2_1 _15680_ (.A(_04335_),
    .B(_02479_),
    .Y(_02498_));
 sky130_fd_sc_hd__o211a_1 _15681_ (.A1(_02477_),
    .A2(_02497_),
    .B1(_02498_),
    .C1(_02481_),
    .X(_01195_));
 sky130_fd_sc_hd__o21a_1 _15682_ (.A1(\timer[6] ),
    .A2(_02495_),
    .B1(\timer[7] ),
    .X(_02499_));
 sky130_fd_sc_hd__or3_2 _15683_ (.A(\timer[0] ),
    .B(_03416_),
    .C(_03427_),
    .X(_02500_));
 sky130_fd_sc_hd__inv_2 _15684_ (.A(_02500_),
    .Y(_02501_));
 sky130_fd_sc_hd__nand2_1 _15685_ (.A(_04382_),
    .B(_02479_),
    .Y(_02502_));
 sky130_fd_sc_hd__o311a_1 _15686_ (.A1(_02477_),
    .A2(_02499_),
    .A3(_02501_),
    .B1(_02502_),
    .C1(_06026_),
    .X(_01196_));
 sky130_fd_sc_hd__or2_1 _15687_ (.A(\timer[0] ),
    .B(_03416_),
    .X(_02503_));
 sky130_fd_sc_hd__a21o_1 _15688_ (.A1(\timer[8] ),
    .A2(_02503_),
    .B1(_02476_),
    .X(_02504_));
 sky130_fd_sc_hd__nor2_1 _15689_ (.A(\timer[8] ),
    .B(_02500_),
    .Y(_02505_));
 sky130_fd_sc_hd__o221a_1 _15690_ (.A1(_04415_),
    .A2(_02486_),
    .B1(_02504_),
    .B2(_02505_),
    .C1(_06026_),
    .X(_01197_));
 sky130_fd_sc_hd__clkbuf_4 _15691_ (.A(_02486_),
    .X(_02506_));
 sky130_fd_sc_hd__o21ai_1 _15692_ (.A1(\timer[8] ),
    .A2(_02503_),
    .B1(\timer[9] ),
    .Y(_02507_));
 sky130_fd_sc_hd__or3_2 _15693_ (.A(\timer[9] ),
    .B(\timer[8] ),
    .C(_02500_),
    .X(_02508_));
 sky130_fd_sc_hd__a31o_1 _15694_ (.A1(_02484_),
    .A2(_02507_),
    .A3(_02508_),
    .B1(_03240_),
    .X(_02509_));
 sky130_fd_sc_hd__o21ba_1 _15695_ (.A1(_04447_),
    .A2(_02506_),
    .B1_N(_02509_),
    .X(_01198_));
 sky130_fd_sc_hd__a21o_1 _15696_ (.A1(\timer[10] ),
    .A2(_02508_),
    .B1(_02476_),
    .X(_02510_));
 sky130_fd_sc_hd__nor2_1 _15697_ (.A(\timer[10] ),
    .B(_02508_),
    .Y(_02511_));
 sky130_fd_sc_hd__o221a_1 _15698_ (.A1(_07371_),
    .A2(_02486_),
    .B1(_02510_),
    .B2(_02511_),
    .C1(_06026_),
    .X(_01199_));
 sky130_fd_sc_hd__xor2_1 _15699_ (.A(\timer[11] ),
    .B(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__nand2_1 _15700_ (.A(_01881_),
    .B(_02479_),
    .Y(_02513_));
 sky130_fd_sc_hd__o211a_1 _15701_ (.A1(_02477_),
    .A2(_02512_),
    .B1(_02513_),
    .C1(_02481_),
    .X(_01200_));
 sky130_fd_sc_hd__or3_1 _15702_ (.A(\timer[11] ),
    .B(\timer[10] ),
    .C(_02508_),
    .X(_02514_));
 sky130_fd_sc_hd__a21oi_1 _15703_ (.A1(\timer[12] ),
    .A2(_02514_),
    .B1(_02475_),
    .Y(_02515_));
 sky130_fd_sc_hd__or2_1 _15704_ (.A(\timer[12] ),
    .B(_02514_),
    .X(_02516_));
 sky130_fd_sc_hd__a22o_1 _15705_ (.A1(_04561_),
    .A2(_02476_),
    .B1(_02515_),
    .B2(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__nor2_1 _15706_ (.A(_08335_),
    .B(_02517_),
    .Y(_01201_));
 sky130_fd_sc_hd__a21oi_1 _15707_ (.A1(\timer[13] ),
    .A2(_02516_),
    .B1(_02488_),
    .Y(_02518_));
 sky130_fd_sc_hd__o21ai_1 _15708_ (.A1(\timer[13] ),
    .A2(_02516_),
    .B1(_02518_),
    .Y(_02519_));
 sky130_fd_sc_hd__o211a_1 _15709_ (.A1(_04593_),
    .A2(_02506_),
    .B1(_02519_),
    .C1(_02481_),
    .X(_01202_));
 sky130_fd_sc_hd__o21ai_1 _15710_ (.A1(\timer[13] ),
    .A2(_02516_),
    .B1(\timer[14] ),
    .Y(_02520_));
 sky130_fd_sc_hd__or3_1 _15711_ (.A(\timer[13] ),
    .B(\timer[14] ),
    .C(_02516_),
    .X(_02521_));
 sky130_fd_sc_hd__and3_1 _15712_ (.A(_02484_),
    .B(_02520_),
    .C(_02521_),
    .X(_02522_));
 sky130_fd_sc_hd__a211oi_1 _15713_ (.A1(_04631_),
    .A2(_02477_),
    .B1(_02522_),
    .C1(_07775_),
    .Y(_01203_));
 sky130_fd_sc_hd__and2_1 _15714_ (.A(\timer[15] ),
    .B(_02521_),
    .X(_02523_));
 sky130_fd_sc_hd__or2_1 _15715_ (.A(\timer[15] ),
    .B(_02521_),
    .X(_02524_));
 sky130_fd_sc_hd__or3b_1 _15716_ (.A(_02476_),
    .B(_02523_),
    .C_N(_02524_),
    .X(_02525_));
 sky130_fd_sc_hd__o211a_1 _15717_ (.A1(_07441_),
    .A2(_02506_),
    .B1(_02525_),
    .C1(_02481_),
    .X(_01204_));
 sky130_fd_sc_hd__a21o_1 _15718_ (.A1(\timer[16] ),
    .A2(_02524_),
    .B1(_02488_),
    .X(_02526_));
 sky130_fd_sc_hd__nor2_1 _15719_ (.A(\timer[16] ),
    .B(_02524_),
    .Y(_02527_));
 sky130_fd_sc_hd__nand2_1 _15720_ (.A(_04702_),
    .B(_02479_),
    .Y(_02528_));
 sky130_fd_sc_hd__o211a_1 _15721_ (.A1(_02526_),
    .A2(_02527_),
    .B1(_02528_),
    .C1(_02481_),
    .X(_01205_));
 sky130_fd_sc_hd__o21a_1 _15722_ (.A1(\timer[16] ),
    .A2(_02524_),
    .B1(\timer[17] ),
    .X(_02529_));
 sky130_fd_sc_hd__and2b_1 _15723_ (.A_N(\timer[17] ),
    .B(_02527_),
    .X(_02530_));
 sky130_fd_sc_hd__nand2_1 _15724_ (.A(_04737_),
    .B(_02479_),
    .Y(_02531_));
 sky130_fd_sc_hd__o311a_1 _15725_ (.A1(_02477_),
    .A2(_02529_),
    .A3(_02530_),
    .B1(_02531_),
    .C1(_06026_),
    .X(_01206_));
 sky130_fd_sc_hd__and2b_1 _15726_ (.A_N(_02530_),
    .B(\timer[18] ),
    .X(_02532_));
 sky130_fd_sc_hd__or4_2 _15727_ (.A(\timer[17] ),
    .B(\timer[16] ),
    .C(\timer[18] ),
    .D(_02524_),
    .X(_02533_));
 sky130_fd_sc_hd__or3b_1 _15728_ (.A(_02476_),
    .B(_02532_),
    .C_N(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__o211a_1 _15729_ (.A1(_04777_),
    .A2(_02506_),
    .B1(_02534_),
    .C1(_02481_),
    .X(_01207_));
 sky130_fd_sc_hd__a21oi_1 _15730_ (.A1(\timer[19] ),
    .A2(_02533_),
    .B1(_02488_),
    .Y(_02535_));
 sky130_fd_sc_hd__o21ai_1 _15731_ (.A1(\timer[19] ),
    .A2(_02533_),
    .B1(_02535_),
    .Y(_02536_));
 sky130_fd_sc_hd__o211a_1 _15732_ (.A1(_04806_),
    .A2(_02506_),
    .B1(_02536_),
    .C1(_02481_),
    .X(_01208_));
 sky130_fd_sc_hd__o21a_1 _15733_ (.A1(\timer[19] ),
    .A2(_02533_),
    .B1(\timer[20] ),
    .X(_02537_));
 sky130_fd_sc_hd__or3_1 _15734_ (.A(\timer[19] ),
    .B(\timer[20] ),
    .C(_02533_),
    .X(_02538_));
 sky130_fd_sc_hd__or3b_1 _15735_ (.A(_02476_),
    .B(_02537_),
    .C_N(_02538_),
    .X(_02539_));
 sky130_fd_sc_hd__o211a_1 _15736_ (.A1(_04842_),
    .A2(_02506_),
    .B1(_02539_),
    .C1(_02481_),
    .X(_01209_));
 sky130_fd_sc_hd__or2_1 _15737_ (.A(\timer[21] ),
    .B(_02538_),
    .X(_02540_));
 sky130_fd_sc_hd__a21oi_1 _15738_ (.A1(\timer[21] ),
    .A2(_02538_),
    .B1(_02488_),
    .Y(_02541_));
 sky130_fd_sc_hd__nand2_1 _15739_ (.A(_02540_),
    .B(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__o211a_1 _15740_ (.A1(_04871_),
    .A2(_02506_),
    .B1(_02542_),
    .C1(_02481_),
    .X(_01210_));
 sky130_fd_sc_hd__a21oi_1 _15741_ (.A1(\timer[22] ),
    .A2(_02540_),
    .B1(_02488_),
    .Y(_02543_));
 sky130_fd_sc_hd__o21ai_1 _15742_ (.A1(\timer[22] ),
    .A2(_02540_),
    .B1(_02543_),
    .Y(_02544_));
 sky130_fd_sc_hd__buf_2 _15743_ (.A(_07778_),
    .X(_02545_));
 sky130_fd_sc_hd__o211a_1 _15744_ (.A1(_04909_),
    .A2(_02506_),
    .B1(_02544_),
    .C1(_02545_),
    .X(_01211_));
 sky130_fd_sc_hd__o21a_1 _15745_ (.A1(\timer[22] ),
    .A2(_02540_),
    .B1(\timer[23] ),
    .X(_02546_));
 sky130_fd_sc_hd__or3_2 _15746_ (.A(\timer[23] ),
    .B(\timer[22] ),
    .C(_02540_),
    .X(_02547_));
 sky130_fd_sc_hd__or3b_1 _15747_ (.A(_02476_),
    .B(_02546_),
    .C_N(_02547_),
    .X(_02548_));
 sky130_fd_sc_hd__o211a_1 _15748_ (.A1(_04941_),
    .A2(_02506_),
    .B1(_02548_),
    .C1(_02545_),
    .X(_01212_));
 sky130_fd_sc_hd__a21oi_1 _15749_ (.A1(\timer[24] ),
    .A2(_02547_),
    .B1(_02488_),
    .Y(_02549_));
 sky130_fd_sc_hd__o21ai_1 _15750_ (.A1(\timer[24] ),
    .A2(_02547_),
    .B1(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__o211a_1 _15751_ (.A1(_04979_),
    .A2(_02506_),
    .B1(_02550_),
    .C1(_02545_),
    .X(_01213_));
 sky130_fd_sc_hd__o21a_1 _15752_ (.A1(\timer[24] ),
    .A2(_02547_),
    .B1(\timer[25] ),
    .X(_02551_));
 sky130_fd_sc_hd__or3_1 _15753_ (.A(\timer[25] ),
    .B(\timer[24] ),
    .C(_02547_),
    .X(_02552_));
 sky130_fd_sc_hd__or3b_1 _15754_ (.A(_02476_),
    .B(_02551_),
    .C_N(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__o211a_1 _15755_ (.A1(_05009_),
    .A2(_02486_),
    .B1(_02553_),
    .C1(_02545_),
    .X(_01214_));
 sky130_fd_sc_hd__nor2_1 _15756_ (.A(\timer[26] ),
    .B(_02552_),
    .Y(_02554_));
 sky130_fd_sc_hd__a21o_1 _15757_ (.A1(\timer[26] ),
    .A2(_02552_),
    .B1(_02479_),
    .X(_02555_));
 sky130_fd_sc_hd__nand2_1 _15758_ (.A(_05037_),
    .B(_02479_),
    .Y(_02556_));
 sky130_fd_sc_hd__o211a_1 _15759_ (.A1(_02554_),
    .A2(_02555_),
    .B1(_02556_),
    .C1(_02545_),
    .X(_01215_));
 sky130_fd_sc_hd__inv_2 _15760_ (.A(\timer[27] ),
    .Y(_02557_));
 sky130_fd_sc_hd__o22ai_1 _15761_ (.A1(_03417_),
    .A2(_02547_),
    .B1(_02554_),
    .B2(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__nand2_1 _15762_ (.A(_05069_),
    .B(_02479_),
    .Y(_02559_));
 sky130_fd_sc_hd__o211a_1 _15763_ (.A1(_02477_),
    .A2(_02558_),
    .B1(_02559_),
    .C1(_02545_),
    .X(_01216_));
 sky130_fd_sc_hd__or2_2 _15764_ (.A(_03423_),
    .B(_02503_),
    .X(_02560_));
 sky130_fd_sc_hd__or3_1 _15765_ (.A(\timer[28] ),
    .B(_03425_),
    .C(_02560_),
    .X(_02561_));
 sky130_fd_sc_hd__inv_2 _15766_ (.A(_02561_),
    .Y(_02562_));
 sky130_fd_sc_hd__a211o_1 _15767_ (.A1(\timer[28] ),
    .A2(_02560_),
    .B1(_02562_),
    .C1(_02488_),
    .X(_02563_));
 sky130_fd_sc_hd__o211a_1 _15768_ (.A1(_05107_),
    .A2(_02486_),
    .B1(_02563_),
    .C1(_02545_),
    .X(_01217_));
 sky130_fd_sc_hd__or2_1 _15769_ (.A(\timer[29] ),
    .B(_02561_),
    .X(_02564_));
 sky130_fd_sc_hd__nand2_1 _15770_ (.A(_02484_),
    .B(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__a21o_1 _15771_ (.A1(\timer[29] ),
    .A2(_02561_),
    .B1(_02565_),
    .X(_02566_));
 sky130_fd_sc_hd__o211a_1 _15772_ (.A1(_05139_),
    .A2(_02486_),
    .B1(_02566_),
    .C1(_02545_),
    .X(_01218_));
 sky130_fd_sc_hd__nor2_1 _15773_ (.A(_03424_),
    .B(_02560_),
    .Y(_02567_));
 sky130_fd_sc_hd__a221o_1 _15774_ (.A1(\timer[31] ),
    .A2(_02567_),
    .B1(_02564_),
    .B2(\timer[30] ),
    .C1(_02476_),
    .X(_02568_));
 sky130_fd_sc_hd__o211a_1 _15775_ (.A1(_05170_),
    .A2(_02486_),
    .B1(_02568_),
    .C1(_02545_),
    .X(_01219_));
 sky130_fd_sc_hd__inv_2 _15776_ (.A(\timer[31] ),
    .Y(_02569_));
 sky130_fd_sc_hd__o21ai_1 _15777_ (.A1(_02569_),
    .A2(_02567_),
    .B1(_02486_),
    .Y(_02570_));
 sky130_fd_sc_hd__o211a_1 _15778_ (.A1(_05201_),
    .A2(_02486_),
    .B1(_02570_),
    .C1(_02545_),
    .X(_01220_));
 sky130_fd_sc_hd__a32o_1 _15779_ (.A1(_03376_),
    .A2(_07899_),
    .A3(_03363_),
    .B1(_07905_),
    .B2(_06186_),
    .X(_01221_));
 sky130_fd_sc_hd__a21o_1 _15780_ (.A1(_06186_),
    .A2(_03298_),
    .B1(_03409_),
    .X(_02571_));
 sky130_fd_sc_hd__and3_1 _15781_ (.A(_07778_),
    .B(_07676_),
    .C(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__clkbuf_1 _15782_ (.A(_02572_),
    .X(_01222_));
 sky130_fd_sc_hd__o21a_1 _15783_ (.A1(_03298_),
    .A2(_04006_),
    .B1(_03389_),
    .X(_02573_));
 sky130_fd_sc_hd__or2b_1 _15784_ (.A(_03630_),
    .B_N(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_02574_));
 sky130_fd_sc_hd__and3_1 _15785_ (.A(_03317_),
    .B(_03364_),
    .C(_07984_),
    .X(_02575_));
 sky130_fd_sc_hd__or3b_1 _15786_ (.A(_03410_),
    .B(_02575_),
    .C_N(_02573_),
    .X(_02576_));
 sky130_fd_sc_hd__a211o_1 _15787_ (.A1(_03384_),
    .A2(_02574_),
    .B1(_02576_),
    .C1(_03226_),
    .X(_02577_));
 sky130_fd_sc_hd__o211a_1 _15788_ (.A1(latched_store),
    .A2(_02573_),
    .B1(_02577_),
    .C1(_06026_),
    .X(_01223_));
 sky130_fd_sc_hd__o221a_1 _15789_ (.A1(_03385_),
    .A2(_03292_),
    .B1(_03318_),
    .B2(_06069_),
    .C1(_06026_),
    .X(_01224_));
 sky130_fd_sc_hd__a31oi_1 _15790_ (.A1(_04156_),
    .A2(_03292_),
    .A3(_03271_),
    .B1(_07680_),
    .Y(_02578_));
 sky130_fd_sc_hd__o211a_1 _15791_ (.A1(is_beq_bne_blt_bge_bltu_bgeu),
    .A2(instr_jalr),
    .B1(_02574_),
    .C1(\cpu_state[3] ),
    .X(_02579_));
 sky130_fd_sc_hd__and3_1 _15792_ (.A(_04156_),
    .B(_06863_),
    .C(_03368_),
    .X(_02580_));
 sky130_fd_sc_hd__or4b_1 _15793_ (.A(_03302_),
    .B(_02579_),
    .C(_02580_),
    .D_N(_02578_),
    .X(_02581_));
 sky130_fd_sc_hd__o211a_1 _15794_ (.A1(latched_branch),
    .A2(_02578_),
    .B1(_02581_),
    .C1(_06026_),
    .X(_01225_));
 sky130_fd_sc_hd__o211a_1 _15795_ (.A1(_03292_),
    .A2(_03226_),
    .B1(_03282_),
    .C1(_03305_),
    .X(_02582_));
 sky130_fd_sc_hd__a22o_1 _15796_ (.A1(instr_lh),
    .A2(_03291_),
    .B1(_02582_),
    .B2(latched_is_lh),
    .X(_01227_));
 sky130_fd_sc_hd__a22o_1 _15797_ (.A1(instr_lb),
    .A2(_03291_),
    .B1(_02582_),
    .B2(latched_is_lb),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _15798_ (.A0(latched_compr),
    .A1(compressed_instr),
    .S(_08033_),
    .X(_02583_));
 sky130_fd_sc_hd__clkbuf_1 _15799_ (.A(_02583_),
    .X(_01229_));
 sky130_fd_sc_hd__and2_1 _15800_ (.A(_08033_),
    .B(_07994_),
    .X(_02584_));
 sky130_fd_sc_hd__clkbuf_1 _15801_ (.A(_02584_),
    .X(_01230_));
 sky130_fd_sc_hd__a21o_1 _15802_ (.A1(\decoded_imm_j[1] ),
    .A2(_05974_),
    .B1(_05978_),
    .X(_01231_));
 sky130_fd_sc_hd__a21o_1 _15803_ (.A1(\decoded_imm_j[2] ),
    .A2(_05974_),
    .B1(_05982_),
    .X(_01232_));
 sky130_fd_sc_hd__a221o_1 _15804_ (.A1(\decoded_imm_j[3] ),
    .A2(_05983_),
    .B1(_03895_),
    .B2(_06016_),
    .C1(_05985_),
    .X(_01233_));
 sky130_fd_sc_hd__and2_1 _15805_ (.A(_05960_),
    .B(_03763_),
    .X(_02585_));
 sky130_fd_sc_hd__o22a_1 _15806_ (.A1(\decoded_imm_j[4] ),
    .A2(_06006_),
    .B1(_02585_),
    .B2(_05988_),
    .X(_01234_));
 sky130_fd_sc_hd__nor2_1 _15807_ (.A(_05960_),
    .B(_05970_),
    .Y(_02586_));
 sky130_fd_sc_hd__buf_2 _15808_ (.A(_02586_),
    .X(_02587_));
 sky130_fd_sc_hd__and3_1 _15809_ (.A(_05960_),
    .B(_03634_),
    .C(_03864_),
    .X(_02588_));
 sky130_fd_sc_hd__a221o_1 _15810_ (.A1(\decoded_imm_j[5] ),
    .A2(_05983_),
    .B1(_03954_),
    .B2(_02587_),
    .C1(_02588_),
    .X(_01235_));
 sky130_fd_sc_hd__and3_1 _15811_ (.A(_05960_),
    .B(_03634_),
    .C(_03822_),
    .X(_02589_));
 sky130_fd_sc_hd__a221o_1 _15812_ (.A1(\decoded_imm_j[6] ),
    .A2(_05983_),
    .B1(_03965_),
    .B2(_02587_),
    .C1(_02589_),
    .X(_01236_));
 sky130_fd_sc_hd__and3_1 _15813_ (.A(_05960_),
    .B(_03634_),
    .C(_03878_),
    .X(_02590_));
 sky130_fd_sc_hd__a221o_1 _15814_ (.A1(\decoded_imm_j[7] ),
    .A2(_05983_),
    .B1(_03977_),
    .B2(_02587_),
    .C1(_02590_),
    .X(_01237_));
 sky130_fd_sc_hd__and2_1 _15815_ (.A(\decoded_imm_j[8] ),
    .B(_05973_),
    .X(_02591_));
 sky130_fd_sc_hd__a221o_1 _15816_ (.A1(_03826_),
    .A2(_06016_),
    .B1(_02587_),
    .B2(_03987_),
    .C1(_02591_),
    .X(_01238_));
 sky130_fd_sc_hd__a22o_1 _15817_ (.A1(_03892_),
    .A2(_06016_),
    .B1(_02587_),
    .B2(_03994_),
    .X(_02592_));
 sky130_fd_sc_hd__a21o_1 _15818_ (.A1(\decoded_imm_j[9] ),
    .A2(_05974_),
    .B1(_02592_),
    .X(_01239_));
 sky130_fd_sc_hd__a22o_1 _15819_ (.A1(_03867_),
    .A2(_06016_),
    .B1(_02586_),
    .B2(_04000_),
    .X(_02593_));
 sky130_fd_sc_hd__a21o_1 _15820_ (.A1(\decoded_imm_j[10] ),
    .A2(_05974_),
    .B1(_02593_),
    .X(_01240_));
 sky130_fd_sc_hd__nand2_1 _15821_ (.A(_05960_),
    .B(_03737_),
    .Y(_02594_));
 sky130_fd_sc_hd__o2bb2a_1 _15822_ (.A1_N(_05971_),
    .A2_N(_02594_),
    .B1(\decoded_imm_j[11] ),
    .B2(_03636_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _15823_ (.A0(\decoded_imm_j[12] ),
    .A1(_03737_),
    .S(_03635_),
    .X(_02595_));
 sky130_fd_sc_hd__clkbuf_1 _15824_ (.A(_02595_),
    .X(_01242_));
 sky130_fd_sc_hd__nor2_2 _15825_ (.A(_05970_),
    .B(_02594_),
    .Y(_02596_));
 sky130_fd_sc_hd__a221o_1 _15826_ (.A1(\decoded_imm_j[13] ),
    .A2(_05983_),
    .B1(_03747_),
    .B2(_02587_),
    .C1(_02596_),
    .X(_01243_));
 sky130_fd_sc_hd__a221o_1 _15827_ (.A1(\decoded_imm_j[14] ),
    .A2(_05987_),
    .B1(_03891_),
    .B2(_02587_),
    .C1(_02596_),
    .X(_01244_));
 sky130_fd_sc_hd__a221o_1 _15828_ (.A1(\decoded_imm_j[15] ),
    .A2(_05987_),
    .B1(_03781_),
    .B2(_02587_),
    .C1(_02596_),
    .X(_01245_));
 sky130_fd_sc_hd__a221o_1 _15829_ (.A1(\decoded_imm_j[16] ),
    .A2(_05987_),
    .B1(_03910_),
    .B2(_02587_),
    .C1(_02596_),
    .X(_01246_));
 sky130_fd_sc_hd__nor2_1 _15830_ (.A(_05987_),
    .B(_06017_),
    .Y(_02597_));
 sky130_fd_sc_hd__a211o_1 _15831_ (.A1(\decoded_imm_j[17] ),
    .A2(_05983_),
    .B1(_02596_),
    .C1(_02597_),
    .X(_01247_));
 sky130_fd_sc_hd__and3_1 _15832_ (.A(_05969_),
    .B(_03634_),
    .C(_03918_),
    .X(_02598_));
 sky130_fd_sc_hd__a211o_1 _15833_ (.A1(\decoded_imm_j[18] ),
    .A2(_05983_),
    .B1(_02596_),
    .C1(_02598_),
    .X(_01248_));
 sky130_fd_sc_hd__and3_1 _15834_ (.A(_05969_),
    .B(_03634_),
    .C(_03920_),
    .X(_02599_));
 sky130_fd_sc_hd__a211o_1 _15835_ (.A1(\decoded_imm_j[19] ),
    .A2(_05983_),
    .B1(_02596_),
    .C1(_02599_),
    .X(_01249_));
 sky130_fd_sc_hd__a221o_1 _15836_ (.A1(_08232_),
    .A2(_05987_),
    .B1(_03756_),
    .B2(_02587_),
    .C1(_02596_),
    .X(_01250_));
 sky130_fd_sc_hd__nand2_1 _15837_ (.A(_03816_),
    .B(_03916_),
    .Y(_02600_));
 sky130_fd_sc_hd__and3_1 _15838_ (.A(_03739_),
    .B(_03869_),
    .C(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__and3b_1 _15839_ (.A_N(_03878_),
    .B(_03885_),
    .C(_03895_),
    .X(_02602_));
 sky130_fd_sc_hd__and3_1 _15840_ (.A(_03215_),
    .B(_03979_),
    .C(_03864_),
    .X(_02603_));
 sky130_fd_sc_hd__and3_1 _15841_ (.A(_03634_),
    .B(_02602_),
    .C(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__a221o_1 _15842_ (.A1(instr_lui),
    .A2(_05987_),
    .B1(_06016_),
    .B2(_02601_),
    .C1(_02604_),
    .X(_01251_));
 sky130_fd_sc_hd__and3_1 _15843_ (.A(_03799_),
    .B(_03885_),
    .C(_02603_),
    .X(_02605_));
 sky130_fd_sc_hd__mux2_1 _15844_ (.A0(instr_auipc),
    .A1(_02605_),
    .S(_03635_),
    .X(_02606_));
 sky130_fd_sc_hd__clkbuf_1 _15845_ (.A(_02606_),
    .X(_01252_));
 sky130_fd_sc_hd__and2b_1 _15846_ (.A_N(_03804_),
    .B(_03794_),
    .X(_02607_));
 sky130_fd_sc_hd__and2_1 _15847_ (.A(_03798_),
    .B(_02607_),
    .X(_02608_));
 sky130_fd_sc_hd__a41o_1 _15848_ (.A1(_05969_),
    .A2(_03810_),
    .A3(_03864_),
    .A4(_02608_),
    .B1(_05973_),
    .X(_02609_));
 sky130_fd_sc_hd__o22a_1 _15849_ (.A1(_03402_),
    .A2(_06006_),
    .B1(_03788_),
    .B2(_02609_),
    .X(_01253_));
 sky130_fd_sc_hd__nor2b_4 _15850_ (.A(decoder_pseudo_trigger),
    .B_N(decoder_trigger),
    .Y(_02610_));
 sky130_fd_sc_hd__buf_2 _15851_ (.A(_02610_),
    .X(_02611_));
 sky130_fd_sc_hd__clkbuf_4 _15852_ (.A(\mem_rdata_q[12] ),
    .X(_02612_));
 sky130_fd_sc_hd__clkbuf_4 _15853_ (.A(\mem_rdata_q[13] ),
    .X(_02613_));
 sky130_fd_sc_hd__nor3_1 _15854_ (.A(_02612_),
    .B(_02613_),
    .C(_03940_),
    .Y(_02614_));
 sky130_fd_sc_hd__and2_1 _15855_ (.A(_03305_),
    .B(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__nor2_2 _15856_ (.A(_03239_),
    .B(_02610_),
    .Y(_02616_));
 sky130_fd_sc_hd__clkbuf_4 _15857_ (.A(_02616_),
    .X(_02617_));
 sky130_fd_sc_hd__a32o_1 _15858_ (.A1(_03309_),
    .A2(_02611_),
    .A3(_02615_),
    .B1(_02617_),
    .B2(instr_beq),
    .X(_01254_));
 sky130_fd_sc_hd__clkbuf_4 _15859_ (.A(_02616_),
    .X(_02618_));
 sky130_fd_sc_hd__or2b_1 _15860_ (.A(_02613_),
    .B_N(_02612_),
    .X(_02619_));
 sky130_fd_sc_hd__nor2_2 _15861_ (.A(_03940_),
    .B(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__and3_1 _15862_ (.A(_03309_),
    .B(_03304_),
    .C(_02610_),
    .X(_02621_));
 sky130_fd_sc_hd__clkbuf_2 _15863_ (.A(_02621_),
    .X(_02622_));
 sky130_fd_sc_hd__a22o_1 _15864_ (.A1(instr_bne),
    .A2(_02618_),
    .B1(_02620_),
    .B2(_02622_),
    .X(_01255_));
 sky130_fd_sc_hd__nor3b_2 _15865_ (.A(_02612_),
    .B(_02613_),
    .C_N(_03940_),
    .Y(_02623_));
 sky130_fd_sc_hd__a22o_1 _15866_ (.A1(instr_blt),
    .A2(_02618_),
    .B1(_02622_),
    .B2(_02623_),
    .X(_01256_));
 sky130_fd_sc_hd__and3b_1 _15867_ (.A_N(_02613_),
    .B(_03940_),
    .C(_02612_),
    .X(_02624_));
 sky130_fd_sc_hd__buf_2 _15868_ (.A(_02624_),
    .X(_02625_));
 sky130_fd_sc_hd__a22o_1 _15869_ (.A1(instr_bge),
    .A2(_02618_),
    .B1(_02622_),
    .B2(_02625_),
    .X(_01257_));
 sky130_fd_sc_hd__and3b_1 _15870_ (.A_N(_02612_),
    .B(_02613_),
    .C(_03940_),
    .X(_02626_));
 sky130_fd_sc_hd__a22o_1 _15871_ (.A1(instr_bltu),
    .A2(_02618_),
    .B1(_02622_),
    .B2(_02626_),
    .X(_01258_));
 sky130_fd_sc_hd__and3_1 _15872_ (.A(_02612_),
    .B(_02613_),
    .C(_03940_),
    .X(_02627_));
 sky130_fd_sc_hd__a22o_1 _15873_ (.A1(instr_bgeu),
    .A2(_02618_),
    .B1(_02622_),
    .B2(_02627_),
    .X(_01259_));
 sky130_fd_sc_hd__nor2_1 _15874_ (.A(_03833_),
    .B(_03770_),
    .Y(_02628_));
 sky130_fd_sc_hd__and4b_1 _15875_ (.A_N(_03768_),
    .B(_03916_),
    .C(_02603_),
    .D(_02608_),
    .X(_02629_));
 sky130_fd_sc_hd__a31o_1 _15876_ (.A1(_03790_),
    .A2(_03816_),
    .A3(_02628_),
    .B1(_02629_),
    .X(_02630_));
 sky130_fd_sc_hd__mux2_1 _15877_ (.A0(instr_jalr),
    .A1(_02630_),
    .S(_03635_),
    .X(_02631_));
 sky130_fd_sc_hd__clkbuf_1 _15878_ (.A(_02631_),
    .X(_01260_));
 sky130_fd_sc_hd__or2b_1 _15879_ (.A(decoder_pseudo_trigger),
    .B_N(decoder_trigger),
    .X(_02632_));
 sky130_fd_sc_hd__clkbuf_4 _15880_ (.A(_02632_),
    .X(_02633_));
 sky130_fd_sc_hd__clkbuf_4 _15881_ (.A(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__buf_4 _15882_ (.A(_02634_),
    .X(_02635_));
 sky130_fd_sc_hd__and2_1 _15883_ (.A(_02611_),
    .B(_02614_),
    .X(_02636_));
 sky130_fd_sc_hd__a22o_1 _15884_ (.A1(instr_lb),
    .A2(_02635_),
    .B1(_02636_),
    .B2(is_lb_lh_lw_lbu_lhu),
    .X(_01261_));
 sky130_fd_sc_hd__and2_1 _15885_ (.A(_02611_),
    .B(_02620_),
    .X(_02637_));
 sky130_fd_sc_hd__a22o_1 _15886_ (.A1(instr_lh),
    .A2(_02635_),
    .B1(_02637_),
    .B2(is_lb_lh_lw_lbu_lhu),
    .X(_01262_));
 sky130_fd_sc_hd__or3b_1 _15887_ (.A(_02612_),
    .B(\mem_rdata_q[14] ),
    .C_N(_02613_),
    .X(_02638_));
 sky130_fd_sc_hd__nor2_1 _15888_ (.A(_02634_),
    .B(_02638_),
    .Y(_02639_));
 sky130_fd_sc_hd__a22o_1 _15889_ (.A1(instr_lw),
    .A2(_02635_),
    .B1(_02639_),
    .B2(is_lb_lh_lw_lbu_lhu),
    .X(_01263_));
 sky130_fd_sc_hd__and2_1 _15890_ (.A(is_lb_lh_lw_lbu_lhu),
    .B(_02611_),
    .X(_02640_));
 sky130_fd_sc_hd__a22o_1 _15891_ (.A1(instr_lbu),
    .A2(_02635_),
    .B1(_02623_),
    .B2(_02640_),
    .X(_01264_));
 sky130_fd_sc_hd__a22o_1 _15892_ (.A1(instr_lhu),
    .A2(_02635_),
    .B1(_02625_),
    .B2(_02640_),
    .X(_01265_));
 sky130_fd_sc_hd__a22o_1 _15893_ (.A1(instr_sb),
    .A2(_02635_),
    .B1(_02636_),
    .B2(is_sb_sh_sw),
    .X(_01266_));
 sky130_fd_sc_hd__a22o_1 _15894_ (.A1(instr_sh),
    .A2(_02635_),
    .B1(_02637_),
    .B2(is_sb_sh_sw),
    .X(_01267_));
 sky130_fd_sc_hd__a32o_1 _15895_ (.A1(is_alu_reg_imm),
    .A2(_02611_),
    .A3(_02615_),
    .B1(_02616_),
    .B2(instr_addi),
    .X(_01268_));
 sky130_fd_sc_hd__nor3b_1 _15896_ (.A(_02612_),
    .B(_03940_),
    .C_N(_02613_),
    .Y(_02641_));
 sky130_fd_sc_hd__and3_1 _15897_ (.A(_03304_),
    .B(is_alu_reg_imm),
    .C(_02610_),
    .X(_02642_));
 sky130_fd_sc_hd__clkbuf_2 _15898_ (.A(_02642_),
    .X(_02643_));
 sky130_fd_sc_hd__a22o_1 _15899_ (.A1(instr_slti),
    .A2(_02618_),
    .B1(_02641_),
    .B2(_02643_),
    .X(_01269_));
 sky130_fd_sc_hd__and3b_1 _15900_ (.A_N(_03940_),
    .B(_02613_),
    .C(_02612_),
    .X(_02644_));
 sky130_fd_sc_hd__a22o_1 _15901_ (.A1(instr_sltiu),
    .A2(_02618_),
    .B1(_02643_),
    .B2(_02644_),
    .X(_01270_));
 sky130_fd_sc_hd__a22o_1 _15902_ (.A1(instr_xori),
    .A2(_02618_),
    .B1(_02623_),
    .B2(_02643_),
    .X(_01271_));
 sky130_fd_sc_hd__a22o_1 _15903_ (.A1(instr_ori),
    .A2(_02618_),
    .B1(_02626_),
    .B2(_02643_),
    .X(_01272_));
 sky130_fd_sc_hd__a22o_1 _15904_ (.A1(instr_andi),
    .A2(_02617_),
    .B1(_02627_),
    .B2(_02643_),
    .X(_01273_));
 sky130_fd_sc_hd__a22o_1 _15905_ (.A1(instr_sw),
    .A2(_02635_),
    .B1(_02639_),
    .B2(is_sb_sh_sw),
    .X(_01274_));
 sky130_fd_sc_hd__or3_1 _15906_ (.A(\mem_rdata_q[29] ),
    .B(\mem_rdata_q[30] ),
    .C(\mem_rdata_q[31] ),
    .X(_02645_));
 sky130_fd_sc_hd__or4_1 _15907_ (.A(\mem_rdata_q[28] ),
    .B(\mem_rdata_q[25] ),
    .C(\mem_rdata_q[26] ),
    .D(\mem_rdata_q[27] ),
    .X(_02646_));
 sky130_fd_sc_hd__nor2_1 _15908_ (.A(_02645_),
    .B(_02646_),
    .Y(_02647_));
 sky130_fd_sc_hd__and4_1 _15909_ (.A(is_alu_reg_imm),
    .B(_02611_),
    .C(_02620_),
    .D(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__a21o_1 _15910_ (.A1(instr_slli),
    .A2(_02635_),
    .B1(_02648_),
    .X(_01275_));
 sky130_fd_sc_hd__and2_1 _15911_ (.A(_02611_),
    .B(_02647_),
    .X(_02649_));
 sky130_fd_sc_hd__buf_4 _15912_ (.A(_02633_),
    .X(_02650_));
 sky130_fd_sc_hd__a32o_1 _15913_ (.A1(is_alu_reg_imm),
    .A2(_02625_),
    .A3(_02649_),
    .B1(_02650_),
    .B2(instr_srli),
    .X(_01276_));
 sky130_fd_sc_hd__and2_1 _15914_ (.A(_03277_),
    .B(is_alu_reg_reg),
    .X(_02651_));
 sky130_fd_sc_hd__and3_1 _15915_ (.A(_02610_),
    .B(_02647_),
    .C(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__buf_2 _15916_ (.A(_02652_),
    .X(_02653_));
 sky130_fd_sc_hd__a22o_1 _15917_ (.A1(instr_add),
    .A2(_02617_),
    .B1(_02614_),
    .B2(_02653_),
    .X(_01277_));
 sky130_fd_sc_hd__nor2_1 _15918_ (.A(\mem_rdata_q[29] ),
    .B(\mem_rdata_q[31] ),
    .Y(_02654_));
 sky130_fd_sc_hd__nor2_1 _15919_ (.A(_02633_),
    .B(_02646_),
    .Y(_02655_));
 sky130_fd_sc_hd__and3_1 _15920_ (.A(\mem_rdata_q[30] ),
    .B(_02654_),
    .C(_02655_),
    .X(_02656_));
 sky130_fd_sc_hd__a32o_1 _15921_ (.A1(is_alu_reg_reg),
    .A2(_02615_),
    .A3(_02656_),
    .B1(_02616_),
    .B2(_05517_),
    .X(_01278_));
 sky130_fd_sc_hd__a22o_1 _15922_ (.A1(instr_sll),
    .A2(_02617_),
    .B1(_02620_),
    .B2(_02653_),
    .X(_01279_));
 sky130_fd_sc_hd__a22o_1 _15923_ (.A1(instr_slt),
    .A2(_02617_),
    .B1(_02641_),
    .B2(_02653_),
    .X(_01280_));
 sky130_fd_sc_hd__a22o_1 _15924_ (.A1(instr_sltu),
    .A2(_02617_),
    .B1(_02644_),
    .B2(_02653_),
    .X(_01281_));
 sky130_fd_sc_hd__a22o_1 _15925_ (.A1(instr_xor),
    .A2(_02617_),
    .B1(_02623_),
    .B2(_02653_),
    .X(_01282_));
 sky130_fd_sc_hd__a32o_1 _15926_ (.A1(_02625_),
    .A2(_02649_),
    .A3(_02651_),
    .B1(_02616_),
    .B2(instr_srl),
    .X(_01283_));
 sky130_fd_sc_hd__a32o_1 _15927_ (.A1(_02625_),
    .A2(_02651_),
    .A3(_02656_),
    .B1(_02616_),
    .B2(instr_sra),
    .X(_01284_));
 sky130_fd_sc_hd__a22o_1 _15928_ (.A1(instr_or),
    .A2(_02617_),
    .B1(_02626_),
    .B2(_02653_),
    .X(_01285_));
 sky130_fd_sc_hd__a22o_1 _15929_ (.A1(instr_and),
    .A2(_02617_),
    .B1(_02627_),
    .B2(_02653_),
    .X(_01286_));
 sky130_fd_sc_hd__and4_1 _15930_ (.A(is_alu_reg_imm),
    .B(_02625_),
    .C(_02654_),
    .D(_02655_),
    .X(_02657_));
 sky130_fd_sc_hd__a22o_1 _15931_ (.A1(instr_srai),
    .A2(_02650_),
    .B1(_02657_),
    .B2(\mem_rdata_q[30] ),
    .X(_01287_));
 sky130_fd_sc_hd__and4bb_1 _15932_ (.A_N(\mem_rdata_q[29] ),
    .B_N(\mem_rdata_q[24] ),
    .C(\mem_rdata_q[31] ),
    .D(\mem_rdata_q[30] ),
    .X(_02658_));
 sky130_fd_sc_hd__and2_2 _15933_ (.A(_02655_),
    .B(_02658_),
    .X(_02659_));
 sky130_fd_sc_hd__or4_1 _15934_ (.A(\mem_rdata_q[2] ),
    .B(\mem_rdata_q[18] ),
    .C(\mem_rdata_q[3] ),
    .D(\mem_rdata_q[19] ),
    .X(_02660_));
 sky130_fd_sc_hd__nand2_1 _15935_ (.A(\mem_rdata_q[0] ),
    .B(\mem_rdata_q[1] ),
    .Y(_02661_));
 sky130_fd_sc_hd__or4_1 _15936_ (.A(\mem_rdata_q[16] ),
    .B(\mem_rdata_q[17] ),
    .C(_02660_),
    .D(_02661_),
    .X(_02662_));
 sky130_fd_sc_hd__and3_1 _15937_ (.A(\mem_rdata_q[5] ),
    .B(\mem_rdata_q[4] ),
    .C(\mem_rdata_q[6] ),
    .X(_02663_));
 sky130_fd_sc_hd__or4b_4 _15938_ (.A(\mem_rdata_q[15] ),
    .B(_02638_),
    .C(_02662_),
    .D_N(_02663_),
    .X(_02664_));
 sky130_fd_sc_hd__nor4_4 _15939_ (.A(\mem_rdata_q[21] ),
    .B(\mem_rdata_q[22] ),
    .C(\mem_rdata_q[23] ),
    .D(_02664_),
    .Y(_02665_));
 sky130_fd_sc_hd__a22o_1 _15940_ (.A1(instr_rdcycle),
    .A2(_02650_),
    .B1(_02659_),
    .B2(_02665_),
    .X(_01288_));
 sky130_fd_sc_hd__or3_1 _15941_ (.A(\mem_rdata_q[28] ),
    .B(\mem_rdata_q[25] ),
    .C(_02632_),
    .X(_02666_));
 sky130_fd_sc_hd__and4bb_4 _15942_ (.A_N(_02666_),
    .B_N(\mem_rdata_q[26] ),
    .C(\mem_rdata_q[27] ),
    .D(_02658_),
    .X(_02667_));
 sky130_fd_sc_hd__a22o_1 _15943_ (.A1(_04018_),
    .A2(_02650_),
    .B1(_02665_),
    .B2(_02667_),
    .X(_01289_));
 sky130_fd_sc_hd__or4b_1 _15944_ (.A(\mem_rdata_q[20] ),
    .B(\mem_rdata_q[22] ),
    .C(\mem_rdata_q[23] ),
    .D_N(\mem_rdata_q[21] ),
    .X(_02668_));
 sky130_fd_sc_hd__nor2_2 _15945_ (.A(_02664_),
    .B(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__a22o_1 _15946_ (.A1(_04012_),
    .A2(_02650_),
    .B1(_02659_),
    .B2(_02669_),
    .X(_01290_));
 sky130_fd_sc_hd__a22o_1 _15947_ (.A1(_04016_),
    .A2(_02650_),
    .B1(_02667_),
    .B2(_02669_),
    .X(_01291_));
 sky130_fd_sc_hd__or4b_1 _15948_ (.A(\mem_rdata_q[5] ),
    .B(\mem_rdata_q[4] ),
    .C(\mem_rdata_q[6] ),
    .D_N(\mem_rdata_q[3] ),
    .X(_02670_));
 sky130_fd_sc_hd__nor2_1 _15949_ (.A(_02661_),
    .B(_02670_),
    .Y(_02671_));
 sky130_fd_sc_hd__and3_1 _15950_ (.A(_03305_),
    .B(\mem_rdata_q[2] ),
    .C(_02671_),
    .X(_02672_));
 sky130_fd_sc_hd__a22o_1 _15951_ (.A1(instr_fence),
    .A2(_02617_),
    .B1(_02636_),
    .B2(_02672_),
    .X(_01292_));
 sky130_fd_sc_hd__nand2_1 _15952_ (.A(net66),
    .B(net299),
    .Y(_02673_));
 sky130_fd_sc_hd__nand2_1 _15953_ (.A(\mem_state[0] ),
    .B(\mem_state[1] ),
    .Y(_02674_));
 sky130_fd_sc_hd__or2_1 _15954_ (.A(_03196_),
    .B(net299),
    .X(_02675_));
 sky130_fd_sc_hd__buf_2 _15955_ (.A(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__inv_2 _15956_ (.A(\mem_state[1] ),
    .Y(_02677_));
 sky130_fd_sc_hd__nand2_1 _15957_ (.A(\mem_state[0] ),
    .B(_02677_),
    .Y(_02678_));
 sky130_fd_sc_hd__or4_1 _15958_ (.A(mem_do_wdata),
    .B(_03218_),
    .C(_03219_),
    .D(_03233_),
    .X(_02679_));
 sky130_fd_sc_hd__o21ai_1 _15959_ (.A1(_03757_),
    .A2(_02678_),
    .B1(_02679_),
    .Y(_02680_));
 sky130_fd_sc_hd__nand2_1 _15960_ (.A(_01821_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__or4_1 _15961_ (.A(\mem_state[0] ),
    .B(_02677_),
    .C(_03227_),
    .D(_02676_),
    .X(_02682_));
 sky130_fd_sc_hd__o211a_1 _15962_ (.A1(_02674_),
    .A2(_02676_),
    .B1(_02681_),
    .C1(_02682_),
    .X(_02683_));
 sky130_fd_sc_hd__o21ai_1 _15963_ (.A1(net65),
    .A2(_02673_),
    .B1(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__inv_2 _15964_ (.A(net224),
    .Y(_02685_));
 sky130_fd_sc_hd__or2_1 _15965_ (.A(_02685_),
    .B(_02678_),
    .X(_02686_));
 sky130_fd_sc_hd__a22o_1 _15966_ (.A1(_03286_),
    .A2(_03198_),
    .B1(_03233_),
    .B2(_02674_),
    .X(_02687_));
 sky130_fd_sc_hd__a21oi_1 _15967_ (.A1(_02686_),
    .A2(_02687_),
    .B1(_02684_),
    .Y(_02688_));
 sky130_fd_sc_hd__a22o_1 _15968_ (.A1(net262),
    .A2(_02684_),
    .B1(_02688_),
    .B2(_01821_),
    .X(_01293_));
 sky130_fd_sc_hd__o21a_1 _15969_ (.A1(_04168_),
    .A2(_03636_),
    .B1(_06003_),
    .X(_01294_));
 sky130_fd_sc_hd__nor2_1 _15970_ (.A(\mem_rdata_q[2] ),
    .B(\mem_rdata_q[28] ),
    .Y(_02689_));
 sky130_fd_sc_hd__and4_1 _15971_ (.A(\mem_rdata_q[25] ),
    .B(_02610_),
    .C(_02671_),
    .D(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__nor2_1 _15972_ (.A(\mem_rdata_q[27] ),
    .B(_02645_),
    .Y(_02691_));
 sky130_fd_sc_hd__a32o_2 _15973_ (.A1(\mem_rdata_q[26] ),
    .A2(_02690_),
    .A3(_02691_),
    .B1(_02650_),
    .B2(_04022_),
    .X(_01295_));
 sky130_fd_sc_hd__or4b_1 _15974_ (.A(_03965_),
    .B(_05999_),
    .C(_06000_),
    .D_N(_03977_),
    .X(_02692_));
 sky130_fd_sc_hd__nor2_1 _15975_ (.A(_05998_),
    .B(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__mux2_1 _15976_ (.A0(instr_waitirq),
    .A1(_02693_),
    .S(_03635_),
    .X(_02694_));
 sky130_fd_sc_hd__clkbuf_1 _15977_ (.A(_02694_),
    .X(_01296_));
 sky130_fd_sc_hd__and4bb_2 _15978_ (.A_N(_02645_),
    .B_N(\mem_rdata_q[26] ),
    .C(\mem_rdata_q[27] ),
    .D(_02690_),
    .X(_02695_));
 sky130_fd_sc_hd__a21o_1 _15979_ (.A1(_04024_),
    .A2(_02635_),
    .B1(_02695_),
    .X(_01297_));
 sky130_fd_sc_hd__a31o_1 _15980_ (.A1(_03891_),
    .A2(_03767_),
    .A3(_02600_),
    .B1(_03862_),
    .X(_02696_));
 sky130_fd_sc_hd__nand2_1 _15981_ (.A(_03783_),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__o21ai_1 _15982_ (.A1(_03743_),
    .A2(_03916_),
    .B1(_03862_),
    .Y(_02698_));
 sky130_fd_sc_hd__nor2_1 _15983_ (.A(_03844_),
    .B(_05963_),
    .Y(_02699_));
 sky130_fd_sc_hd__a21bo_1 _15984_ (.A1(_03856_),
    .A2(_02698_),
    .B1_N(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__and3_1 _15985_ (.A(_03228_),
    .B(_02697_),
    .C(_02700_),
    .X(_02701_));
 sky130_fd_sc_hd__nand2_1 _15986_ (.A(_05990_),
    .B(_02701_),
    .Y(_02702_));
 sky130_fd_sc_hd__a22o_1 _15987_ (.A1(_03767_),
    .A2(_03788_),
    .B1(_03864_),
    .B2(_03880_),
    .X(_02703_));
 sky130_fd_sc_hd__a41o_1 _15988_ (.A1(_03816_),
    .A2(_03737_),
    .A3(_02628_),
    .A4(_02699_),
    .B1(_02703_),
    .X(_02704_));
 sky130_fd_sc_hd__a22o_1 _15989_ (.A1(\decoded_rd[0] ),
    .A2(_05973_),
    .B1(_06016_),
    .B2(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__a31o_1 _15990_ (.A1(_03636_),
    .A2(_03822_),
    .A3(_02702_),
    .B1(_02705_),
    .X(_01298_));
 sky130_fd_sc_hd__nor2_1 _15991_ (.A(_05970_),
    .B(_02701_),
    .Y(_02706_));
 sky130_fd_sc_hd__a21o_1 _15992_ (.A1(_06016_),
    .A2(_05991_),
    .B1(_02706_),
    .X(_02707_));
 sky130_fd_sc_hd__a22o_1 _15993_ (.A1(\decoded_rd[1] ),
    .A2(_05987_),
    .B1(_03880_),
    .B2(_05977_),
    .X(_02708_));
 sky130_fd_sc_hd__a21o_1 _15994_ (.A1(_03867_),
    .A2(_02707_),
    .B1(_02708_),
    .X(_01299_));
 sky130_fd_sc_hd__a221o_1 _15995_ (.A1(_03885_),
    .A2(_03880_),
    .B1(_02702_),
    .B2(_03826_),
    .C1(_05973_),
    .X(_02709_));
 sky130_fd_sc_hd__o21a_1 _15996_ (.A1(\decoded_rd[2] ),
    .A2(_03636_),
    .B1(_02709_),
    .X(_01300_));
 sky130_fd_sc_hd__a21oi_1 _15997_ (.A1(_03893_),
    .A2(_05990_),
    .B1(_05976_),
    .Y(_02710_));
 sky130_fd_sc_hd__a221o_1 _15998_ (.A1(\decoded_rd[3] ),
    .A2(_05987_),
    .B1(_03892_),
    .B2(_02706_),
    .C1(_02710_),
    .X(_01301_));
 sky130_fd_sc_hd__a22o_1 _15999_ (.A1(\decoded_rd[4] ),
    .A2(_05974_),
    .B1(_03763_),
    .B2(_02706_),
    .X(_01302_));
 sky130_fd_sc_hd__o21a_1 _16000_ (.A1(\cpuregs.raddr1[0] ),
    .A2(_03636_),
    .B1(_06005_),
    .X(_01303_));
 sky130_fd_sc_hd__o211a_1 _16001_ (.A1(\cpuregs.raddr1[1] ),
    .A2(_06006_),
    .B1(_06014_),
    .C1(_06015_),
    .X(_01304_));
 sky130_fd_sc_hd__a31o_1 _16002_ (.A1(_03826_),
    .A2(_06016_),
    .A3(_05996_),
    .B1(_06018_),
    .X(_01305_));
 sky130_fd_sc_hd__o22a_1 _16003_ (.A1(\cpuregs.raddr1[3] ),
    .A2(_06006_),
    .B1(_06020_),
    .B2(_06022_),
    .X(_01306_));
 sky130_fd_sc_hd__a41o_1 _16004_ (.A1(_03635_),
    .A2(_03763_),
    .A3(_05995_),
    .A4(_06023_),
    .B1(_06025_),
    .X(_01307_));
 sky130_fd_sc_hd__o22a_1 _16005_ (.A1(\cpuregs.raddr2[0] ),
    .A2(_06006_),
    .B1(_05968_),
    .B2(_05972_),
    .X(_01308_));
 sky130_fd_sc_hd__a22o_1 _16006_ (.A1(\cpuregs.raddr2[1] ),
    .A2(_05974_),
    .B1(_05975_),
    .B2(_05978_),
    .X(_01309_));
 sky130_fd_sc_hd__a22o_1 _16007_ (.A1(\cpuregs.raddr2[2] ),
    .A2(_05974_),
    .B1(_05980_),
    .B2(_05982_),
    .X(_01310_));
 sky130_fd_sc_hd__a211o_1 _16008_ (.A1(\cpuregs.raddr2[3] ),
    .A2(_05983_),
    .B1(_05984_),
    .C1(_05985_),
    .X(_01311_));
 sky130_fd_sc_hd__o22a_1 _16009_ (.A1(\cpuregs.raddr2[4] ),
    .A2(_06006_),
    .B1(_05986_),
    .B2(_05988_),
    .X(_01312_));
 sky130_fd_sc_hd__clkbuf_4 _16010_ (.A(_02611_),
    .X(_02711_));
 sky130_fd_sc_hd__or3_2 _16011_ (.A(instr_jalr),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(is_alu_reg_imm),
    .X(_02712_));
 sky130_fd_sc_hd__a221o_1 _16012_ (.A1(is_sb_sh_sw),
    .A2(\mem_rdata_q[7] ),
    .B1(_02712_),
    .B2(\mem_rdata_q[20] ),
    .C1(_02634_),
    .X(_02713_));
 sky130_fd_sc_hd__o21a_1 _16013_ (.A1(\decoded_imm[0] ),
    .A2(_02711_),
    .B1(_02713_),
    .X(_01313_));
 sky130_fd_sc_hd__and2_1 _16014_ (.A(\mem_rdata_q[21] ),
    .B(_02712_),
    .X(_02714_));
 sky130_fd_sc_hd__buf_2 _16015_ (.A(instr_jal),
    .X(_02715_));
 sky130_fd_sc_hd__or2_1 _16016_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(is_sb_sh_sw),
    .X(_02716_));
 sky130_fd_sc_hd__a221o_1 _16017_ (.A1(_02715_),
    .A2(\decoded_imm_j[1] ),
    .B1(\mem_rdata_q[8] ),
    .B2(_02716_),
    .C1(_02633_),
    .X(_02717_));
 sky130_fd_sc_hd__o22a_1 _16018_ (.A1(\decoded_imm[1] ),
    .A2(_02711_),
    .B1(_02714_),
    .B2(_02717_),
    .X(_01314_));
 sky130_fd_sc_hd__and2_1 _16019_ (.A(\mem_rdata_q[22] ),
    .B(_02712_),
    .X(_02718_));
 sky130_fd_sc_hd__a221o_1 _16020_ (.A1(_02715_),
    .A2(\decoded_imm_j[2] ),
    .B1(_02716_),
    .B2(\mem_rdata_q[9] ),
    .C1(_02633_),
    .X(_02719_));
 sky130_fd_sc_hd__o22a_1 _16021_ (.A1(\decoded_imm[2] ),
    .A2(_02711_),
    .B1(_02718_),
    .B2(_02719_),
    .X(_01315_));
 sky130_fd_sc_hd__clkbuf_4 _16022_ (.A(_02611_),
    .X(_02720_));
 sky130_fd_sc_hd__and2_1 _16023_ (.A(\mem_rdata_q[23] ),
    .B(_02712_),
    .X(_02721_));
 sky130_fd_sc_hd__a221o_1 _16024_ (.A1(_02715_),
    .A2(\decoded_imm_j[3] ),
    .B1(_02716_),
    .B2(\mem_rdata_q[10] ),
    .C1(_02633_),
    .X(_02722_));
 sky130_fd_sc_hd__o22a_1 _16025_ (.A1(\decoded_imm[3] ),
    .A2(_02720_),
    .B1(_02721_),
    .B2(_02722_),
    .X(_01316_));
 sky130_fd_sc_hd__and2_1 _16026_ (.A(\mem_rdata_q[24] ),
    .B(_02712_),
    .X(_02723_));
 sky130_fd_sc_hd__a221o_1 _16027_ (.A1(_02715_),
    .A2(\decoded_imm_j[4] ),
    .B1(_02716_),
    .B2(\mem_rdata_q[11] ),
    .C1(_02633_),
    .X(_02724_));
 sky130_fd_sc_hd__o22a_1 _16028_ (.A1(\decoded_imm[4] ),
    .A2(_02720_),
    .B1(_02723_),
    .B2(_02724_),
    .X(_01317_));
 sky130_fd_sc_hd__or2_1 _16029_ (.A(_02712_),
    .B(_02716_),
    .X(_02725_));
 sky130_fd_sc_hd__buf_2 _16030_ (.A(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__and3_1 _16031_ (.A(instr_jal),
    .B(\decoded_imm_j[5] ),
    .C(_02610_),
    .X(_02727_));
 sky130_fd_sc_hd__a21o_1 _16032_ (.A1(\decoded_imm[5] ),
    .A2(_02634_),
    .B1(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__a31o_1 _16033_ (.A1(\mem_rdata_q[25] ),
    .A2(_02711_),
    .A3(_02726_),
    .B1(_02728_),
    .X(_01318_));
 sky130_fd_sc_hd__a221o_1 _16034_ (.A1(_02715_),
    .A2(\decoded_imm_j[6] ),
    .B1(_02726_),
    .B2(\mem_rdata_q[26] ),
    .C1(_02634_),
    .X(_02729_));
 sky130_fd_sc_hd__o21a_1 _16035_ (.A1(\decoded_imm[6] ),
    .A2(_02711_),
    .B1(_02729_),
    .X(_01319_));
 sky130_fd_sc_hd__a221o_1 _16036_ (.A1(_02715_),
    .A2(\decoded_imm_j[7] ),
    .B1(_02726_),
    .B2(\mem_rdata_q[27] ),
    .C1(_02634_),
    .X(_02730_));
 sky130_fd_sc_hd__o21a_1 _16037_ (.A1(\decoded_imm[7] ),
    .A2(_02711_),
    .B1(_02730_),
    .X(_01320_));
 sky130_fd_sc_hd__a221o_1 _16038_ (.A1(_02715_),
    .A2(\decoded_imm_j[8] ),
    .B1(_02726_),
    .B2(\mem_rdata_q[28] ),
    .C1(_02634_),
    .X(_02731_));
 sky130_fd_sc_hd__o21a_1 _16039_ (.A1(\decoded_imm[8] ),
    .A2(_02711_),
    .B1(_02731_),
    .X(_01321_));
 sky130_fd_sc_hd__a221o_1 _16040_ (.A1(_02715_),
    .A2(\decoded_imm_j[9] ),
    .B1(_02726_),
    .B2(\mem_rdata_q[29] ),
    .C1(_02634_),
    .X(_02732_));
 sky130_fd_sc_hd__o21a_1 _16041_ (.A1(\decoded_imm[9] ),
    .A2(_02711_),
    .B1(_02732_),
    .X(_01322_));
 sky130_fd_sc_hd__a221o_1 _16042_ (.A1(_02715_),
    .A2(\decoded_imm_j[10] ),
    .B1(_02726_),
    .B2(\mem_rdata_q[30] ),
    .C1(_02634_),
    .X(_02733_));
 sky130_fd_sc_hd__o21a_1 _16043_ (.A1(\decoded_imm[10] ),
    .A2(_02711_),
    .B1(_02733_),
    .X(_01323_));
 sky130_fd_sc_hd__o21a_1 _16044_ (.A1(is_sb_sh_sw),
    .A2(_02712_),
    .B1(\mem_rdata_q[31] ),
    .X(_02734_));
 sky130_fd_sc_hd__a221o_1 _16045_ (.A1(_02715_),
    .A2(\decoded_imm_j[11] ),
    .B1(\mem_rdata_q[7] ),
    .B2(_03309_),
    .C1(_02633_),
    .X(_02735_));
 sky130_fd_sc_hd__o22a_1 _16046_ (.A1(\decoded_imm[11] ),
    .A2(_02720_),
    .B1(_02734_),
    .B2(_02735_),
    .X(_01324_));
 sky130_fd_sc_hd__a21o_2 _16047_ (.A1(\mem_rdata_q[31] ),
    .A2(_02726_),
    .B1(_02633_),
    .X(_02736_));
 sky130_fd_sc_hd__a22o_1 _16048_ (.A1(_03402_),
    .A2(\decoded_imm_j[12] ),
    .B1(_03403_),
    .B2(_02612_),
    .X(_02737_));
 sky130_fd_sc_hd__o22a_1 _16049_ (.A1(\decoded_imm[12] ),
    .A2(_02720_),
    .B1(_02736_),
    .B2(_02737_),
    .X(_01325_));
 sky130_fd_sc_hd__a22o_1 _16050_ (.A1(_03402_),
    .A2(\decoded_imm_j[13] ),
    .B1(_03403_),
    .B2(_02613_),
    .X(_02738_));
 sky130_fd_sc_hd__o22a_1 _16051_ (.A1(\decoded_imm[13] ),
    .A2(_02720_),
    .B1(_02736_),
    .B2(_02738_),
    .X(_01326_));
 sky130_fd_sc_hd__a22o_1 _16052_ (.A1(_03402_),
    .A2(\decoded_imm_j[14] ),
    .B1(_03403_),
    .B2(_03940_),
    .X(_02739_));
 sky130_fd_sc_hd__o22a_1 _16053_ (.A1(\decoded_imm[14] ),
    .A2(_02720_),
    .B1(_02736_),
    .B2(_02739_),
    .X(_01327_));
 sky130_fd_sc_hd__a22o_1 _16054_ (.A1(_03402_),
    .A2(\decoded_imm_j[15] ),
    .B1(_03403_),
    .B2(\mem_rdata_q[15] ),
    .X(_02740_));
 sky130_fd_sc_hd__o22a_1 _16055_ (.A1(\decoded_imm[15] ),
    .A2(_02720_),
    .B1(_02736_),
    .B2(_02740_),
    .X(_01328_));
 sky130_fd_sc_hd__a22o_1 _16056_ (.A1(_03402_),
    .A2(\decoded_imm_j[16] ),
    .B1(_03403_),
    .B2(\mem_rdata_q[16] ),
    .X(_02741_));
 sky130_fd_sc_hd__o22a_1 _16057_ (.A1(\decoded_imm[16] ),
    .A2(_02720_),
    .B1(_02736_),
    .B2(_02741_),
    .X(_01329_));
 sky130_fd_sc_hd__a22o_1 _16058_ (.A1(_03402_),
    .A2(\decoded_imm_j[17] ),
    .B1(_03403_),
    .B2(\mem_rdata_q[17] ),
    .X(_02742_));
 sky130_fd_sc_hd__o22a_1 _16059_ (.A1(\decoded_imm[17] ),
    .A2(_02720_),
    .B1(_02736_),
    .B2(_02742_),
    .X(_01330_));
 sky130_fd_sc_hd__a22o_1 _16060_ (.A1(_03402_),
    .A2(\decoded_imm_j[18] ),
    .B1(_03403_),
    .B2(\mem_rdata_q[18] ),
    .X(_02743_));
 sky130_fd_sc_hd__o22a_1 _16061_ (.A1(\decoded_imm[18] ),
    .A2(_02720_),
    .B1(_02736_),
    .B2(_02743_),
    .X(_01331_));
 sky130_fd_sc_hd__a22o_1 _16062_ (.A1(_03402_),
    .A2(\decoded_imm_j[19] ),
    .B1(_03403_),
    .B2(\mem_rdata_q[19] ),
    .X(_02744_));
 sky130_fd_sc_hd__o22a_1 _16063_ (.A1(\decoded_imm[19] ),
    .A2(_02611_),
    .B1(_02736_),
    .B2(_02744_),
    .X(_01332_));
 sky130_fd_sc_hd__and2_1 _16064_ (.A(_03403_),
    .B(_02610_),
    .X(_02745_));
 sky130_fd_sc_hd__buf_2 _16065_ (.A(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__a22o_1 _16066_ (.A1(instr_jal),
    .A2(_08232_),
    .B1(_02726_),
    .B2(\mem_rdata_q[31] ),
    .X(_02747_));
 sky130_fd_sc_hd__and2_1 _16067_ (.A(_02610_),
    .B(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__buf_2 _16068_ (.A(_02748_),
    .X(_02749_));
 sky130_fd_sc_hd__a221o_1 _16069_ (.A1(\decoded_imm[20] ),
    .A2(_02650_),
    .B1(_02746_),
    .B2(\mem_rdata_q[20] ),
    .C1(_02749_),
    .X(_01333_));
 sky130_fd_sc_hd__a221o_1 _16070_ (.A1(\decoded_imm[21] ),
    .A2(_02650_),
    .B1(_02746_),
    .B2(\mem_rdata_q[21] ),
    .C1(_02749_),
    .X(_01334_));
 sky130_fd_sc_hd__buf_2 _16071_ (.A(_02633_),
    .X(_02750_));
 sky130_fd_sc_hd__a221o_1 _16072_ (.A1(\decoded_imm[22] ),
    .A2(_02750_),
    .B1(_02746_),
    .B2(\mem_rdata_q[22] ),
    .C1(_02749_),
    .X(_01335_));
 sky130_fd_sc_hd__a221o_1 _16073_ (.A1(\decoded_imm[23] ),
    .A2(_02750_),
    .B1(_02746_),
    .B2(\mem_rdata_q[23] ),
    .C1(_02749_),
    .X(_01336_));
 sky130_fd_sc_hd__a221o_1 _16074_ (.A1(\decoded_imm[24] ),
    .A2(_02750_),
    .B1(_02746_),
    .B2(\mem_rdata_q[24] ),
    .C1(_02749_),
    .X(_01337_));
 sky130_fd_sc_hd__a221o_1 _16075_ (.A1(\decoded_imm[25] ),
    .A2(_02750_),
    .B1(_02746_),
    .B2(\mem_rdata_q[25] ),
    .C1(_02749_),
    .X(_01338_));
 sky130_fd_sc_hd__a221o_1 _16076_ (.A1(\decoded_imm[26] ),
    .A2(_02750_),
    .B1(_02746_),
    .B2(\mem_rdata_q[26] ),
    .C1(_02749_),
    .X(_01339_));
 sky130_fd_sc_hd__a221o_1 _16077_ (.A1(\decoded_imm[27] ),
    .A2(_02750_),
    .B1(_02746_),
    .B2(\mem_rdata_q[27] ),
    .C1(_02749_),
    .X(_01340_));
 sky130_fd_sc_hd__a221o_1 _16078_ (.A1(\decoded_imm[28] ),
    .A2(_02750_),
    .B1(_02746_),
    .B2(\mem_rdata_q[28] ),
    .C1(_02749_),
    .X(_01341_));
 sky130_fd_sc_hd__a221o_1 _16079_ (.A1(\decoded_imm[29] ),
    .A2(_02750_),
    .B1(_02746_),
    .B2(\mem_rdata_q[29] ),
    .C1(_02749_),
    .X(_01342_));
 sky130_fd_sc_hd__a221o_1 _16080_ (.A1(\decoded_imm[30] ),
    .A2(_02750_),
    .B1(_02745_),
    .B2(\mem_rdata_q[30] ),
    .C1(_02748_),
    .X(_01343_));
 sky130_fd_sc_hd__a221o_1 _16081_ (.A1(\decoded_imm[31] ),
    .A2(_02750_),
    .B1(_02745_),
    .B2(\mem_rdata_q[31] ),
    .C1(_02748_),
    .X(_01344_));
 sky130_fd_sc_hd__a21o_1 _16082_ (.A1(compressed_instr),
    .A2(_05974_),
    .B1(_06016_),
    .X(_01345_));
 sky130_fd_sc_hd__nand2_1 _16083_ (.A(_03213_),
    .B(_03833_),
    .Y(_02751_));
 sky130_fd_sc_hd__a32o_1 _16084_ (.A1(_03767_),
    .A2(_03935_),
    .A3(_02751_),
    .B1(_03816_),
    .B2(_03215_),
    .X(_02752_));
 sky130_fd_sc_hd__mux2_1 _16085_ (.A0(is_lb_lh_lw_lbu_lhu),
    .A1(_02752_),
    .S(_03635_),
    .X(_02753_));
 sky130_fd_sc_hd__clkbuf_1 _16086_ (.A(_02753_),
    .X(_01346_));
 sky130_fd_sc_hd__a211o_1 _16087_ (.A1(is_slli_srli_srai),
    .A2(_02650_),
    .B1(_02648_),
    .C1(_02657_),
    .X(_01347_));
 sky130_fd_sc_hd__a211o_1 _16088_ (.A1(is_alu_reg_imm),
    .A2(_02619_),
    .B1(_02634_),
    .C1(instr_jalr),
    .X(_02754_));
 sky130_fd_sc_hd__o21a_1 _16089_ (.A1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .A2(_02711_),
    .B1(_02754_),
    .X(_01348_));
 sky130_fd_sc_hd__nor2_1 _16090_ (.A(_03228_),
    .B(_03815_),
    .Y(_02755_));
 sky130_fd_sc_hd__and4b_1 _16091_ (.A_N(_03878_),
    .B(_02607_),
    .C(_02755_),
    .D(_03783_),
    .X(_02756_));
 sky130_fd_sc_hd__a211o_1 _16092_ (.A1(_03781_),
    .A2(_03935_),
    .B1(_02756_),
    .C1(_05987_),
    .X(_02757_));
 sky130_fd_sc_hd__o21a_1 _16093_ (.A1(is_sb_sh_sw),
    .A2(_03636_),
    .B1(_02757_),
    .X(_01349_));
 sky130_fd_sc_hd__a211o_1 _16094_ (.A1(_02608_),
    .A2(_02755_),
    .B1(_05973_),
    .C1(_03845_),
    .X(_02758_));
 sky130_fd_sc_hd__o211a_1 _16095_ (.A1(_03309_),
    .A2(_06006_),
    .B1(_02758_),
    .C1(_06026_),
    .X(_01350_));
 sky130_fd_sc_hd__o21a_1 _16096_ (.A1(_03762_),
    .A2(_03736_),
    .B1(_03776_),
    .X(_02759_));
 sky130_fd_sc_hd__o221a_1 _16097_ (.A1(_03747_),
    .A2(_03781_),
    .B1(_03768_),
    .B2(_02759_),
    .C1(_06009_),
    .X(_02760_));
 sky130_fd_sc_hd__a311o_1 _16098_ (.A1(_03799_),
    .A2(_03833_),
    .A3(_03916_),
    .B1(_03893_),
    .C1(_03891_),
    .X(_02761_));
 sky130_fd_sc_hd__o211a_1 _16099_ (.A1(_03854_),
    .A2(_02760_),
    .B1(_02761_),
    .C1(_05993_),
    .X(_02762_));
 sky130_fd_sc_hd__a2bb2o_1 _16100_ (.A1_N(_02762_),
    .A2_N(_05976_),
    .B1(_05973_),
    .B2(is_alu_reg_imm),
    .X(_02763_));
 sky130_fd_sc_hd__a41o_1 _16101_ (.A1(_03635_),
    .A2(_03799_),
    .A3(_03885_),
    .A4(_02755_),
    .B1(_02763_),
    .X(_01351_));
 sky130_fd_sc_hd__o21ba_1 _16102_ (.A1(_03783_),
    .A2(_03856_),
    .B1_N(_05961_),
    .X(_02764_));
 sky130_fd_sc_hd__a21oi_1 _16103_ (.A1(_02602_),
    .A2(_02755_),
    .B1(_06023_),
    .Y(_02765_));
 sky130_fd_sc_hd__a21oi_1 _16104_ (.A1(_06023_),
    .A2(_02764_),
    .B1(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__mux2_1 _16105_ (.A0(is_alu_reg_reg),
    .A1(_02766_),
    .S(_03635_),
    .X(_02767_));
 sky130_fd_sc_hd__clkbuf_1 _16106_ (.A(_02767_),
    .X(_01352_));
 sky130_fd_sc_hd__o21a_1 _16107_ (.A1(_03309_),
    .A2(_03255_),
    .B1(_02618_),
    .X(_01353_));
 sky130_fd_sc_hd__and3_1 _16108_ (.A(_03286_),
    .B(_03220_),
    .C(_01821_),
    .X(_02768_));
 sky130_fd_sc_hd__and3_1 _16109_ (.A(mem_do_wdata),
    .B(_03220_),
    .C(_01821_),
    .X(_02769_));
 sky130_fd_sc_hd__buf_2 _16110_ (.A(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__buf_4 _16111_ (.A(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__o21ba_1 _16112_ (.A1(_03221_),
    .A2(_02676_),
    .B1_N(_02771_),
    .X(_02772_));
 sky130_fd_sc_hd__a22o_1 _16113_ (.A1(_05829_),
    .A2(_02768_),
    .B1(_02772_),
    .B2(net193),
    .X(_01354_));
 sky130_fd_sc_hd__o31a_1 _16114_ (.A1(_03199_),
    .A2(_02674_),
    .A3(_02676_),
    .B1(_02673_),
    .X(_02773_));
 sky130_fd_sc_hd__and3_1 _16115_ (.A(_02681_),
    .B(_02682_),
    .C(_02773_),
    .X(_02774_));
 sky130_fd_sc_hd__and2_1 _16116_ (.A(_02686_),
    .B(_02774_),
    .X(_02775_));
 sky130_fd_sc_hd__o41a_1 _16117_ (.A1(_03218_),
    .A2(_03199_),
    .A3(_02676_),
    .A4(_02678_),
    .B1(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__inv_2 _16118_ (.A(_02776_),
    .Y(_02777_));
 sky130_fd_sc_hd__o22a_1 _16119_ (.A1(\mem_state[0] ),
    .A2(_02774_),
    .B1(_02777_),
    .B2(_02768_),
    .X(_01355_));
 sky130_fd_sc_hd__o22a_1 _16120_ (.A1(\mem_state[1] ),
    .A2(_02775_),
    .B1(_02777_),
    .B2(_02771_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _16121_ (.A0(net263),
    .A1(_05324_),
    .S(_02771_),
    .X(_02778_));
 sky130_fd_sc_hd__clkbuf_1 _16122_ (.A(_02778_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _16123_ (.A0(net274),
    .A1(_05286_),
    .S(_02771_),
    .X(_02779_));
 sky130_fd_sc_hd__clkbuf_1 _16124_ (.A(_02779_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _16125_ (.A0(net285),
    .A1(_05413_),
    .S(_02771_),
    .X(_02780_));
 sky130_fd_sc_hd__clkbuf_1 _16126_ (.A(_02780_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _16127_ (.A0(net288),
    .A1(_05414_),
    .S(_02771_),
    .X(_02781_));
 sky130_fd_sc_hd__clkbuf_1 _16128_ (.A(_02781_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _16129_ (.A0(net289),
    .A1(_05255_),
    .S(_02771_),
    .X(_02782_));
 sky130_fd_sc_hd__clkbuf_1 _16130_ (.A(_02782_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _16131_ (.A0(net290),
    .A1(net126),
    .S(_02771_),
    .X(_02783_));
 sky130_fd_sc_hd__clkbuf_1 _16132_ (.A(_02783_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _16133_ (.A0(net291),
    .A1(net127),
    .S(_02771_),
    .X(_02784_));
 sky130_fd_sc_hd__clkbuf_1 _16134_ (.A(_02784_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _16135_ (.A0(net292),
    .A1(net128),
    .S(_02771_),
    .X(_02785_));
 sky130_fd_sc_hd__clkbuf_1 _16136_ (.A(_02785_),
    .X(_01364_));
 sky130_fd_sc_hd__clkbuf_4 _16137_ (.A(_02770_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_1 _16138_ (.A0(net293),
    .A1(net255),
    .S(_02786_),
    .X(_02787_));
 sky130_fd_sc_hd__clkbuf_1 _16139_ (.A(_02787_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _16140_ (.A0(net294),
    .A1(net256),
    .S(_02786_),
    .X(_02788_));
 sky130_fd_sc_hd__clkbuf_1 _16141_ (.A(_02788_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _16142_ (.A0(net264),
    .A1(net226),
    .S(_02786_),
    .X(_02789_));
 sky130_fd_sc_hd__clkbuf_1 _16143_ (.A(_02789_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _16144_ (.A0(net265),
    .A1(net227),
    .S(_02786_),
    .X(_02790_));
 sky130_fd_sc_hd__clkbuf_1 _16145_ (.A(_02790_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _16146_ (.A0(net266),
    .A1(net228),
    .S(_02786_),
    .X(_02791_));
 sky130_fd_sc_hd__clkbuf_1 _16147_ (.A(_02791_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _16148_ (.A0(net267),
    .A1(net229),
    .S(_02786_),
    .X(_02792_));
 sky130_fd_sc_hd__clkbuf_1 _16149_ (.A(_02792_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _16150_ (.A0(net268),
    .A1(net230),
    .S(_02786_),
    .X(_02793_));
 sky130_fd_sc_hd__clkbuf_1 _16151_ (.A(_02793_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _16152_ (.A0(net269),
    .A1(net231),
    .S(_02786_),
    .X(_02794_));
 sky130_fd_sc_hd__clkbuf_1 _16153_ (.A(_02794_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _16154_ (.A0(net270),
    .A1(net232),
    .S(_02786_),
    .X(_02795_));
 sky130_fd_sc_hd__clkbuf_1 _16155_ (.A(_02795_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _16156_ (.A0(net271),
    .A1(net233),
    .S(_02786_),
    .X(_02796_));
 sky130_fd_sc_hd__clkbuf_1 _16157_ (.A(_02796_),
    .X(_01374_));
 sky130_fd_sc_hd__clkbuf_4 _16158_ (.A(_02770_),
    .X(_02797_));
 sky130_fd_sc_hd__mux2_1 _16159_ (.A0(net272),
    .A1(net234),
    .S(_02797_),
    .X(_02798_));
 sky130_fd_sc_hd__clkbuf_1 _16160_ (.A(_02798_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _16161_ (.A0(net273),
    .A1(net235),
    .S(_02797_),
    .X(_02799_));
 sky130_fd_sc_hd__clkbuf_1 _16162_ (.A(_02799_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _16163_ (.A0(net275),
    .A1(net237),
    .S(_02797_),
    .X(_02800_));
 sky130_fd_sc_hd__clkbuf_1 _16164_ (.A(_02800_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _16165_ (.A0(net276),
    .A1(net238),
    .S(_02797_),
    .X(_02801_));
 sky130_fd_sc_hd__clkbuf_1 _16166_ (.A(_02801_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _16167_ (.A0(net277),
    .A1(net239),
    .S(_02797_),
    .X(_02802_));
 sky130_fd_sc_hd__clkbuf_1 _16168_ (.A(_02802_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _16169_ (.A0(net278),
    .A1(net240),
    .S(_02797_),
    .X(_02803_));
 sky130_fd_sc_hd__clkbuf_1 _16170_ (.A(_02803_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _16171_ (.A0(net279),
    .A1(net241),
    .S(_02797_),
    .X(_02804_));
 sky130_fd_sc_hd__clkbuf_1 _16172_ (.A(_02804_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _16173_ (.A0(net280),
    .A1(net242),
    .S(_02797_),
    .X(_02805_));
 sky130_fd_sc_hd__clkbuf_1 _16174_ (.A(_02805_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _16175_ (.A0(net281),
    .A1(net243),
    .S(_02797_),
    .X(_02806_));
 sky130_fd_sc_hd__clkbuf_1 _16176_ (.A(_02806_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _16177_ (.A0(net282),
    .A1(net244),
    .S(_02797_),
    .X(_02807_));
 sky130_fd_sc_hd__clkbuf_1 _16178_ (.A(_02807_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _16179_ (.A0(net283),
    .A1(net245),
    .S(_02770_),
    .X(_02808_));
 sky130_fd_sc_hd__clkbuf_1 _16180_ (.A(_02808_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _16181_ (.A0(net284),
    .A1(net246),
    .S(_02770_),
    .X(_02809_));
 sky130_fd_sc_hd__clkbuf_1 _16182_ (.A(_02809_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _16183_ (.A0(net286),
    .A1(net248),
    .S(_02770_),
    .X(_02810_));
 sky130_fd_sc_hd__clkbuf_1 _16184_ (.A(_02810_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _16185_ (.A0(net287),
    .A1(net249),
    .S(_02770_),
    .X(_02811_));
 sky130_fd_sc_hd__clkbuf_1 _16186_ (.A(_02811_),
    .X(_01388_));
 sky130_fd_sc_hd__or2_1 _16187_ (.A(net295),
    .B(_01822_),
    .X(_02812_));
 sky130_fd_sc_hd__a21bo_1 _16188_ (.A1(net257),
    .A2(net258),
    .B1_N(_01822_),
    .X(_02813_));
 sky130_fd_sc_hd__and2_1 _16189_ (.A(_03221_),
    .B(_01821_),
    .X(_02814_));
 sky130_fd_sc_hd__a32o_1 _16190_ (.A1(_02812_),
    .A2(_02813_),
    .A3(_02814_),
    .B1(_02676_),
    .B2(net295),
    .X(_01389_));
 sky130_fd_sc_hd__or2_1 _16191_ (.A(net296),
    .B(_01822_),
    .X(_02815_));
 sky130_fd_sc_hd__a21bo_1 _16192_ (.A1(net257),
    .A2(net259),
    .B1_N(_01822_),
    .X(_02816_));
 sky130_fd_sc_hd__a32o_1 _16193_ (.A1(_02814_),
    .A2(_02815_),
    .A3(_02816_),
    .B1(_02676_),
    .B2(net296),
    .X(_01390_));
 sky130_fd_sc_hd__or2_1 _16194_ (.A(net297),
    .B(_01822_),
    .X(_02817_));
 sky130_fd_sc_hd__a21bo_1 _16195_ (.A1(net257),
    .A2(net260),
    .B1_N(_01822_),
    .X(_02818_));
 sky130_fd_sc_hd__a32o_1 _16196_ (.A1(_02814_),
    .A2(_02817_),
    .A3(_02818_),
    .B1(_02676_),
    .B2(net297),
    .X(_01391_));
 sky130_fd_sc_hd__a21bo_1 _16197_ (.A1(net257),
    .A2(net261),
    .B1_N(_01822_),
    .X(_02819_));
 sky130_fd_sc_hd__or2_1 _16198_ (.A(net298),
    .B(_01822_),
    .X(_02820_));
 sky130_fd_sc_hd__a32o_1 _16199_ (.A1(_02814_),
    .A2(_02819_),
    .A3(_02820_),
    .B1(_02676_),
    .B2(net298),
    .X(_01392_));
 sky130_fd_sc_hd__nor2_1 _16200_ (.A(_03730_),
    .B(_02678_),
    .Y(_02821_));
 sky130_fd_sc_hd__nand2_1 _16201_ (.A(_02685_),
    .B(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__o211a_1 _16202_ (.A1(_03849_),
    .A2(_02821_),
    .B1(_02822_),
    .C1(_01821_),
    .X(_01393_));
 sky130_fd_sc_hd__nor2_1 _16203_ (.A(_03218_),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__nor2_1 _16204_ (.A(prefetched_high_word),
    .B(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__a41o_1 _16205_ (.A1(_03187_),
    .A2(net33),
    .A3(net44),
    .A4(_02823_),
    .B1(clear_prefetched_high_word),
    .X(_02825_));
 sky130_fd_sc_hd__nor3_1 _16206_ (.A(net299),
    .B(_02824_),
    .C(_02825_),
    .Y(_01394_));
 sky130_fd_sc_hd__and3_1 _16207_ (.A(_04156_),
    .B(_07898_),
    .C(_06863_),
    .X(_02826_));
 sky130_fd_sc_hd__a22o_1 _16208_ (.A1(_06082_),
    .A2(_06862_),
    .B1(_02826_),
    .B2(\decoded_rd[3] ),
    .X(_01395_));
 sky130_fd_sc_hd__a22o_1 _16209_ (.A1(_06081_),
    .A2(_06862_),
    .B1(_02826_),
    .B2(\decoded_rd[4] ),
    .X(_01396_));
 sky130_fd_sc_hd__and4_1 _16210_ (.A(_03187_),
    .B(_03198_),
    .C(_03215_),
    .D(_03217_),
    .X(_02827_));
 sky130_fd_sc_hd__nand2_1 _16211_ (.A(net33),
    .B(net44),
    .Y(_02828_));
 sky130_fd_sc_hd__o311ai_1 _16212_ (.A1(_03753_),
    .A2(_03223_),
    .A3(_02828_),
    .B1(_02821_),
    .C1(_01821_),
    .Y(_02829_));
 sky130_fd_sc_hd__a211o_2 _16213_ (.A1(_03218_),
    .A2(_02685_),
    .B1(_02827_),
    .C1(_02829_),
    .X(_02830_));
 sky130_fd_sc_hd__clkbuf_4 _16214_ (.A(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__mux2_1 _16215_ (.A0(net40),
    .A1(\mem_16bit_buffer[0] ),
    .S(_02831_),
    .X(_02832_));
 sky130_fd_sc_hd__clkbuf_1 _16216_ (.A(_02832_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _16217_ (.A0(net41),
    .A1(\mem_16bit_buffer[1] ),
    .S(_02831_),
    .X(_02833_));
 sky130_fd_sc_hd__clkbuf_1 _16218_ (.A(_02833_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _16219_ (.A0(net42),
    .A1(\mem_16bit_buffer[2] ),
    .S(_02831_),
    .X(_02834_));
 sky130_fd_sc_hd__clkbuf_1 _16220_ (.A(_02834_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _16221_ (.A0(net43),
    .A1(\mem_16bit_buffer[3] ),
    .S(_02831_),
    .X(_02835_));
 sky130_fd_sc_hd__clkbuf_1 _16222_ (.A(_02835_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _16223_ (.A0(net45),
    .A1(\mem_16bit_buffer[4] ),
    .S(_02831_),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_1 _16224_ (.A(_02836_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _16225_ (.A0(net46),
    .A1(\mem_16bit_buffer[5] ),
    .S(_02831_),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_1 _16226_ (.A(_02837_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _16227_ (.A0(net47),
    .A1(\mem_16bit_buffer[6] ),
    .S(_02831_),
    .X(_02838_));
 sky130_fd_sc_hd__clkbuf_1 _16228_ (.A(_02838_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _16229_ (.A0(net48),
    .A1(\mem_16bit_buffer[7] ),
    .S(_02831_),
    .X(_02839_));
 sky130_fd_sc_hd__clkbuf_1 _16230_ (.A(_02839_),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _16231_ (.A0(net49),
    .A1(\mem_16bit_buffer[8] ),
    .S(_02831_),
    .X(_02840_));
 sky130_fd_sc_hd__clkbuf_1 _16232_ (.A(_02840_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _16233_ (.A0(net50),
    .A1(\mem_16bit_buffer[9] ),
    .S(_02831_),
    .X(_02841_));
 sky130_fd_sc_hd__clkbuf_1 _16234_ (.A(_02841_),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _16235_ (.A0(net51),
    .A1(\mem_16bit_buffer[10] ),
    .S(_02830_),
    .X(_02842_));
 sky130_fd_sc_hd__clkbuf_1 _16236_ (.A(_02842_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _16237_ (.A0(net52),
    .A1(\mem_16bit_buffer[11] ),
    .S(_02830_),
    .X(_02843_));
 sky130_fd_sc_hd__clkbuf_1 _16238_ (.A(_02843_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _16239_ (.A0(net53),
    .A1(\mem_16bit_buffer[12] ),
    .S(_02830_),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _16240_ (.A(_02844_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _16241_ (.A0(net54),
    .A1(\mem_16bit_buffer[13] ),
    .S(_02830_),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_1 _16242_ (.A(_02845_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _16243_ (.A0(net56),
    .A1(\mem_16bit_buffer[14] ),
    .S(_02830_),
    .X(_02846_));
 sky130_fd_sc_hd__clkbuf_1 _16244_ (.A(_02846_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _16245_ (.A0(net57),
    .A1(\mem_16bit_buffer[15] ),
    .S(_02830_),
    .X(_02847_));
 sky130_fd_sc_hd__clkbuf_1 _16246_ (.A(_02847_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _16247_ (.A0(\mem_rdata_q[0] ),
    .A1(_03783_),
    .S(_03914_),
    .X(_02848_));
 sky130_fd_sc_hd__clkbuf_1 _16248_ (.A(_02848_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _16249_ (.A0(\mem_rdata_q[1] ),
    .A1(_03213_),
    .S(_03914_),
    .X(_02849_));
 sky130_fd_sc_hd__clkbuf_1 _16250_ (.A(_02849_),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _16251_ (.A0(\mem_rdata_q[2] ),
    .A1(_03864_),
    .S(_03914_),
    .X(_02850_));
 sky130_fd_sc_hd__clkbuf_1 _16252_ (.A(_02850_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _16253_ (.A0(\mem_rdata_q[3] ),
    .A1(_03810_),
    .S(_03914_),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_1 _16254_ (.A(_02851_),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _16255_ (.A0(\mem_rdata_q[4] ),
    .A1(_03885_),
    .S(_03914_),
    .X(_02852_));
 sky130_fd_sc_hd__clkbuf_1 _16256_ (.A(_02852_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _16257_ (.A0(\mem_rdata_q[5] ),
    .A1(_03895_),
    .S(_03914_),
    .X(_02853_));
 sky130_fd_sc_hd__clkbuf_1 _16258_ (.A(_02853_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _16259_ (.A0(\mem_rdata_q[6] ),
    .A1(_03878_),
    .S(_03914_),
    .X(_02854_));
 sky130_fd_sc_hd__clkbuf_1 _16260_ (.A(_02854_),
    .X(_01419_));
 sky130_fd_sc_hd__and2_1 _16261_ (.A(_07737_),
    .B(_03216_),
    .X(_02855_));
 sky130_fd_sc_hd__clkbuf_1 _16262_ (.A(_02855_),
    .X(_01420_));
 sky130_fd_sc_hd__a21o_1 _16263_ (.A1(_05941_),
    .A2(_07944_),
    .B1(_03292_),
    .X(_02856_));
 sky130_fd_sc_hd__and3_1 _16264_ (.A(\reg_next_pc[0] ),
    .B(_07778_),
    .C(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__clkbuf_1 _16265_ (.A(_02857_),
    .X(_01421_));
 sky130_fd_sc_hd__nand2_2 _16266_ (.A(_06346_),
    .B(_06823_),
    .Y(_02858_));
 sky130_fd_sc_hd__buf_6 _16267_ (.A(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__mux2_1 _16268_ (.A0(_06941_),
    .A1(\cpuregs.regs[15][0] ),
    .S(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__clkbuf_1 _16269_ (.A(_02860_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _16270_ (.A0(_06945_),
    .A1(\cpuregs.regs[15][1] ),
    .S(_02859_),
    .X(_02861_));
 sky130_fd_sc_hd__clkbuf_1 _16271_ (.A(_02861_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _16272_ (.A0(_06947_),
    .A1(\cpuregs.regs[15][2] ),
    .S(_02859_),
    .X(_02862_));
 sky130_fd_sc_hd__clkbuf_1 _16273_ (.A(_02862_),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _16274_ (.A0(_06949_),
    .A1(\cpuregs.regs[15][3] ),
    .S(_02859_),
    .X(_02863_));
 sky130_fd_sc_hd__clkbuf_1 _16275_ (.A(_02863_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _16276_ (.A0(_06951_),
    .A1(\cpuregs.regs[15][4] ),
    .S(_02859_),
    .X(_02864_));
 sky130_fd_sc_hd__clkbuf_1 _16277_ (.A(_02864_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _16278_ (.A0(_06953_),
    .A1(\cpuregs.regs[15][5] ),
    .S(_02859_),
    .X(_02865_));
 sky130_fd_sc_hd__clkbuf_1 _16279_ (.A(_02865_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _16280_ (.A0(_06955_),
    .A1(\cpuregs.regs[15][6] ),
    .S(_02859_),
    .X(_02866_));
 sky130_fd_sc_hd__clkbuf_1 _16281_ (.A(_02866_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _16282_ (.A0(_06957_),
    .A1(\cpuregs.regs[15][7] ),
    .S(_02859_),
    .X(_02867_));
 sky130_fd_sc_hd__clkbuf_1 _16283_ (.A(_02867_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _16284_ (.A0(_06959_),
    .A1(\cpuregs.regs[15][8] ),
    .S(_02859_),
    .X(_02868_));
 sky130_fd_sc_hd__clkbuf_1 _16285_ (.A(_02868_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _16286_ (.A0(_06961_),
    .A1(\cpuregs.regs[15][9] ),
    .S(_02859_),
    .X(_02869_));
 sky130_fd_sc_hd__clkbuf_1 _16287_ (.A(_02869_),
    .X(_01431_));
 sky130_fd_sc_hd__buf_6 _16288_ (.A(_02858_),
    .X(_02870_));
 sky130_fd_sc_hd__mux2_1 _16289_ (.A0(_06963_),
    .A1(\cpuregs.regs[15][10] ),
    .S(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__clkbuf_1 _16290_ (.A(_02871_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _16291_ (.A0(_06966_),
    .A1(\cpuregs.regs[15][11] ),
    .S(_02870_),
    .X(_02872_));
 sky130_fd_sc_hd__clkbuf_1 _16292_ (.A(_02872_),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _16293_ (.A0(_06968_),
    .A1(\cpuregs.regs[15][12] ),
    .S(_02870_),
    .X(_02873_));
 sky130_fd_sc_hd__clkbuf_1 _16294_ (.A(_02873_),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _16295_ (.A0(_06970_),
    .A1(\cpuregs.regs[15][13] ),
    .S(_02870_),
    .X(_02874_));
 sky130_fd_sc_hd__clkbuf_1 _16296_ (.A(_02874_),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _16297_ (.A0(_06972_),
    .A1(\cpuregs.regs[15][14] ),
    .S(_02870_),
    .X(_02875_));
 sky130_fd_sc_hd__clkbuf_1 _16298_ (.A(_02875_),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _16299_ (.A0(_06974_),
    .A1(\cpuregs.regs[15][15] ),
    .S(_02870_),
    .X(_02876_));
 sky130_fd_sc_hd__clkbuf_1 _16300_ (.A(_02876_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _16301_ (.A0(_06976_),
    .A1(\cpuregs.regs[15][16] ),
    .S(_02870_),
    .X(_02877_));
 sky130_fd_sc_hd__clkbuf_1 _16302_ (.A(_02877_),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _16303_ (.A0(_06978_),
    .A1(\cpuregs.regs[15][17] ),
    .S(_02870_),
    .X(_02878_));
 sky130_fd_sc_hd__clkbuf_1 _16304_ (.A(_02878_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _16305_ (.A0(_06980_),
    .A1(\cpuregs.regs[15][18] ),
    .S(_02870_),
    .X(_02879_));
 sky130_fd_sc_hd__clkbuf_1 _16306_ (.A(_02879_),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _16307_ (.A0(_06982_),
    .A1(\cpuregs.regs[15][19] ),
    .S(_02870_),
    .X(_02880_));
 sky130_fd_sc_hd__clkbuf_1 _16308_ (.A(_02880_),
    .X(_01441_));
 sky130_fd_sc_hd__clkbuf_8 _16309_ (.A(_02858_),
    .X(_02881_));
 sky130_fd_sc_hd__mux2_1 _16310_ (.A0(_06984_),
    .A1(\cpuregs.regs[15][20] ),
    .S(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__clkbuf_1 _16311_ (.A(_02882_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _16312_ (.A0(_06987_),
    .A1(\cpuregs.regs[15][21] ),
    .S(_02881_),
    .X(_02883_));
 sky130_fd_sc_hd__clkbuf_1 _16313_ (.A(_02883_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _16314_ (.A0(_06989_),
    .A1(\cpuregs.regs[15][22] ),
    .S(_02881_),
    .X(_02884_));
 sky130_fd_sc_hd__clkbuf_1 _16315_ (.A(_02884_),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _16316_ (.A0(_06991_),
    .A1(\cpuregs.regs[15][23] ),
    .S(_02881_),
    .X(_02885_));
 sky130_fd_sc_hd__clkbuf_1 _16317_ (.A(_02885_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _16318_ (.A0(_06993_),
    .A1(\cpuregs.regs[15][24] ),
    .S(_02881_),
    .X(_02886_));
 sky130_fd_sc_hd__clkbuf_1 _16319_ (.A(_02886_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _16320_ (.A0(_06995_),
    .A1(\cpuregs.regs[15][25] ),
    .S(_02881_),
    .X(_02887_));
 sky130_fd_sc_hd__clkbuf_1 _16321_ (.A(_02887_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _16322_ (.A0(_06997_),
    .A1(\cpuregs.regs[15][26] ),
    .S(_02881_),
    .X(_02888_));
 sky130_fd_sc_hd__clkbuf_1 _16323_ (.A(_02888_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _16324_ (.A0(_06999_),
    .A1(\cpuregs.regs[15][27] ),
    .S(_02881_),
    .X(_02889_));
 sky130_fd_sc_hd__clkbuf_1 _16325_ (.A(_02889_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _16326_ (.A0(_07001_),
    .A1(\cpuregs.regs[15][28] ),
    .S(_02881_),
    .X(_02890_));
 sky130_fd_sc_hd__clkbuf_1 _16327_ (.A(_02890_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _16328_ (.A0(_07003_),
    .A1(\cpuregs.regs[15][29] ),
    .S(_02881_),
    .X(_02891_));
 sky130_fd_sc_hd__clkbuf_1 _16329_ (.A(_02891_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _16330_ (.A0(_07005_),
    .A1(\cpuregs.regs[15][30] ),
    .S(_02858_),
    .X(_02892_));
 sky130_fd_sc_hd__clkbuf_1 _16331_ (.A(_02892_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _16332_ (.A0(_07007_),
    .A1(\cpuregs.regs[15][31] ),
    .S(_02858_),
    .X(_02893_));
 sky130_fd_sc_hd__clkbuf_1 _16333_ (.A(_02893_),
    .X(_01453_));
 sky130_fd_sc_hd__and4bb_4 _16334_ (.A_N(\cpuregs.waddr[2] ),
    .B_N(_06082_),
    .C(_06083_),
    .D(_06081_),
    .X(_02894_));
 sky130_fd_sc_hd__nand2_4 _16335_ (.A(_06383_),
    .B(_02894_),
    .Y(_02895_));
 sky130_fd_sc_hd__clkbuf_8 _16336_ (.A(_02895_),
    .X(_02896_));
 sky130_fd_sc_hd__mux2_1 _16337_ (.A0(_06941_),
    .A1(\cpuregs.regs[16][0] ),
    .S(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__clkbuf_1 _16338_ (.A(_02897_),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _16339_ (.A0(_06945_),
    .A1(\cpuregs.regs[16][1] ),
    .S(_02896_),
    .X(_02898_));
 sky130_fd_sc_hd__clkbuf_1 _16340_ (.A(_02898_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _16341_ (.A0(_06947_),
    .A1(\cpuregs.regs[16][2] ),
    .S(_02896_),
    .X(_02899_));
 sky130_fd_sc_hd__clkbuf_1 _16342_ (.A(_02899_),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _16343_ (.A0(_06949_),
    .A1(\cpuregs.regs[16][3] ),
    .S(_02896_),
    .X(_02900_));
 sky130_fd_sc_hd__clkbuf_1 _16344_ (.A(_02900_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _16345_ (.A0(_06951_),
    .A1(\cpuregs.regs[16][4] ),
    .S(_02896_),
    .X(_02901_));
 sky130_fd_sc_hd__clkbuf_1 _16346_ (.A(_02901_),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _16347_ (.A0(_06953_),
    .A1(\cpuregs.regs[16][5] ),
    .S(_02896_),
    .X(_02902_));
 sky130_fd_sc_hd__clkbuf_1 _16348_ (.A(_02902_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _16349_ (.A0(_06955_),
    .A1(\cpuregs.regs[16][6] ),
    .S(_02896_),
    .X(_02903_));
 sky130_fd_sc_hd__clkbuf_1 _16350_ (.A(_02903_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _16351_ (.A0(_06957_),
    .A1(\cpuregs.regs[16][7] ),
    .S(_02896_),
    .X(_02904_));
 sky130_fd_sc_hd__clkbuf_1 _16352_ (.A(_02904_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _16353_ (.A0(_06959_),
    .A1(\cpuregs.regs[16][8] ),
    .S(_02896_),
    .X(_02905_));
 sky130_fd_sc_hd__clkbuf_1 _16354_ (.A(_02905_),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _16355_ (.A0(_06961_),
    .A1(\cpuregs.regs[16][9] ),
    .S(_02896_),
    .X(_02906_));
 sky130_fd_sc_hd__clkbuf_1 _16356_ (.A(_02906_),
    .X(_01463_));
 sky130_fd_sc_hd__clkbuf_8 _16357_ (.A(_02895_),
    .X(_02907_));
 sky130_fd_sc_hd__mux2_1 _16358_ (.A0(_06963_),
    .A1(\cpuregs.regs[16][10] ),
    .S(_02907_),
    .X(_02908_));
 sky130_fd_sc_hd__clkbuf_1 _16359_ (.A(_02908_),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _16360_ (.A0(_06966_),
    .A1(\cpuregs.regs[16][11] ),
    .S(_02907_),
    .X(_02909_));
 sky130_fd_sc_hd__clkbuf_1 _16361_ (.A(_02909_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _16362_ (.A0(_06968_),
    .A1(\cpuregs.regs[16][12] ),
    .S(_02907_),
    .X(_02910_));
 sky130_fd_sc_hd__clkbuf_1 _16363_ (.A(_02910_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _16364_ (.A0(_06970_),
    .A1(\cpuregs.regs[16][13] ),
    .S(_02907_),
    .X(_02911_));
 sky130_fd_sc_hd__clkbuf_1 _16365_ (.A(_02911_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _16366_ (.A0(_06972_),
    .A1(\cpuregs.regs[16][14] ),
    .S(_02907_),
    .X(_02912_));
 sky130_fd_sc_hd__clkbuf_1 _16367_ (.A(_02912_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _16368_ (.A0(_06974_),
    .A1(\cpuregs.regs[16][15] ),
    .S(_02907_),
    .X(_02913_));
 sky130_fd_sc_hd__clkbuf_1 _16369_ (.A(_02913_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _16370_ (.A0(_06976_),
    .A1(\cpuregs.regs[16][16] ),
    .S(_02907_),
    .X(_02914_));
 sky130_fd_sc_hd__clkbuf_1 _16371_ (.A(_02914_),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _16372_ (.A0(_06978_),
    .A1(\cpuregs.regs[16][17] ),
    .S(_02907_),
    .X(_02915_));
 sky130_fd_sc_hd__clkbuf_1 _16373_ (.A(_02915_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _16374_ (.A0(_06980_),
    .A1(\cpuregs.regs[16][18] ),
    .S(_02907_),
    .X(_02916_));
 sky130_fd_sc_hd__clkbuf_1 _16375_ (.A(_02916_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _16376_ (.A0(_06982_),
    .A1(\cpuregs.regs[16][19] ),
    .S(_02907_),
    .X(_02917_));
 sky130_fd_sc_hd__clkbuf_1 _16377_ (.A(_02917_),
    .X(_01473_));
 sky130_fd_sc_hd__buf_6 _16378_ (.A(_02895_),
    .X(_02918_));
 sky130_fd_sc_hd__mux2_1 _16379_ (.A0(_06984_),
    .A1(\cpuregs.regs[16][20] ),
    .S(_02918_),
    .X(_02919_));
 sky130_fd_sc_hd__clkbuf_1 _16380_ (.A(_02919_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _16381_ (.A0(_06987_),
    .A1(\cpuregs.regs[16][21] ),
    .S(_02918_),
    .X(_02920_));
 sky130_fd_sc_hd__clkbuf_1 _16382_ (.A(_02920_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _16383_ (.A0(_06989_),
    .A1(\cpuregs.regs[16][22] ),
    .S(_02918_),
    .X(_02921_));
 sky130_fd_sc_hd__clkbuf_1 _16384_ (.A(_02921_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _16385_ (.A0(_06991_),
    .A1(\cpuregs.regs[16][23] ),
    .S(_02918_),
    .X(_02922_));
 sky130_fd_sc_hd__clkbuf_1 _16386_ (.A(_02922_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _16387_ (.A0(_06993_),
    .A1(\cpuregs.regs[16][24] ),
    .S(_02918_),
    .X(_02923_));
 sky130_fd_sc_hd__clkbuf_1 _16388_ (.A(_02923_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _16389_ (.A0(_06995_),
    .A1(\cpuregs.regs[16][25] ),
    .S(_02918_),
    .X(_02924_));
 sky130_fd_sc_hd__clkbuf_1 _16390_ (.A(_02924_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _16391_ (.A0(_06997_),
    .A1(\cpuregs.regs[16][26] ),
    .S(_02918_),
    .X(_02925_));
 sky130_fd_sc_hd__clkbuf_1 _16392_ (.A(_02925_),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _16393_ (.A0(_06999_),
    .A1(\cpuregs.regs[16][27] ),
    .S(_02918_),
    .X(_02926_));
 sky130_fd_sc_hd__clkbuf_1 _16394_ (.A(_02926_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _16395_ (.A0(_07001_),
    .A1(\cpuregs.regs[16][28] ),
    .S(_02918_),
    .X(_02927_));
 sky130_fd_sc_hd__clkbuf_1 _16396_ (.A(_02927_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _16397_ (.A0(_07003_),
    .A1(\cpuregs.regs[16][29] ),
    .S(_02918_),
    .X(_02928_));
 sky130_fd_sc_hd__clkbuf_1 _16398_ (.A(_02928_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _16399_ (.A0(_07005_),
    .A1(\cpuregs.regs[16][30] ),
    .S(_02895_),
    .X(_02929_));
 sky130_fd_sc_hd__clkbuf_1 _16400_ (.A(_02929_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _16401_ (.A0(_07007_),
    .A1(\cpuregs.regs[16][31] ),
    .S(_02895_),
    .X(_02930_));
 sky130_fd_sc_hd__clkbuf_1 _16402_ (.A(_02930_),
    .X(_01485_));
 sky130_fd_sc_hd__nand2_4 _16403_ (.A(_06422_),
    .B(_06713_),
    .Y(_02931_));
 sky130_fd_sc_hd__buf_6 _16404_ (.A(_02931_),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_1 _16405_ (.A0(_06941_),
    .A1(\cpuregs.regs[29][0] ),
    .S(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__clkbuf_1 _16406_ (.A(_02933_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _16407_ (.A0(_06945_),
    .A1(\cpuregs.regs[29][1] ),
    .S(_02932_),
    .X(_02934_));
 sky130_fd_sc_hd__clkbuf_1 _16408_ (.A(_02934_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _16409_ (.A0(_06947_),
    .A1(\cpuregs.regs[29][2] ),
    .S(_02932_),
    .X(_02935_));
 sky130_fd_sc_hd__clkbuf_1 _16410_ (.A(_02935_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _16411_ (.A0(_06949_),
    .A1(\cpuregs.regs[29][3] ),
    .S(_02932_),
    .X(_02936_));
 sky130_fd_sc_hd__clkbuf_1 _16412_ (.A(_02936_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _16413_ (.A0(_06951_),
    .A1(\cpuregs.regs[29][4] ),
    .S(_02932_),
    .X(_02937_));
 sky130_fd_sc_hd__clkbuf_1 _16414_ (.A(_02937_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _16415_ (.A0(_06953_),
    .A1(\cpuregs.regs[29][5] ),
    .S(_02932_),
    .X(_02938_));
 sky130_fd_sc_hd__clkbuf_1 _16416_ (.A(_02938_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _16417_ (.A0(_06955_),
    .A1(\cpuregs.regs[29][6] ),
    .S(_02932_),
    .X(_02939_));
 sky130_fd_sc_hd__clkbuf_1 _16418_ (.A(_02939_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _16419_ (.A0(_06957_),
    .A1(\cpuregs.regs[29][7] ),
    .S(_02932_),
    .X(_02940_));
 sky130_fd_sc_hd__clkbuf_1 _16420_ (.A(_02940_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _16421_ (.A0(_06959_),
    .A1(\cpuregs.regs[29][8] ),
    .S(_02932_),
    .X(_02941_));
 sky130_fd_sc_hd__clkbuf_1 _16422_ (.A(_02941_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _16423_ (.A0(_06961_),
    .A1(\cpuregs.regs[29][9] ),
    .S(_02932_),
    .X(_02942_));
 sky130_fd_sc_hd__clkbuf_1 _16424_ (.A(_02942_),
    .X(_01495_));
 sky130_fd_sc_hd__buf_6 _16425_ (.A(_02931_),
    .X(_02943_));
 sky130_fd_sc_hd__mux2_1 _16426_ (.A0(_06963_),
    .A1(\cpuregs.regs[29][10] ),
    .S(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__clkbuf_1 _16427_ (.A(_02944_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _16428_ (.A0(_06966_),
    .A1(\cpuregs.regs[29][11] ),
    .S(_02943_),
    .X(_02945_));
 sky130_fd_sc_hd__clkbuf_1 _16429_ (.A(_02945_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _16430_ (.A0(_06968_),
    .A1(\cpuregs.regs[29][12] ),
    .S(_02943_),
    .X(_02946_));
 sky130_fd_sc_hd__clkbuf_1 _16431_ (.A(_02946_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _16432_ (.A0(_06970_),
    .A1(\cpuregs.regs[29][13] ),
    .S(_02943_),
    .X(_02947_));
 sky130_fd_sc_hd__clkbuf_1 _16433_ (.A(_02947_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _16434_ (.A0(_06972_),
    .A1(\cpuregs.regs[29][14] ),
    .S(_02943_),
    .X(_02948_));
 sky130_fd_sc_hd__clkbuf_1 _16435_ (.A(_02948_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _16436_ (.A0(_06974_),
    .A1(\cpuregs.regs[29][15] ),
    .S(_02943_),
    .X(_02949_));
 sky130_fd_sc_hd__clkbuf_1 _16437_ (.A(_02949_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _16438_ (.A0(_06976_),
    .A1(\cpuregs.regs[29][16] ),
    .S(_02943_),
    .X(_02950_));
 sky130_fd_sc_hd__clkbuf_1 _16439_ (.A(_02950_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _16440_ (.A0(_06978_),
    .A1(\cpuregs.regs[29][17] ),
    .S(_02943_),
    .X(_02951_));
 sky130_fd_sc_hd__clkbuf_1 _16441_ (.A(_02951_),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _16442_ (.A0(_06980_),
    .A1(\cpuregs.regs[29][18] ),
    .S(_02943_),
    .X(_02952_));
 sky130_fd_sc_hd__clkbuf_1 _16443_ (.A(_02952_),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _16444_ (.A0(_06982_),
    .A1(\cpuregs.regs[29][19] ),
    .S(_02943_),
    .X(_02953_));
 sky130_fd_sc_hd__clkbuf_1 _16445_ (.A(_02953_),
    .X(_01505_));
 sky130_fd_sc_hd__buf_6 _16446_ (.A(_02931_),
    .X(_02954_));
 sky130_fd_sc_hd__mux2_1 _16447_ (.A0(_06984_),
    .A1(\cpuregs.regs[29][20] ),
    .S(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__clkbuf_1 _16448_ (.A(_02955_),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _16449_ (.A0(_06987_),
    .A1(\cpuregs.regs[29][21] ),
    .S(_02954_),
    .X(_02956_));
 sky130_fd_sc_hd__clkbuf_1 _16450_ (.A(_02956_),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _16451_ (.A0(_06989_),
    .A1(\cpuregs.regs[29][22] ),
    .S(_02954_),
    .X(_02957_));
 sky130_fd_sc_hd__clkbuf_1 _16452_ (.A(_02957_),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _16453_ (.A0(_06991_),
    .A1(\cpuregs.regs[29][23] ),
    .S(_02954_),
    .X(_02958_));
 sky130_fd_sc_hd__clkbuf_1 _16454_ (.A(_02958_),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _16455_ (.A0(_06993_),
    .A1(\cpuregs.regs[29][24] ),
    .S(_02954_),
    .X(_02959_));
 sky130_fd_sc_hd__clkbuf_1 _16456_ (.A(_02959_),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _16457_ (.A0(_06995_),
    .A1(\cpuregs.regs[29][25] ),
    .S(_02954_),
    .X(_02960_));
 sky130_fd_sc_hd__clkbuf_1 _16458_ (.A(_02960_),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _16459_ (.A0(_06997_),
    .A1(\cpuregs.regs[29][26] ),
    .S(_02954_),
    .X(_02961_));
 sky130_fd_sc_hd__clkbuf_1 _16460_ (.A(_02961_),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _16461_ (.A0(_06999_),
    .A1(\cpuregs.regs[29][27] ),
    .S(_02954_),
    .X(_02962_));
 sky130_fd_sc_hd__clkbuf_1 _16462_ (.A(_02962_),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _16463_ (.A0(_07001_),
    .A1(\cpuregs.regs[29][28] ),
    .S(_02954_),
    .X(_02963_));
 sky130_fd_sc_hd__clkbuf_1 _16464_ (.A(_02963_),
    .X(_01514_));
 sky130_fd_sc_hd__mux2_1 _16465_ (.A0(_07003_),
    .A1(\cpuregs.regs[29][29] ),
    .S(_02954_),
    .X(_02964_));
 sky130_fd_sc_hd__clkbuf_1 _16466_ (.A(_02964_),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _16467_ (.A0(_07005_),
    .A1(\cpuregs.regs[29][30] ),
    .S(_02931_),
    .X(_02965_));
 sky130_fd_sc_hd__clkbuf_1 _16468_ (.A(_02965_),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _16469_ (.A0(_07007_),
    .A1(\cpuregs.regs[29][31] ),
    .S(_02931_),
    .X(_02966_));
 sky130_fd_sc_hd__clkbuf_1 _16470_ (.A(_02966_),
    .X(_01517_));
 sky130_fd_sc_hd__and4bb_4 _16471_ (.A_N(\cpuregs.waddr[2] ),
    .B_N(_06082_),
    .C(_06601_),
    .D(_06081_),
    .X(_02967_));
 sky130_fd_sc_hd__buf_6 _16472_ (.A(_02967_),
    .X(_02968_));
 sky130_fd_sc_hd__mux2_1 _16473_ (.A0(\cpuregs.regs[17][0] ),
    .A1(_06531_),
    .S(_02968_),
    .X(_02969_));
 sky130_fd_sc_hd__clkbuf_1 _16474_ (.A(_02969_),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _16475_ (.A0(\cpuregs.regs[17][1] ),
    .A1(_06536_),
    .S(_02968_),
    .X(_02970_));
 sky130_fd_sc_hd__clkbuf_1 _16476_ (.A(_02970_),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _16477_ (.A0(\cpuregs.regs[17][2] ),
    .A1(_06538_),
    .S(_02968_),
    .X(_02971_));
 sky130_fd_sc_hd__clkbuf_1 _16478_ (.A(_02971_),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _16479_ (.A0(\cpuregs.regs[17][3] ),
    .A1(_06540_),
    .S(_02968_),
    .X(_02972_));
 sky130_fd_sc_hd__clkbuf_1 _16480_ (.A(_02972_),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _16481_ (.A0(\cpuregs.regs[17][4] ),
    .A1(_06542_),
    .S(_02968_),
    .X(_02973_));
 sky130_fd_sc_hd__clkbuf_1 _16482_ (.A(_02973_),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _16483_ (.A0(\cpuregs.regs[17][5] ),
    .A1(_06544_),
    .S(_02968_),
    .X(_02974_));
 sky130_fd_sc_hd__clkbuf_1 _16484_ (.A(_02974_),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _16485_ (.A0(\cpuregs.regs[17][6] ),
    .A1(_06546_),
    .S(_02968_),
    .X(_02975_));
 sky130_fd_sc_hd__clkbuf_1 _16486_ (.A(_02975_),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _16487_ (.A0(\cpuregs.regs[17][7] ),
    .A1(_06548_),
    .S(_02968_),
    .X(_02976_));
 sky130_fd_sc_hd__clkbuf_1 _16488_ (.A(_02976_),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _16489_ (.A0(\cpuregs.regs[17][8] ),
    .A1(_06550_),
    .S(_02968_),
    .X(_02977_));
 sky130_fd_sc_hd__clkbuf_1 _16490_ (.A(_02977_),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _16491_ (.A0(\cpuregs.regs[17][9] ),
    .A1(_06552_),
    .S(_02968_),
    .X(_02978_));
 sky130_fd_sc_hd__clkbuf_1 _16492_ (.A(_02978_),
    .X(_01527_));
 sky130_fd_sc_hd__clkbuf_8 _16493_ (.A(_02967_),
    .X(_02979_));
 sky130_fd_sc_hd__mux2_1 _16494_ (.A0(\cpuregs.regs[17][10] ),
    .A1(_06554_),
    .S(_02979_),
    .X(_02980_));
 sky130_fd_sc_hd__clkbuf_1 _16495_ (.A(_02980_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _16496_ (.A0(\cpuregs.regs[17][11] ),
    .A1(_06557_),
    .S(_02979_),
    .X(_02981_));
 sky130_fd_sc_hd__clkbuf_1 _16497_ (.A(_02981_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _16498_ (.A0(\cpuregs.regs[17][12] ),
    .A1(_06559_),
    .S(_02979_),
    .X(_02982_));
 sky130_fd_sc_hd__clkbuf_1 _16499_ (.A(_02982_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _16500_ (.A0(\cpuregs.regs[17][13] ),
    .A1(_06561_),
    .S(_02979_),
    .X(_02983_));
 sky130_fd_sc_hd__clkbuf_1 _16501_ (.A(_02983_),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _16502_ (.A0(\cpuregs.regs[17][14] ),
    .A1(_06563_),
    .S(_02979_),
    .X(_02984_));
 sky130_fd_sc_hd__clkbuf_1 _16503_ (.A(_02984_),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _16504_ (.A0(\cpuregs.regs[17][15] ),
    .A1(_06565_),
    .S(_02979_),
    .X(_02985_));
 sky130_fd_sc_hd__clkbuf_1 _16505_ (.A(_02985_),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _16506_ (.A0(\cpuregs.regs[17][16] ),
    .A1(_06567_),
    .S(_02979_),
    .X(_02986_));
 sky130_fd_sc_hd__clkbuf_1 _16507_ (.A(_02986_),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _16508_ (.A0(\cpuregs.regs[17][17] ),
    .A1(_06569_),
    .S(_02979_),
    .X(_02987_));
 sky130_fd_sc_hd__clkbuf_1 _16509_ (.A(_02987_),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _16510_ (.A0(\cpuregs.regs[17][18] ),
    .A1(_06571_),
    .S(_02979_),
    .X(_02988_));
 sky130_fd_sc_hd__clkbuf_1 _16511_ (.A(_02988_),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _16512_ (.A0(\cpuregs.regs[17][19] ),
    .A1(_06573_),
    .S(_02979_),
    .X(_02989_));
 sky130_fd_sc_hd__clkbuf_1 _16513_ (.A(_02989_),
    .X(_01537_));
 sky130_fd_sc_hd__clkbuf_8 _16514_ (.A(_02967_),
    .X(_02990_));
 sky130_fd_sc_hd__mux2_1 _16515_ (.A0(\cpuregs.regs[17][20] ),
    .A1(_06575_),
    .S(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__clkbuf_1 _16516_ (.A(_02991_),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _16517_ (.A0(\cpuregs.regs[17][21] ),
    .A1(_06578_),
    .S(_02990_),
    .X(_02992_));
 sky130_fd_sc_hd__clkbuf_1 _16518_ (.A(_02992_),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _16519_ (.A0(\cpuregs.regs[17][22] ),
    .A1(_06580_),
    .S(_02990_),
    .X(_02993_));
 sky130_fd_sc_hd__clkbuf_1 _16520_ (.A(_02993_),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _16521_ (.A0(\cpuregs.regs[17][23] ),
    .A1(_06582_),
    .S(_02990_),
    .X(_02994_));
 sky130_fd_sc_hd__clkbuf_1 _16522_ (.A(_02994_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _16523_ (.A0(\cpuregs.regs[17][24] ),
    .A1(_06584_),
    .S(_02990_),
    .X(_02995_));
 sky130_fd_sc_hd__clkbuf_1 _16524_ (.A(_02995_),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _16525_ (.A0(\cpuregs.regs[17][25] ),
    .A1(_06586_),
    .S(_02990_),
    .X(_02996_));
 sky130_fd_sc_hd__clkbuf_1 _16526_ (.A(_02996_),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _16527_ (.A0(\cpuregs.regs[17][26] ),
    .A1(_06588_),
    .S(_02990_),
    .X(_02997_));
 sky130_fd_sc_hd__clkbuf_1 _16528_ (.A(_02997_),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _16529_ (.A0(\cpuregs.regs[17][27] ),
    .A1(_06590_),
    .S(_02990_),
    .X(_02998_));
 sky130_fd_sc_hd__clkbuf_1 _16530_ (.A(_02998_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _16531_ (.A0(\cpuregs.regs[17][28] ),
    .A1(_06592_),
    .S(_02990_),
    .X(_02999_));
 sky130_fd_sc_hd__clkbuf_1 _16532_ (.A(_02999_),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _16533_ (.A0(\cpuregs.regs[17][29] ),
    .A1(_06594_),
    .S(_02990_),
    .X(_03000_));
 sky130_fd_sc_hd__clkbuf_1 _16534_ (.A(_03000_),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _16535_ (.A0(\cpuregs.regs[17][30] ),
    .A1(_06596_),
    .S(_02967_),
    .X(_03001_));
 sky130_fd_sc_hd__clkbuf_1 _16536_ (.A(_03001_),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _16537_ (.A0(\cpuregs.regs[17][31] ),
    .A1(_06598_),
    .S(_02967_),
    .X(_03002_));
 sky130_fd_sc_hd__clkbuf_1 _16538_ (.A(_03002_),
    .X(_01549_));
 sky130_fd_sc_hd__nand2_4 _16539_ (.A(_06080_),
    .B(_02894_),
    .Y(_03003_));
 sky130_fd_sc_hd__clkbuf_8 _16540_ (.A(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__mux2_1 _16541_ (.A0(_06941_),
    .A1(\cpuregs.regs[18][0] ),
    .S(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__clkbuf_1 _16542_ (.A(_03005_),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _16543_ (.A0(_06945_),
    .A1(\cpuregs.regs[18][1] ),
    .S(_03004_),
    .X(_03006_));
 sky130_fd_sc_hd__clkbuf_1 _16544_ (.A(_03006_),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _16545_ (.A0(_06947_),
    .A1(\cpuregs.regs[18][2] ),
    .S(_03004_),
    .X(_03007_));
 sky130_fd_sc_hd__clkbuf_1 _16546_ (.A(_03007_),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _16547_ (.A0(_06949_),
    .A1(\cpuregs.regs[18][3] ),
    .S(_03004_),
    .X(_03008_));
 sky130_fd_sc_hd__clkbuf_1 _16548_ (.A(_03008_),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _16549_ (.A0(_06951_),
    .A1(\cpuregs.regs[18][4] ),
    .S(_03004_),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_1 _16550_ (.A(_03009_),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _16551_ (.A0(_06953_),
    .A1(\cpuregs.regs[18][5] ),
    .S(_03004_),
    .X(_03010_));
 sky130_fd_sc_hd__clkbuf_1 _16552_ (.A(_03010_),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _16553_ (.A0(_06955_),
    .A1(\cpuregs.regs[18][6] ),
    .S(_03004_),
    .X(_03011_));
 sky130_fd_sc_hd__clkbuf_1 _16554_ (.A(_03011_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _16555_ (.A0(_06957_),
    .A1(\cpuregs.regs[18][7] ),
    .S(_03004_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_1 _16556_ (.A(_03012_),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _16557_ (.A0(_06959_),
    .A1(\cpuregs.regs[18][8] ),
    .S(_03004_),
    .X(_03013_));
 sky130_fd_sc_hd__clkbuf_1 _16558_ (.A(_03013_),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _16559_ (.A0(_06961_),
    .A1(\cpuregs.regs[18][9] ),
    .S(_03004_),
    .X(_03014_));
 sky130_fd_sc_hd__clkbuf_1 _16560_ (.A(_03014_),
    .X(_01559_));
 sky130_fd_sc_hd__clkbuf_8 _16561_ (.A(_03003_),
    .X(_03015_));
 sky130_fd_sc_hd__mux2_1 _16562_ (.A0(_06963_),
    .A1(\cpuregs.regs[18][10] ),
    .S(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__clkbuf_1 _16563_ (.A(_03016_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _16564_ (.A0(_06966_),
    .A1(\cpuregs.regs[18][11] ),
    .S(_03015_),
    .X(_03017_));
 sky130_fd_sc_hd__clkbuf_1 _16565_ (.A(_03017_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _16566_ (.A0(_06968_),
    .A1(\cpuregs.regs[18][12] ),
    .S(_03015_),
    .X(_03018_));
 sky130_fd_sc_hd__clkbuf_1 _16567_ (.A(_03018_),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _16568_ (.A0(_06970_),
    .A1(\cpuregs.regs[18][13] ),
    .S(_03015_),
    .X(_03019_));
 sky130_fd_sc_hd__clkbuf_1 _16569_ (.A(_03019_),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _16570_ (.A0(_06972_),
    .A1(\cpuregs.regs[18][14] ),
    .S(_03015_),
    .X(_03020_));
 sky130_fd_sc_hd__clkbuf_1 _16571_ (.A(_03020_),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _16572_ (.A0(_06974_),
    .A1(\cpuregs.regs[18][15] ),
    .S(_03015_),
    .X(_03021_));
 sky130_fd_sc_hd__clkbuf_1 _16573_ (.A(_03021_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _16574_ (.A0(_06976_),
    .A1(\cpuregs.regs[18][16] ),
    .S(_03015_),
    .X(_03022_));
 sky130_fd_sc_hd__clkbuf_1 _16575_ (.A(_03022_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _16576_ (.A0(_06978_),
    .A1(\cpuregs.regs[18][17] ),
    .S(_03015_),
    .X(_03023_));
 sky130_fd_sc_hd__clkbuf_1 _16577_ (.A(_03023_),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _16578_ (.A0(_06980_),
    .A1(\cpuregs.regs[18][18] ),
    .S(_03015_),
    .X(_03024_));
 sky130_fd_sc_hd__clkbuf_1 _16579_ (.A(_03024_),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _16580_ (.A0(_06982_),
    .A1(\cpuregs.regs[18][19] ),
    .S(_03015_),
    .X(_03025_));
 sky130_fd_sc_hd__clkbuf_1 _16581_ (.A(_03025_),
    .X(_01569_));
 sky130_fd_sc_hd__buf_6 _16582_ (.A(_03003_),
    .X(_03026_));
 sky130_fd_sc_hd__mux2_1 _16583_ (.A0(_06984_),
    .A1(\cpuregs.regs[18][20] ),
    .S(_03026_),
    .X(_03027_));
 sky130_fd_sc_hd__clkbuf_1 _16584_ (.A(_03027_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _16585_ (.A0(_06987_),
    .A1(\cpuregs.regs[18][21] ),
    .S(_03026_),
    .X(_03028_));
 sky130_fd_sc_hd__clkbuf_1 _16586_ (.A(_03028_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _16587_ (.A0(_06989_),
    .A1(\cpuregs.regs[18][22] ),
    .S(_03026_),
    .X(_03029_));
 sky130_fd_sc_hd__clkbuf_1 _16588_ (.A(_03029_),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _16589_ (.A0(_06991_),
    .A1(\cpuregs.regs[18][23] ),
    .S(_03026_),
    .X(_03030_));
 sky130_fd_sc_hd__clkbuf_1 _16590_ (.A(_03030_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _16591_ (.A0(_06993_),
    .A1(\cpuregs.regs[18][24] ),
    .S(_03026_),
    .X(_03031_));
 sky130_fd_sc_hd__clkbuf_1 _16592_ (.A(_03031_),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _16593_ (.A0(_06995_),
    .A1(\cpuregs.regs[18][25] ),
    .S(_03026_),
    .X(_03032_));
 sky130_fd_sc_hd__clkbuf_1 _16594_ (.A(_03032_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _16595_ (.A0(_06997_),
    .A1(\cpuregs.regs[18][26] ),
    .S(_03026_),
    .X(_03033_));
 sky130_fd_sc_hd__clkbuf_1 _16596_ (.A(_03033_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _16597_ (.A0(_06999_),
    .A1(\cpuregs.regs[18][27] ),
    .S(_03026_),
    .X(_03034_));
 sky130_fd_sc_hd__clkbuf_1 _16598_ (.A(_03034_),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _16599_ (.A0(_07001_),
    .A1(\cpuregs.regs[18][28] ),
    .S(_03026_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_1 _16600_ (.A(_03035_),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _16601_ (.A0(_07003_),
    .A1(\cpuregs.regs[18][29] ),
    .S(_03026_),
    .X(_03036_));
 sky130_fd_sc_hd__clkbuf_1 _16602_ (.A(_03036_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _16603_ (.A0(_07005_),
    .A1(\cpuregs.regs[18][30] ),
    .S(_03003_),
    .X(_03037_));
 sky130_fd_sc_hd__clkbuf_1 _16604_ (.A(_03037_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _16605_ (.A0(_07007_),
    .A1(\cpuregs.regs[18][31] ),
    .S(_03003_),
    .X(_03038_));
 sky130_fd_sc_hd__clkbuf_1 _16606_ (.A(_03038_),
    .X(_01581_));
 sky130_fd_sc_hd__nor3b_4 _16607_ (.A(_06750_),
    .B(\cpuregs.waddr[1] ),
    .C_N(\cpuregs.waddr[0] ),
    .Y(_03039_));
 sky130_fd_sc_hd__buf_6 _16608_ (.A(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__mux2_1 _16609_ (.A0(\cpuregs.regs[1][0] ),
    .A1(_06077_),
    .S(_03040_),
    .X(_03041_));
 sky130_fd_sc_hd__clkbuf_1 _16610_ (.A(_03041_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _16611_ (.A0(\cpuregs.regs[1][1] ),
    .A1(_06095_),
    .S(_03040_),
    .X(_03042_));
 sky130_fd_sc_hd__clkbuf_1 _16612_ (.A(_03042_),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _16613_ (.A0(\cpuregs.regs[1][2] ),
    .A1(_06104_),
    .S(_03040_),
    .X(_03043_));
 sky130_fd_sc_hd__clkbuf_1 _16614_ (.A(_03043_),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _16615_ (.A0(\cpuregs.regs[1][3] ),
    .A1(_06113_),
    .S(_03040_),
    .X(_03044_));
 sky130_fd_sc_hd__clkbuf_1 _16616_ (.A(_03044_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _16617_ (.A0(\cpuregs.regs[1][4] ),
    .A1(_06124_),
    .S(_03040_),
    .X(_03045_));
 sky130_fd_sc_hd__clkbuf_1 _16618_ (.A(_03045_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _16619_ (.A0(\cpuregs.regs[1][5] ),
    .A1(_06131_),
    .S(_03040_),
    .X(_03046_));
 sky130_fd_sc_hd__clkbuf_1 _16620_ (.A(_03046_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _16621_ (.A0(\cpuregs.regs[1][6] ),
    .A1(_06140_),
    .S(_03040_),
    .X(_03047_));
 sky130_fd_sc_hd__clkbuf_1 _16622_ (.A(_03047_),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _16623_ (.A0(\cpuregs.regs[1][7] ),
    .A1(_06149_),
    .S(_03040_),
    .X(_03048_));
 sky130_fd_sc_hd__clkbuf_1 _16624_ (.A(_03048_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _16625_ (.A0(\cpuregs.regs[1][8] ),
    .A1(_06156_),
    .S(_03040_),
    .X(_03049_));
 sky130_fd_sc_hd__clkbuf_1 _16626_ (.A(_03049_),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _16627_ (.A0(\cpuregs.regs[1][9] ),
    .A1(_06165_),
    .S(_03040_),
    .X(_03050_));
 sky130_fd_sc_hd__clkbuf_1 _16628_ (.A(_03050_),
    .X(_01591_));
 sky130_fd_sc_hd__clkbuf_8 _16629_ (.A(_03039_),
    .X(_03051_));
 sky130_fd_sc_hd__mux2_1 _16630_ (.A0(\cpuregs.regs[1][10] ),
    .A1(_06174_),
    .S(_03051_),
    .X(_03052_));
 sky130_fd_sc_hd__clkbuf_1 _16631_ (.A(_03052_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _16632_ (.A0(\cpuregs.regs[1][11] ),
    .A1(_06183_),
    .S(_03051_),
    .X(_03053_));
 sky130_fd_sc_hd__clkbuf_1 _16633_ (.A(_03053_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _16634_ (.A0(\cpuregs.regs[1][12] ),
    .A1(_06192_),
    .S(_03051_),
    .X(_03054_));
 sky130_fd_sc_hd__clkbuf_1 _16635_ (.A(_03054_),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _16636_ (.A0(\cpuregs.regs[1][13] ),
    .A1(_06200_),
    .S(_03051_),
    .X(_03055_));
 sky130_fd_sc_hd__clkbuf_1 _16637_ (.A(_03055_),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _16638_ (.A0(\cpuregs.regs[1][14] ),
    .A1(_06207_),
    .S(_03051_),
    .X(_03056_));
 sky130_fd_sc_hd__clkbuf_1 _16639_ (.A(_03056_),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _16640_ (.A0(\cpuregs.regs[1][15] ),
    .A1(_06215_),
    .S(_03051_),
    .X(_03057_));
 sky130_fd_sc_hd__clkbuf_1 _16641_ (.A(_03057_),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _16642_ (.A0(\cpuregs.regs[1][16] ),
    .A1(_06223_),
    .S(_03051_),
    .X(_03058_));
 sky130_fd_sc_hd__clkbuf_1 _16643_ (.A(_03058_),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _16644_ (.A0(\cpuregs.regs[1][17] ),
    .A1(_06231_),
    .S(_03051_),
    .X(_03059_));
 sky130_fd_sc_hd__clkbuf_1 _16645_ (.A(_03059_),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _16646_ (.A0(\cpuregs.regs[1][18] ),
    .A1(_06239_),
    .S(_03051_),
    .X(_03060_));
 sky130_fd_sc_hd__clkbuf_1 _16647_ (.A(_03060_),
    .X(_01600_));
 sky130_fd_sc_hd__mux2_1 _16648_ (.A0(\cpuregs.regs[1][19] ),
    .A1(_06247_),
    .S(_03051_),
    .X(_03061_));
 sky130_fd_sc_hd__clkbuf_1 _16649_ (.A(_03061_),
    .X(_01601_));
 sky130_fd_sc_hd__buf_6 _16650_ (.A(_03039_),
    .X(_03062_));
 sky130_fd_sc_hd__mux2_1 _16651_ (.A0(\cpuregs.regs[1][20] ),
    .A1(_06256_),
    .S(_03062_),
    .X(_03063_));
 sky130_fd_sc_hd__clkbuf_1 _16652_ (.A(_03063_),
    .X(_01602_));
 sky130_fd_sc_hd__mux2_1 _16653_ (.A0(\cpuregs.regs[1][21] ),
    .A1(_06265_),
    .S(_03062_),
    .X(_03064_));
 sky130_fd_sc_hd__clkbuf_1 _16654_ (.A(_03064_),
    .X(_01603_));
 sky130_fd_sc_hd__mux2_1 _16655_ (.A0(\cpuregs.regs[1][22] ),
    .A1(_06273_),
    .S(_03062_),
    .X(_03065_));
 sky130_fd_sc_hd__clkbuf_1 _16656_ (.A(_03065_),
    .X(_01604_));
 sky130_fd_sc_hd__mux2_1 _16657_ (.A0(\cpuregs.regs[1][23] ),
    .A1(_06280_),
    .S(_03062_),
    .X(_03066_));
 sky130_fd_sc_hd__clkbuf_1 _16658_ (.A(_03066_),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _16659_ (.A0(\cpuregs.regs[1][24] ),
    .A1(_06288_),
    .S(_03062_),
    .X(_03067_));
 sky130_fd_sc_hd__clkbuf_1 _16660_ (.A(_03067_),
    .X(_01606_));
 sky130_fd_sc_hd__mux2_1 _16661_ (.A0(\cpuregs.regs[1][25] ),
    .A1(_06296_),
    .S(_03062_),
    .X(_03068_));
 sky130_fd_sc_hd__clkbuf_1 _16662_ (.A(_03068_),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_1 _16663_ (.A0(\cpuregs.regs[1][26] ),
    .A1(_06303_),
    .S(_03062_),
    .X(_03069_));
 sky130_fd_sc_hd__clkbuf_1 _16664_ (.A(_03069_),
    .X(_01608_));
 sky130_fd_sc_hd__mux2_1 _16665_ (.A0(\cpuregs.regs[1][27] ),
    .A1(_06311_),
    .S(_03062_),
    .X(_03070_));
 sky130_fd_sc_hd__clkbuf_1 _16666_ (.A(_03070_),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _16667_ (.A0(\cpuregs.regs[1][28] ),
    .A1(_06319_),
    .S(_03062_),
    .X(_03071_));
 sky130_fd_sc_hd__clkbuf_1 _16668_ (.A(_03071_),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _16669_ (.A0(\cpuregs.regs[1][29] ),
    .A1(_06327_),
    .S(_03062_),
    .X(_03072_));
 sky130_fd_sc_hd__clkbuf_1 _16670_ (.A(_03072_),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _16671_ (.A0(\cpuregs.regs[1][30] ),
    .A1(_06335_),
    .S(_03039_),
    .X(_03073_));
 sky130_fd_sc_hd__clkbuf_1 _16672_ (.A(_03073_),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_1 _16673_ (.A0(\cpuregs.regs[1][31] ),
    .A1(_06342_),
    .S(_03039_),
    .X(_03074_));
 sky130_fd_sc_hd__clkbuf_1 _16674_ (.A(_03074_),
    .X(_01613_));
 sky130_fd_sc_hd__nand2_4 _16675_ (.A(_06346_),
    .B(_02894_),
    .Y(_03075_));
 sky130_fd_sc_hd__clkbuf_8 _16676_ (.A(_03075_),
    .X(_03076_));
 sky130_fd_sc_hd__mux2_1 _16677_ (.A0(_06941_),
    .A1(\cpuregs.regs[19][0] ),
    .S(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__clkbuf_1 _16678_ (.A(_03077_),
    .X(_01614_));
 sky130_fd_sc_hd__mux2_1 _16679_ (.A0(_06945_),
    .A1(\cpuregs.regs[19][1] ),
    .S(_03076_),
    .X(_03078_));
 sky130_fd_sc_hd__clkbuf_1 _16680_ (.A(_03078_),
    .X(_01615_));
 sky130_fd_sc_hd__mux2_1 _16681_ (.A0(_06947_),
    .A1(\cpuregs.regs[19][2] ),
    .S(_03076_),
    .X(_03079_));
 sky130_fd_sc_hd__clkbuf_1 _16682_ (.A(_03079_),
    .X(_01616_));
 sky130_fd_sc_hd__mux2_1 _16683_ (.A0(_06949_),
    .A1(\cpuregs.regs[19][3] ),
    .S(_03076_),
    .X(_03080_));
 sky130_fd_sc_hd__clkbuf_1 _16684_ (.A(_03080_),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _16685_ (.A0(_06951_),
    .A1(\cpuregs.regs[19][4] ),
    .S(_03076_),
    .X(_03081_));
 sky130_fd_sc_hd__clkbuf_1 _16686_ (.A(_03081_),
    .X(_01618_));
 sky130_fd_sc_hd__mux2_1 _16687_ (.A0(_06953_),
    .A1(\cpuregs.regs[19][5] ),
    .S(_03076_),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_1 _16688_ (.A(_03082_),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _16689_ (.A0(_06955_),
    .A1(\cpuregs.regs[19][6] ),
    .S(_03076_),
    .X(_03083_));
 sky130_fd_sc_hd__clkbuf_1 _16690_ (.A(_03083_),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _16691_ (.A0(_06957_),
    .A1(\cpuregs.regs[19][7] ),
    .S(_03076_),
    .X(_03084_));
 sky130_fd_sc_hd__clkbuf_1 _16692_ (.A(_03084_),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _16693_ (.A0(_06959_),
    .A1(\cpuregs.regs[19][8] ),
    .S(_03076_),
    .X(_03085_));
 sky130_fd_sc_hd__clkbuf_1 _16694_ (.A(_03085_),
    .X(_01622_));
 sky130_fd_sc_hd__mux2_1 _16695_ (.A0(_06961_),
    .A1(\cpuregs.regs[19][9] ),
    .S(_03076_),
    .X(_03086_));
 sky130_fd_sc_hd__clkbuf_1 _16696_ (.A(_03086_),
    .X(_01623_));
 sky130_fd_sc_hd__clkbuf_8 _16697_ (.A(_03075_),
    .X(_03087_));
 sky130_fd_sc_hd__mux2_1 _16698_ (.A0(_06963_),
    .A1(\cpuregs.regs[19][10] ),
    .S(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__clkbuf_1 _16699_ (.A(_03088_),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _16700_ (.A0(_06966_),
    .A1(\cpuregs.regs[19][11] ),
    .S(_03087_),
    .X(_03089_));
 sky130_fd_sc_hd__clkbuf_1 _16701_ (.A(_03089_),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _16702_ (.A0(_06968_),
    .A1(\cpuregs.regs[19][12] ),
    .S(_03087_),
    .X(_03090_));
 sky130_fd_sc_hd__clkbuf_1 _16703_ (.A(_03090_),
    .X(_01626_));
 sky130_fd_sc_hd__mux2_1 _16704_ (.A0(_06970_),
    .A1(\cpuregs.regs[19][13] ),
    .S(_03087_),
    .X(_03091_));
 sky130_fd_sc_hd__clkbuf_1 _16705_ (.A(_03091_),
    .X(_01627_));
 sky130_fd_sc_hd__mux2_1 _16706_ (.A0(_06972_),
    .A1(\cpuregs.regs[19][14] ),
    .S(_03087_),
    .X(_03092_));
 sky130_fd_sc_hd__clkbuf_1 _16707_ (.A(_03092_),
    .X(_01628_));
 sky130_fd_sc_hd__mux2_1 _16708_ (.A0(_06974_),
    .A1(\cpuregs.regs[19][15] ),
    .S(_03087_),
    .X(_03093_));
 sky130_fd_sc_hd__clkbuf_1 _16709_ (.A(_03093_),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _16710_ (.A0(_06976_),
    .A1(\cpuregs.regs[19][16] ),
    .S(_03087_),
    .X(_03094_));
 sky130_fd_sc_hd__clkbuf_1 _16711_ (.A(_03094_),
    .X(_01630_));
 sky130_fd_sc_hd__mux2_1 _16712_ (.A0(_06978_),
    .A1(\cpuregs.regs[19][17] ),
    .S(_03087_),
    .X(_03095_));
 sky130_fd_sc_hd__clkbuf_1 _16713_ (.A(_03095_),
    .X(_01631_));
 sky130_fd_sc_hd__mux2_1 _16714_ (.A0(_06980_),
    .A1(\cpuregs.regs[19][18] ),
    .S(_03087_),
    .X(_03096_));
 sky130_fd_sc_hd__clkbuf_1 _16715_ (.A(_03096_),
    .X(_01632_));
 sky130_fd_sc_hd__mux2_1 _16716_ (.A0(_06982_),
    .A1(\cpuregs.regs[19][19] ),
    .S(_03087_),
    .X(_03097_));
 sky130_fd_sc_hd__clkbuf_1 _16717_ (.A(_03097_),
    .X(_01633_));
 sky130_fd_sc_hd__buf_6 _16718_ (.A(_03075_),
    .X(_03098_));
 sky130_fd_sc_hd__mux2_1 _16719_ (.A0(_06984_),
    .A1(\cpuregs.regs[19][20] ),
    .S(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__clkbuf_1 _16720_ (.A(_03099_),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_1 _16721_ (.A0(_06987_),
    .A1(\cpuregs.regs[19][21] ),
    .S(_03098_),
    .X(_03100_));
 sky130_fd_sc_hd__clkbuf_1 _16722_ (.A(_03100_),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _16723_ (.A0(_06989_),
    .A1(\cpuregs.regs[19][22] ),
    .S(_03098_),
    .X(_03101_));
 sky130_fd_sc_hd__clkbuf_1 _16724_ (.A(_03101_),
    .X(_01636_));
 sky130_fd_sc_hd__mux2_1 _16725_ (.A0(_06991_),
    .A1(\cpuregs.regs[19][23] ),
    .S(_03098_),
    .X(_03102_));
 sky130_fd_sc_hd__clkbuf_1 _16726_ (.A(_03102_),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _16727_ (.A0(_06993_),
    .A1(\cpuregs.regs[19][24] ),
    .S(_03098_),
    .X(_03103_));
 sky130_fd_sc_hd__clkbuf_1 _16728_ (.A(_03103_),
    .X(_01638_));
 sky130_fd_sc_hd__mux2_1 _16729_ (.A0(_06995_),
    .A1(\cpuregs.regs[19][25] ),
    .S(_03098_),
    .X(_03104_));
 sky130_fd_sc_hd__clkbuf_1 _16730_ (.A(_03104_),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_1 _16731_ (.A0(_06997_),
    .A1(\cpuregs.regs[19][26] ),
    .S(_03098_),
    .X(_03105_));
 sky130_fd_sc_hd__clkbuf_1 _16732_ (.A(_03105_),
    .X(_01640_));
 sky130_fd_sc_hd__mux2_1 _16733_ (.A0(_06999_),
    .A1(\cpuregs.regs[19][27] ),
    .S(_03098_),
    .X(_03106_));
 sky130_fd_sc_hd__clkbuf_1 _16734_ (.A(_03106_),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _16735_ (.A0(_07001_),
    .A1(\cpuregs.regs[19][28] ),
    .S(_03098_),
    .X(_03107_));
 sky130_fd_sc_hd__clkbuf_1 _16736_ (.A(_03107_),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _16737_ (.A0(_07003_),
    .A1(\cpuregs.regs[19][29] ),
    .S(_03098_),
    .X(_03108_));
 sky130_fd_sc_hd__clkbuf_1 _16738_ (.A(_03108_),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _16739_ (.A0(_07005_),
    .A1(\cpuregs.regs[19][30] ),
    .S(_03075_),
    .X(_03109_));
 sky130_fd_sc_hd__clkbuf_1 _16740_ (.A(_03109_),
    .X(_01644_));
 sky130_fd_sc_hd__mux2_1 _16741_ (.A0(_07007_),
    .A1(\cpuregs.regs[19][31] ),
    .S(_03075_),
    .X(_03110_));
 sky130_fd_sc_hd__clkbuf_1 _16742_ (.A(_03110_),
    .X(_01645_));
 sky130_fd_sc_hd__o22a_1 _16743_ (.A1(\reg_sh[0] ),
    .A2(_03314_),
    .B1(_01929_),
    .B2(_03638_),
    .X(_03111_));
 sky130_fd_sc_hd__a21bo_1 _16744_ (.A1(\reg_sh[0] ),
    .A2(_07274_),
    .B1_N(_03111_),
    .X(_01646_));
 sky130_fd_sc_hd__nor2_1 _16745_ (.A(_03680_),
    .B(_01955_),
    .Y(_03112_));
 sky130_fd_sc_hd__o211a_1 _16746_ (.A1(\reg_sh[0] ),
    .A2(_03399_),
    .B1(_04046_),
    .C1(\reg_sh[1] ),
    .X(_03113_));
 sky130_fd_sc_hd__or3_1 _16747_ (.A(_03316_),
    .B(_03112_),
    .C(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__clkbuf_1 _16748_ (.A(_03114_),
    .X(_01647_));
 sky130_fd_sc_hd__nand2_2 _16749_ (.A(_06422_),
    .B(_06823_),
    .Y(_03115_));
 sky130_fd_sc_hd__buf_6 _16750_ (.A(_03115_),
    .X(_03116_));
 sky130_fd_sc_hd__mux2_1 _16751_ (.A0(_06531_),
    .A1(\cpuregs.regs[13][0] ),
    .S(_03116_),
    .X(_03117_));
 sky130_fd_sc_hd__clkbuf_1 _16752_ (.A(_03117_),
    .X(_01648_));
 sky130_fd_sc_hd__mux2_1 _16753_ (.A0(_06536_),
    .A1(\cpuregs.regs[13][1] ),
    .S(_03116_),
    .X(_03118_));
 sky130_fd_sc_hd__clkbuf_1 _16754_ (.A(_03118_),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _16755_ (.A0(_06538_),
    .A1(\cpuregs.regs[13][2] ),
    .S(_03116_),
    .X(_03119_));
 sky130_fd_sc_hd__clkbuf_1 _16756_ (.A(_03119_),
    .X(_01650_));
 sky130_fd_sc_hd__mux2_1 _16757_ (.A0(_06540_),
    .A1(\cpuregs.regs[13][3] ),
    .S(_03116_),
    .X(_03120_));
 sky130_fd_sc_hd__clkbuf_1 _16758_ (.A(_03120_),
    .X(_01651_));
 sky130_fd_sc_hd__mux2_1 _16759_ (.A0(_06542_),
    .A1(\cpuregs.regs[13][4] ),
    .S(_03116_),
    .X(_03121_));
 sky130_fd_sc_hd__clkbuf_1 _16760_ (.A(_03121_),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _16761_ (.A0(_06544_),
    .A1(\cpuregs.regs[13][5] ),
    .S(_03116_),
    .X(_03122_));
 sky130_fd_sc_hd__clkbuf_1 _16762_ (.A(_03122_),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _16763_ (.A0(_06546_),
    .A1(\cpuregs.regs[13][6] ),
    .S(_03116_),
    .X(_03123_));
 sky130_fd_sc_hd__clkbuf_1 _16764_ (.A(_03123_),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_1 _16765_ (.A0(_06548_),
    .A1(\cpuregs.regs[13][7] ),
    .S(_03116_),
    .X(_03124_));
 sky130_fd_sc_hd__clkbuf_1 _16766_ (.A(_03124_),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _16767_ (.A0(_06550_),
    .A1(\cpuregs.regs[13][8] ),
    .S(_03116_),
    .X(_03125_));
 sky130_fd_sc_hd__clkbuf_1 _16768_ (.A(_03125_),
    .X(_01656_));
 sky130_fd_sc_hd__mux2_1 _16769_ (.A0(_06552_),
    .A1(\cpuregs.regs[13][9] ),
    .S(_03116_),
    .X(_03126_));
 sky130_fd_sc_hd__clkbuf_1 _16770_ (.A(_03126_),
    .X(_01657_));
 sky130_fd_sc_hd__buf_6 _16771_ (.A(_03115_),
    .X(_03127_));
 sky130_fd_sc_hd__mux2_1 _16772_ (.A0(_06554_),
    .A1(\cpuregs.regs[13][10] ),
    .S(_03127_),
    .X(_03128_));
 sky130_fd_sc_hd__clkbuf_1 _16773_ (.A(_03128_),
    .X(_01658_));
 sky130_fd_sc_hd__mux2_1 _16774_ (.A0(_06557_),
    .A1(\cpuregs.regs[13][11] ),
    .S(_03127_),
    .X(_03129_));
 sky130_fd_sc_hd__clkbuf_1 _16775_ (.A(_03129_),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _16776_ (.A0(_06559_),
    .A1(\cpuregs.regs[13][12] ),
    .S(_03127_),
    .X(_03130_));
 sky130_fd_sc_hd__clkbuf_1 _16777_ (.A(_03130_),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_1 _16778_ (.A0(_06561_),
    .A1(\cpuregs.regs[13][13] ),
    .S(_03127_),
    .X(_03131_));
 sky130_fd_sc_hd__clkbuf_1 _16779_ (.A(_03131_),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _16780_ (.A0(_06563_),
    .A1(\cpuregs.regs[13][14] ),
    .S(_03127_),
    .X(_03132_));
 sky130_fd_sc_hd__clkbuf_1 _16781_ (.A(_03132_),
    .X(_01662_));
 sky130_fd_sc_hd__mux2_1 _16782_ (.A0(_06565_),
    .A1(\cpuregs.regs[13][15] ),
    .S(_03127_),
    .X(_03133_));
 sky130_fd_sc_hd__clkbuf_1 _16783_ (.A(_03133_),
    .X(_01663_));
 sky130_fd_sc_hd__mux2_1 _16784_ (.A0(_06567_),
    .A1(\cpuregs.regs[13][16] ),
    .S(_03127_),
    .X(_03134_));
 sky130_fd_sc_hd__clkbuf_1 _16785_ (.A(_03134_),
    .X(_01664_));
 sky130_fd_sc_hd__mux2_1 _16786_ (.A0(_06569_),
    .A1(\cpuregs.regs[13][17] ),
    .S(_03127_),
    .X(_03135_));
 sky130_fd_sc_hd__clkbuf_1 _16787_ (.A(_03135_),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _16788_ (.A0(_06571_),
    .A1(\cpuregs.regs[13][18] ),
    .S(_03127_),
    .X(_03136_));
 sky130_fd_sc_hd__clkbuf_1 _16789_ (.A(_03136_),
    .X(_01666_));
 sky130_fd_sc_hd__mux2_1 _16790_ (.A0(_06573_),
    .A1(\cpuregs.regs[13][19] ),
    .S(_03127_),
    .X(_03137_));
 sky130_fd_sc_hd__clkbuf_1 _16791_ (.A(_03137_),
    .X(_01667_));
 sky130_fd_sc_hd__buf_4 _16792_ (.A(_03115_),
    .X(_03138_));
 sky130_fd_sc_hd__mux2_1 _16793_ (.A0(_06575_),
    .A1(\cpuregs.regs[13][20] ),
    .S(_03138_),
    .X(_03139_));
 sky130_fd_sc_hd__clkbuf_1 _16794_ (.A(_03139_),
    .X(_01668_));
 sky130_fd_sc_hd__mux2_1 _16795_ (.A0(_06578_),
    .A1(\cpuregs.regs[13][21] ),
    .S(_03138_),
    .X(_03140_));
 sky130_fd_sc_hd__clkbuf_1 _16796_ (.A(_03140_),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _16797_ (.A0(_06580_),
    .A1(\cpuregs.regs[13][22] ),
    .S(_03138_),
    .X(_03141_));
 sky130_fd_sc_hd__clkbuf_1 _16798_ (.A(_03141_),
    .X(_01670_));
 sky130_fd_sc_hd__mux2_1 _16799_ (.A0(_06582_),
    .A1(\cpuregs.regs[13][23] ),
    .S(_03138_),
    .X(_03142_));
 sky130_fd_sc_hd__clkbuf_1 _16800_ (.A(_03142_),
    .X(_01671_));
 sky130_fd_sc_hd__mux2_1 _16801_ (.A0(_06584_),
    .A1(\cpuregs.regs[13][24] ),
    .S(_03138_),
    .X(_03143_));
 sky130_fd_sc_hd__clkbuf_1 _16802_ (.A(_03143_),
    .X(_01672_));
 sky130_fd_sc_hd__mux2_1 _16803_ (.A0(_06586_),
    .A1(\cpuregs.regs[13][25] ),
    .S(_03138_),
    .X(_03144_));
 sky130_fd_sc_hd__clkbuf_1 _16804_ (.A(_03144_),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _16805_ (.A0(_06588_),
    .A1(\cpuregs.regs[13][26] ),
    .S(_03138_),
    .X(_03145_));
 sky130_fd_sc_hd__clkbuf_1 _16806_ (.A(_03145_),
    .X(_01674_));
 sky130_fd_sc_hd__mux2_1 _16807_ (.A0(_06590_),
    .A1(\cpuregs.regs[13][27] ),
    .S(_03138_),
    .X(_03146_));
 sky130_fd_sc_hd__clkbuf_1 _16808_ (.A(_03146_),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_1 _16809_ (.A0(_06592_),
    .A1(\cpuregs.regs[13][28] ),
    .S(_03138_),
    .X(_03147_));
 sky130_fd_sc_hd__clkbuf_1 _16810_ (.A(_03147_),
    .X(_01676_));
 sky130_fd_sc_hd__mux2_1 _16811_ (.A0(_06594_),
    .A1(\cpuregs.regs[13][29] ),
    .S(_03138_),
    .X(_03148_));
 sky130_fd_sc_hd__clkbuf_1 _16812_ (.A(_03148_),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _16813_ (.A0(_06596_),
    .A1(\cpuregs.regs[13][30] ),
    .S(_03115_),
    .X(_03149_));
 sky130_fd_sc_hd__clkbuf_1 _16814_ (.A(_03149_),
    .X(_01678_));
 sky130_fd_sc_hd__mux2_1 _16815_ (.A0(_06598_),
    .A1(\cpuregs.regs[13][31] ),
    .S(_03115_),
    .X(_03150_));
 sky130_fd_sc_hd__clkbuf_1 _16816_ (.A(_03150_),
    .X(_01679_));
 sky130_fd_sc_hd__nand2_4 _16817_ (.A(_06080_),
    .B(_06823_),
    .Y(_03151_));
 sky130_fd_sc_hd__buf_6 _16818_ (.A(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__mux2_1 _16819_ (.A0(_06531_),
    .A1(\cpuregs.regs[14][0] ),
    .S(_03152_),
    .X(_03153_));
 sky130_fd_sc_hd__clkbuf_1 _16820_ (.A(_03153_),
    .X(_01680_));
 sky130_fd_sc_hd__mux2_1 _16821_ (.A0(_06536_),
    .A1(\cpuregs.regs[14][1] ),
    .S(_03152_),
    .X(_03154_));
 sky130_fd_sc_hd__clkbuf_1 _16822_ (.A(_03154_),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _16823_ (.A0(_06538_),
    .A1(\cpuregs.regs[14][2] ),
    .S(_03152_),
    .X(_03155_));
 sky130_fd_sc_hd__clkbuf_1 _16824_ (.A(_03155_),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_1 _16825_ (.A0(_06540_),
    .A1(\cpuregs.regs[14][3] ),
    .S(_03152_),
    .X(_03156_));
 sky130_fd_sc_hd__clkbuf_1 _16826_ (.A(_03156_),
    .X(_01683_));
 sky130_fd_sc_hd__mux2_1 _16827_ (.A0(_06542_),
    .A1(\cpuregs.regs[14][4] ),
    .S(_03152_),
    .X(_03157_));
 sky130_fd_sc_hd__clkbuf_1 _16828_ (.A(_03157_),
    .X(_01684_));
 sky130_fd_sc_hd__mux2_1 _16829_ (.A0(_06544_),
    .A1(\cpuregs.regs[14][5] ),
    .S(_03152_),
    .X(_03158_));
 sky130_fd_sc_hd__clkbuf_1 _16830_ (.A(_03158_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _16831_ (.A0(_06546_),
    .A1(\cpuregs.regs[14][6] ),
    .S(_03152_),
    .X(_03159_));
 sky130_fd_sc_hd__clkbuf_1 _16832_ (.A(_03159_),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_1 _16833_ (.A0(_06548_),
    .A1(\cpuregs.regs[14][7] ),
    .S(_03152_),
    .X(_03160_));
 sky130_fd_sc_hd__clkbuf_1 _16834_ (.A(_03160_),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_1 _16835_ (.A0(_06550_),
    .A1(\cpuregs.regs[14][8] ),
    .S(_03152_),
    .X(_03161_));
 sky130_fd_sc_hd__clkbuf_1 _16836_ (.A(_03161_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _16837_ (.A0(_06552_),
    .A1(\cpuregs.regs[14][9] ),
    .S(_03152_),
    .X(_03162_));
 sky130_fd_sc_hd__clkbuf_1 _16838_ (.A(_03162_),
    .X(_01689_));
 sky130_fd_sc_hd__buf_6 _16839_ (.A(_03151_),
    .X(_03163_));
 sky130_fd_sc_hd__mux2_1 _16840_ (.A0(_06554_),
    .A1(\cpuregs.regs[14][10] ),
    .S(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__clkbuf_1 _16841_ (.A(_03164_),
    .X(_01690_));
 sky130_fd_sc_hd__mux2_1 _16842_ (.A0(_06557_),
    .A1(\cpuregs.regs[14][11] ),
    .S(_03163_),
    .X(_03165_));
 sky130_fd_sc_hd__clkbuf_1 _16843_ (.A(_03165_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _16844_ (.A0(_06559_),
    .A1(\cpuregs.regs[14][12] ),
    .S(_03163_),
    .X(_03166_));
 sky130_fd_sc_hd__clkbuf_1 _16845_ (.A(_03166_),
    .X(_01692_));
 sky130_fd_sc_hd__mux2_1 _16846_ (.A0(_06561_),
    .A1(\cpuregs.regs[14][13] ),
    .S(_03163_),
    .X(_03167_));
 sky130_fd_sc_hd__clkbuf_1 _16847_ (.A(_03167_),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _16848_ (.A0(_06563_),
    .A1(\cpuregs.regs[14][14] ),
    .S(_03163_),
    .X(_03168_));
 sky130_fd_sc_hd__clkbuf_1 _16849_ (.A(_03168_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _16850_ (.A0(_06565_),
    .A1(\cpuregs.regs[14][15] ),
    .S(_03163_),
    .X(_03169_));
 sky130_fd_sc_hd__clkbuf_1 _16851_ (.A(_03169_),
    .X(_01695_));
 sky130_fd_sc_hd__mux2_1 _16852_ (.A0(_06567_),
    .A1(\cpuregs.regs[14][16] ),
    .S(_03163_),
    .X(_03170_));
 sky130_fd_sc_hd__clkbuf_1 _16853_ (.A(_03170_),
    .X(_01696_));
 sky130_fd_sc_hd__mux2_1 _16854_ (.A0(_06569_),
    .A1(\cpuregs.regs[14][17] ),
    .S(_03163_),
    .X(_03171_));
 sky130_fd_sc_hd__clkbuf_1 _16855_ (.A(_03171_),
    .X(_01697_));
 sky130_fd_sc_hd__mux2_1 _16856_ (.A0(_06571_),
    .A1(\cpuregs.regs[14][18] ),
    .S(_03163_),
    .X(_03172_));
 sky130_fd_sc_hd__clkbuf_1 _16857_ (.A(_03172_),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_1 _16858_ (.A0(_06573_),
    .A1(\cpuregs.regs[14][19] ),
    .S(_03163_),
    .X(_03173_));
 sky130_fd_sc_hd__clkbuf_1 _16859_ (.A(_03173_),
    .X(_01699_));
 sky130_fd_sc_hd__clkbuf_8 _16860_ (.A(_03151_),
    .X(_03174_));
 sky130_fd_sc_hd__mux2_1 _16861_ (.A0(_06575_),
    .A1(\cpuregs.regs[14][20] ),
    .S(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__clkbuf_1 _16862_ (.A(_03175_),
    .X(_01700_));
 sky130_fd_sc_hd__mux2_1 _16863_ (.A0(_06578_),
    .A1(\cpuregs.regs[14][21] ),
    .S(_03174_),
    .X(_03176_));
 sky130_fd_sc_hd__clkbuf_1 _16864_ (.A(_03176_),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_1 _16865_ (.A0(_06580_),
    .A1(\cpuregs.regs[14][22] ),
    .S(_03174_),
    .X(_03177_));
 sky130_fd_sc_hd__clkbuf_1 _16866_ (.A(_03177_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _16867_ (.A0(_06582_),
    .A1(\cpuregs.regs[14][23] ),
    .S(_03174_),
    .X(_03178_));
 sky130_fd_sc_hd__clkbuf_1 _16868_ (.A(_03178_),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _16869_ (.A0(_06584_),
    .A1(\cpuregs.regs[14][24] ),
    .S(_03174_),
    .X(_03179_));
 sky130_fd_sc_hd__clkbuf_1 _16870_ (.A(_03179_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _16871_ (.A0(_06586_),
    .A1(\cpuregs.regs[14][25] ),
    .S(_03174_),
    .X(_03180_));
 sky130_fd_sc_hd__clkbuf_1 _16872_ (.A(_03180_),
    .X(_01705_));
 sky130_fd_sc_hd__mux2_1 _16873_ (.A0(_06588_),
    .A1(\cpuregs.regs[14][26] ),
    .S(_03174_),
    .X(_03181_));
 sky130_fd_sc_hd__clkbuf_1 _16874_ (.A(_03181_),
    .X(_01706_));
 sky130_fd_sc_hd__mux2_1 _16875_ (.A0(_06590_),
    .A1(\cpuregs.regs[14][27] ),
    .S(_03174_),
    .X(_03182_));
 sky130_fd_sc_hd__clkbuf_1 _16876_ (.A(_03182_),
    .X(_01707_));
 sky130_fd_sc_hd__mux2_1 _16877_ (.A0(_06592_),
    .A1(\cpuregs.regs[14][28] ),
    .S(_03174_),
    .X(_03183_));
 sky130_fd_sc_hd__clkbuf_1 _16878_ (.A(_03183_),
    .X(_01708_));
 sky130_fd_sc_hd__mux2_1 _16879_ (.A0(_06594_),
    .A1(\cpuregs.regs[14][29] ),
    .S(_03174_),
    .X(_03184_));
 sky130_fd_sc_hd__clkbuf_1 _16880_ (.A(_03184_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _16881_ (.A0(_06596_),
    .A1(\cpuregs.regs[14][30] ),
    .S(_03151_),
    .X(_03185_));
 sky130_fd_sc_hd__clkbuf_1 _16882_ (.A(_03185_),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _16883_ (.A0(_06598_),
    .A1(\cpuregs.regs[14][31] ),
    .S(_03151_),
    .X(_03186_));
 sky130_fd_sc_hd__clkbuf_1 _16884_ (.A(_03186_),
    .X(_01711_));
 sky130_fd_sc_hd__dfxtp_1 _16885_ (.CLK(clknet_leaf_41_clk),
    .D(_00081_),
    .Q(\mem_wordsize[0] ));
 sky130_fd_sc_hd__dfxtp_2 _16886_ (.CLK(clknet_leaf_39_clk),
    .D(_00082_),
    .Q(\mem_wordsize[1] ));
 sky130_fd_sc_hd__dfxtp_2 _16887_ (.CLK(clknet_leaf_43_clk),
    .D(_00083_),
    .Q(\mem_wordsize[2] ));
 sky130_fd_sc_hd__dfxtp_1 _16888_ (.CLK(clknet_leaf_33_clk),
    .D(_00058_),
    .Q(\mem_rdata_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _16889_ (.CLK(clknet_leaf_33_clk),
    .D(_00059_),
    .Q(\mem_rdata_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _16890_ (.CLK(clknet_leaf_33_clk),
    .D(_00060_),
    .Q(\mem_rdata_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _16891_ (.CLK(clknet_leaf_31_clk),
    .D(_00036_),
    .Q(\mem_rdata_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _16892_ (.CLK(clknet_leaf_31_clk),
    .D(_00037_),
    .Q(\mem_rdata_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _16893_ (.CLK(clknet_leaf_35_clk),
    .D(_00038_),
    .Q(\mem_rdata_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _16894_ (.CLK(clknet_leaf_35_clk),
    .D(_00039_),
    .Q(\mem_rdata_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _16895_ (.CLK(clknet_leaf_34_clk),
    .D(_00040_),
    .Q(\mem_rdata_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _16896_ (.CLK(clknet_leaf_30_clk),
    .D(_00041_),
    .Q(\mem_rdata_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _16897_ (.CLK(clknet_leaf_30_clk),
    .D(_00042_),
    .Q(\mem_rdata_q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _16898_ (.CLK(clknet_leaf_29_clk),
    .D(_00043_),
    .Q(\mem_rdata_q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _16899_ (.CLK(clknet_leaf_30_clk),
    .D(_00044_),
    .Q(\mem_rdata_q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _16900_ (.CLK(clknet_leaf_31_clk),
    .D(_00045_),
    .Q(\mem_rdata_q[19] ));
 sky130_fd_sc_hd__dfxtp_2 _16901_ (.CLK(clknet_leaf_33_clk),
    .D(_00046_),
    .Q(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__dfxtp_2 _16902_ (.CLK(clknet_leaf_33_clk),
    .D(_00047_),
    .Q(\mem_rdata_q[21] ));
 sky130_fd_sc_hd__dfxtp_2 _16903_ (.CLK(clknet_leaf_33_clk),
    .D(_00048_),
    .Q(\mem_rdata_q[22] ));
 sky130_fd_sc_hd__dfxtp_2 _16904_ (.CLK(clknet_leaf_33_clk),
    .D(_00049_),
    .Q(\mem_rdata_q[23] ));
 sky130_fd_sc_hd__dfxtp_2 _16905_ (.CLK(clknet_leaf_34_clk),
    .D(_00050_),
    .Q(\mem_rdata_q[24] ));
 sky130_fd_sc_hd__dfxtp_2 _16906_ (.CLK(clknet_leaf_35_clk),
    .D(_00051_),
    .Q(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__dfxtp_4 _16907_ (.CLK(clknet_leaf_7_clk),
    .D(_00052_),
    .Q(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__dfxtp_4 _16908_ (.CLK(clknet_leaf_7_clk),
    .D(_00053_),
    .Q(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__dfxtp_2 _16909_ (.CLK(clknet_leaf_6_clk),
    .D(_00054_),
    .Q(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__dfxtp_2 _16910_ (.CLK(clknet_leaf_35_clk),
    .D(_00055_),
    .Q(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__dfxtp_2 _16911_ (.CLK(clknet_leaf_34_clk),
    .D(_00056_),
    .Q(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__dfxtp_2 _16912_ (.CLK(clknet_leaf_34_clk),
    .D(_00057_),
    .Q(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _16913_ (.CLK(clknet_leaf_40_clk),
    .D(_00094_),
    .Q(last_mem_valid));
 sky130_fd_sc_hd__dfxtp_1 _16914_ (.CLK(clknet_leaf_17_clk),
    .D(_00095_),
    .Q(\cpuregs.regs[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16915_ (.CLK(clknet_leaf_190_clk),
    .D(_00096_),
    .Q(\cpuregs.regs[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16916_ (.CLK(clknet_leaf_15_clk),
    .D(_00097_),
    .Q(\cpuregs.regs[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16917_ (.CLK(clknet_leaf_10_clk),
    .D(_00098_),
    .Q(\cpuregs.regs[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16918_ (.CLK(clknet_leaf_187_clk),
    .D(_00099_),
    .Q(\cpuregs.regs[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16919_ (.CLK(clknet_leaf_18_clk),
    .D(_00100_),
    .Q(\cpuregs.regs[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16920_ (.CLK(clknet_leaf_180_clk),
    .D(_00101_),
    .Q(\cpuregs.regs[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16921_ (.CLK(clknet_leaf_172_clk),
    .D(_00102_),
    .Q(\cpuregs.regs[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16922_ (.CLK(clknet_leaf_183_clk),
    .D(_00103_),
    .Q(\cpuregs.regs[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16923_ (.CLK(clknet_leaf_183_clk),
    .D(_00104_),
    .Q(\cpuregs.regs[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16924_ (.CLK(clknet_leaf_130_clk),
    .D(_00105_),
    .Q(\cpuregs.regs[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16925_ (.CLK(clknet_leaf_115_clk),
    .D(_00106_),
    .Q(\cpuregs.regs[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16926_ (.CLK(clknet_leaf_149_clk),
    .D(_00107_),
    .Q(\cpuregs.regs[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16927_ (.CLK(clknet_leaf_138_clk),
    .D(_00108_),
    .Q(\cpuregs.regs[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16928_ (.CLK(clknet_leaf_145_clk),
    .D(_00109_),
    .Q(\cpuregs.regs[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16929_ (.CLK(clknet_leaf_130_clk),
    .D(_00110_),
    .Q(\cpuregs.regs[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16930_ (.CLK(clknet_leaf_142_clk),
    .D(_00111_),
    .Q(\cpuregs.regs[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _16931_ (.CLK(clknet_leaf_140_clk),
    .D(_00112_),
    .Q(\cpuregs.regs[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _16932_ (.CLK(clknet_leaf_153_clk),
    .D(_00113_),
    .Q(\cpuregs.regs[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _16933_ (.CLK(clknet_leaf_179_clk),
    .D(_00114_),
    .Q(\cpuregs.regs[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _16934_ (.CLK(clknet_leaf_101_clk),
    .D(_00115_),
    .Q(\cpuregs.regs[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _16935_ (.CLK(clknet_leaf_101_clk),
    .D(_00116_),
    .Q(\cpuregs.regs[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _16936_ (.CLK(clknet_leaf_120_clk),
    .D(_00117_),
    .Q(\cpuregs.regs[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _16937_ (.CLK(clknet_leaf_164_clk),
    .D(_00118_),
    .Q(\cpuregs.regs[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _16938_ (.CLK(clknet_leaf_161_clk),
    .D(_00119_),
    .Q(\cpuregs.regs[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _16939_ (.CLK(clknet_leaf_110_clk),
    .D(_00120_),
    .Q(\cpuregs.regs[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _16940_ (.CLK(clknet_leaf_166_clk),
    .D(_00121_),
    .Q(\cpuregs.regs[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _16941_ (.CLK(clknet_leaf_105_clk),
    .D(_00122_),
    .Q(\cpuregs.regs[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _16942_ (.CLK(clknet_leaf_119_clk),
    .D(_00123_),
    .Q(\cpuregs.regs[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _16943_ (.CLK(clknet_leaf_117_clk),
    .D(_00124_),
    .Q(\cpuregs.regs[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _16944_ (.CLK(clknet_leaf_163_clk),
    .D(_00125_),
    .Q(\cpuregs.regs[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _16945_ (.CLK(clknet_leaf_169_clk),
    .D(_00126_),
    .Q(\cpuregs.regs[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _16946_ (.CLK(clknet_leaf_53_clk),
    .D(_00074_),
    .Q(\cpu_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _16947_ (.CLK(clknet_leaf_61_clk),
    .D(_00075_),
    .Q(\cpu_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _16948_ (.CLK(clknet_leaf_53_clk),
    .D(_00076_),
    .Q(\cpu_state[2] ));
 sky130_fd_sc_hd__dfxtp_4 _16949_ (.CLK(clknet_leaf_53_clk),
    .D(_00077_),
    .Q(\cpu_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _16950_ (.CLK(clknet_leaf_53_clk),
    .D(_00078_),
    .Q(\cpu_state[4] ));
 sky130_fd_sc_hd__dfxtp_2 _16951_ (.CLK(clknet_leaf_53_clk),
    .D(_00079_),
    .Q(\cpu_state[5] ));
 sky130_fd_sc_hd__dfxtp_4 _16952_ (.CLK(clknet_leaf_53_clk),
    .D(_00080_),
    .Q(\cpu_state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _16953_ (.CLK(clknet_leaf_17_clk),
    .D(_00127_),
    .Q(\cpuregs.regs[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16954_ (.CLK(clknet_leaf_190_clk),
    .D(_00128_),
    .Q(\cpuregs.regs[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16955_ (.CLK(clknet_leaf_10_clk),
    .D(_00129_),
    .Q(\cpuregs.regs[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16956_ (.CLK(clknet_leaf_10_clk),
    .D(_00130_),
    .Q(\cpuregs.regs[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16957_ (.CLK(clknet_leaf_187_clk),
    .D(_00131_),
    .Q(\cpuregs.regs[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16958_ (.CLK(clknet_leaf_18_clk),
    .D(_00132_),
    .Q(\cpuregs.regs[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16959_ (.CLK(clknet_leaf_180_clk),
    .D(_00133_),
    .Q(\cpuregs.regs[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16960_ (.CLK(clknet_leaf_172_clk),
    .D(_00134_),
    .Q(\cpuregs.regs[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16961_ (.CLK(clknet_leaf_183_clk),
    .D(_00135_),
    .Q(\cpuregs.regs[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16962_ (.CLK(clknet_leaf_182_clk),
    .D(_00136_),
    .Q(\cpuregs.regs[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16963_ (.CLK(clknet_leaf_130_clk),
    .D(_00137_),
    .Q(\cpuregs.regs[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16964_ (.CLK(clknet_leaf_115_clk),
    .D(_00138_),
    .Q(\cpuregs.regs[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16965_ (.CLK(clknet_leaf_149_clk),
    .D(_00139_),
    .Q(\cpuregs.regs[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16966_ (.CLK(clknet_leaf_138_clk),
    .D(_00140_),
    .Q(\cpuregs.regs[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16967_ (.CLK(clknet_leaf_145_clk),
    .D(_00141_),
    .Q(\cpuregs.regs[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16968_ (.CLK(clknet_leaf_129_clk),
    .D(_00142_),
    .Q(\cpuregs.regs[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16969_ (.CLK(clknet_leaf_142_clk),
    .D(_00143_),
    .Q(\cpuregs.regs[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _16970_ (.CLK(clknet_leaf_140_clk),
    .D(_00144_),
    .Q(\cpuregs.regs[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _16971_ (.CLK(clknet_leaf_153_clk),
    .D(_00145_),
    .Q(\cpuregs.regs[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _16972_ (.CLK(clknet_leaf_179_clk),
    .D(_00146_),
    .Q(\cpuregs.regs[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _16973_ (.CLK(clknet_leaf_101_clk),
    .D(_00147_),
    .Q(\cpuregs.regs[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _16974_ (.CLK(clknet_leaf_101_clk),
    .D(_00148_),
    .Q(\cpuregs.regs[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _16975_ (.CLK(clknet_leaf_120_clk),
    .D(_00149_),
    .Q(\cpuregs.regs[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _16976_ (.CLK(clknet_leaf_164_clk),
    .D(_00150_),
    .Q(\cpuregs.regs[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _16977_ (.CLK(clknet_leaf_161_clk),
    .D(_00151_),
    .Q(\cpuregs.regs[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _16978_ (.CLK(clknet_leaf_111_clk),
    .D(_00152_),
    .Q(\cpuregs.regs[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _16979_ (.CLK(clknet_leaf_166_clk),
    .D(_00153_),
    .Q(\cpuregs.regs[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _16980_ (.CLK(clknet_leaf_105_clk),
    .D(_00154_),
    .Q(\cpuregs.regs[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _16981_ (.CLK(clknet_leaf_119_clk),
    .D(_00155_),
    .Q(\cpuregs.regs[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _16982_ (.CLK(clknet_leaf_116_clk),
    .D(_00156_),
    .Q(\cpuregs.regs[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _16983_ (.CLK(clknet_leaf_163_clk),
    .D(_00157_),
    .Q(\cpuregs.regs[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _16984_ (.CLK(clknet_leaf_169_clk),
    .D(_00158_),
    .Q(\cpuregs.regs[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _16985_ (.CLK(clknet_leaf_172_clk),
    .D(_00159_),
    .Q(\cpuregs.regs[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16986_ (.CLK(clknet_leaf_189_clk),
    .D(_00160_),
    .Q(\cpuregs.regs[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16987_ (.CLK(clknet_leaf_12_clk),
    .D(_00161_),
    .Q(\cpuregs.regs[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16988_ (.CLK(clknet_leaf_3_clk),
    .D(_00162_),
    .Q(\cpuregs.regs[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16989_ (.CLK(clknet_leaf_1_clk),
    .D(_00163_),
    .Q(\cpuregs.regs[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16990_ (.CLK(clknet_leaf_170_clk),
    .D(_00164_),
    .Q(\cpuregs.regs[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16991_ (.CLK(clknet_leaf_181_clk),
    .D(_00165_),
    .Q(\cpuregs.regs[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16992_ (.CLK(clknet_leaf_186_clk),
    .D(_00166_),
    .Q(\cpuregs.regs[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16993_ (.CLK(clknet_leaf_183_clk),
    .D(_00167_),
    .Q(\cpuregs.regs[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16994_ (.CLK(clknet_leaf_181_clk),
    .D(_00168_),
    .Q(\cpuregs.regs[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16995_ (.CLK(clknet_leaf_131_clk),
    .D(_00169_),
    .Q(\cpuregs.regs[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16996_ (.CLK(clknet_leaf_158_clk),
    .D(_00170_),
    .Q(\cpuregs.regs[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16997_ (.CLK(clknet_leaf_157_clk),
    .D(_00171_),
    .Q(\cpuregs.regs[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16998_ (.CLK(clknet_leaf_139_clk),
    .D(_00172_),
    .Q(\cpuregs.regs[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16999_ (.CLK(clknet_leaf_147_clk),
    .D(_00173_),
    .Q(\cpuregs.regs[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17000_ (.CLK(clknet_leaf_142_clk),
    .D(_00174_),
    .Q(\cpuregs.regs[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17001_ (.CLK(clknet_leaf_141_clk),
    .D(_00175_),
    .Q(\cpuregs.regs[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17002_ (.CLK(clknet_leaf_139_clk),
    .D(_00176_),
    .Q(\cpuregs.regs[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17003_ (.CLK(clknet_leaf_154_clk),
    .D(_00177_),
    .Q(\cpuregs.regs[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17004_ (.CLK(clknet_leaf_180_clk),
    .D(_00178_),
    .Q(\cpuregs.regs[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17005_ (.CLK(clknet_leaf_120_clk),
    .D(_00179_),
    .Q(\cpuregs.regs[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17006_ (.CLK(clknet_leaf_123_clk),
    .D(_00180_),
    .Q(\cpuregs.regs[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17007_ (.CLK(clknet_leaf_124_clk),
    .D(_00181_),
    .Q(\cpuregs.regs[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17008_ (.CLK(clknet_leaf_164_clk),
    .D(_00182_),
    .Q(\cpuregs.regs[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17009_ (.CLK(clknet_leaf_160_clk),
    .D(_00183_),
    .Q(\cpuregs.regs[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17010_ (.CLK(clknet_leaf_111_clk),
    .D(_00184_),
    .Q(\cpuregs.regs[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17011_ (.CLK(clknet_leaf_20_clk),
    .D(_00185_),
    .Q(\cpuregs.regs[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17012_ (.CLK(clknet_leaf_112_clk),
    .D(_00186_),
    .Q(\cpuregs.regs[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17013_ (.CLK(clknet_leaf_117_clk),
    .D(_00187_),
    .Q(\cpuregs.regs[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17014_ (.CLK(clknet_leaf_126_clk),
    .D(_00188_),
    .Q(\cpuregs.regs[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17015_ (.CLK(clknet_leaf_177_clk),
    .D(_00189_),
    .Q(\cpuregs.regs[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17016_ (.CLK(clknet_leaf_169_clk),
    .D(_00190_),
    .Q(\cpuregs.regs[20][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17017_ (.CLK(clknet_leaf_172_clk),
    .D(_00191_),
    .Q(\cpuregs.regs[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17018_ (.CLK(clknet_leaf_190_clk),
    .D(_00192_),
    .Q(\cpuregs.regs[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17019_ (.CLK(clknet_leaf_2_clk),
    .D(_00193_),
    .Q(\cpuregs.regs[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17020_ (.CLK(clknet_leaf_3_clk),
    .D(_00194_),
    .Q(\cpuregs.regs[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17021_ (.CLK(clknet_leaf_1_clk),
    .D(_00195_),
    .Q(\cpuregs.regs[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17022_ (.CLK(clknet_leaf_171_clk),
    .D(_00196_),
    .Q(\cpuregs.regs[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17023_ (.CLK(clknet_leaf_181_clk),
    .D(_00197_),
    .Q(\cpuregs.regs[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17024_ (.CLK(clknet_leaf_186_clk),
    .D(_00198_),
    .Q(\cpuregs.regs[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17025_ (.CLK(clknet_leaf_183_clk),
    .D(_00199_),
    .Q(\cpuregs.regs[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17026_ (.CLK(clknet_leaf_181_clk),
    .D(_00200_),
    .Q(\cpuregs.regs[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17027_ (.CLK(clknet_leaf_130_clk),
    .D(_00201_),
    .Q(\cpuregs.regs[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17028_ (.CLK(clknet_leaf_157_clk),
    .D(_00202_),
    .Q(\cpuregs.regs[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17029_ (.CLK(clknet_leaf_156_clk),
    .D(_00203_),
    .Q(\cpuregs.regs[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17030_ (.CLK(clknet_leaf_139_clk),
    .D(_00204_),
    .Q(\cpuregs.regs[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17031_ (.CLK(clknet_leaf_147_clk),
    .D(_00205_),
    .Q(\cpuregs.regs[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17032_ (.CLK(clknet_leaf_142_clk),
    .D(_00206_),
    .Q(\cpuregs.regs[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17033_ (.CLK(clknet_leaf_141_clk),
    .D(_00207_),
    .Q(\cpuregs.regs[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17034_ (.CLK(clknet_leaf_139_clk),
    .D(_00208_),
    .Q(\cpuregs.regs[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17035_ (.CLK(clknet_leaf_177_clk),
    .D(_00209_),
    .Q(\cpuregs.regs[21][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17036_ (.CLK(clknet_leaf_180_clk),
    .D(_00210_),
    .Q(\cpuregs.regs[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17037_ (.CLK(clknet_leaf_120_clk),
    .D(_00211_),
    .Q(\cpuregs.regs[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17038_ (.CLK(clknet_leaf_123_clk),
    .D(_00212_),
    .Q(\cpuregs.regs[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17039_ (.CLK(clknet_leaf_124_clk),
    .D(_00213_),
    .Q(\cpuregs.regs[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17040_ (.CLK(clknet_leaf_164_clk),
    .D(_00214_),
    .Q(\cpuregs.regs[21][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17041_ (.CLK(clknet_leaf_160_clk),
    .D(_00215_),
    .Q(\cpuregs.regs[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17042_ (.CLK(clknet_leaf_111_clk),
    .D(_00216_),
    .Q(\cpuregs.regs[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17043_ (.CLK(clknet_leaf_20_clk),
    .D(_00217_),
    .Q(\cpuregs.regs[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17044_ (.CLK(clknet_leaf_112_clk),
    .D(_00218_),
    .Q(\cpuregs.regs[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17045_ (.CLK(clknet_leaf_116_clk),
    .D(_00219_),
    .Q(\cpuregs.regs[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17046_ (.CLK(clknet_leaf_126_clk),
    .D(_00220_),
    .Q(\cpuregs.regs[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17047_ (.CLK(clknet_leaf_169_clk),
    .D(_00221_),
    .Q(\cpuregs.regs[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17048_ (.CLK(clknet_leaf_176_clk),
    .D(_00222_),
    .Q(\cpuregs.regs[21][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17049_ (.CLK(clknet_leaf_13_clk),
    .D(_00223_),
    .Q(\cpuregs.regs[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17050_ (.CLK(clknet_leaf_190_clk),
    .D(_00224_),
    .Q(\cpuregs.regs[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17051_ (.CLK(clknet_leaf_3_clk),
    .D(_00225_),
    .Q(\cpuregs.regs[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17052_ (.CLK(clknet_leaf_3_clk),
    .D(_00226_),
    .Q(\cpuregs.regs[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17053_ (.CLK(clknet_leaf_1_clk),
    .D(_00227_),
    .Q(\cpuregs.regs[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17054_ (.CLK(clknet_leaf_172_clk),
    .D(_00228_),
    .Q(\cpuregs.regs[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17055_ (.CLK(clknet_leaf_181_clk),
    .D(_00229_),
    .Q(\cpuregs.regs[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17056_ (.CLK(clknet_leaf_186_clk),
    .D(_00230_),
    .Q(\cpuregs.regs[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17057_ (.CLK(clknet_leaf_183_clk),
    .D(_00231_),
    .Q(\cpuregs.regs[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17058_ (.CLK(clknet_leaf_183_clk),
    .D(_00232_),
    .Q(\cpuregs.regs[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17059_ (.CLK(clknet_leaf_142_clk),
    .D(_00233_),
    .Q(\cpuregs.regs[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17060_ (.CLK(clknet_leaf_157_clk),
    .D(_00234_),
    .Q(\cpuregs.regs[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17061_ (.CLK(clknet_leaf_156_clk),
    .D(_00235_),
    .Q(\cpuregs.regs[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17062_ (.CLK(clknet_leaf_139_clk),
    .D(_00236_),
    .Q(\cpuregs.regs[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17063_ (.CLK(clknet_leaf_147_clk),
    .D(_00237_),
    .Q(\cpuregs.regs[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17064_ (.CLK(clknet_leaf_144_clk),
    .D(_00238_),
    .Q(\cpuregs.regs[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17065_ (.CLK(clknet_leaf_142_clk),
    .D(_00239_),
    .Q(\cpuregs.regs[22][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17066_ (.CLK(clknet_leaf_139_clk),
    .D(_00240_),
    .Q(\cpuregs.regs[22][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17067_ (.CLK(clknet_leaf_178_clk),
    .D(_00241_),
    .Q(\cpuregs.regs[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17068_ (.CLK(clknet_leaf_180_clk),
    .D(_00242_),
    .Q(\cpuregs.regs[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17069_ (.CLK(clknet_leaf_120_clk),
    .D(_00243_),
    .Q(\cpuregs.regs[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17070_ (.CLK(clknet_leaf_123_clk),
    .D(_00244_),
    .Q(\cpuregs.regs[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17071_ (.CLK(clknet_leaf_122_clk),
    .D(_00245_),
    .Q(\cpuregs.regs[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17072_ (.CLK(clknet_leaf_164_clk),
    .D(_00246_),
    .Q(\cpuregs.regs[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17073_ (.CLK(clknet_leaf_162_clk),
    .D(_00247_),
    .Q(\cpuregs.regs[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17074_ (.CLK(clknet_leaf_110_clk),
    .D(_00248_),
    .Q(\cpuregs.regs[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17075_ (.CLK(clknet_leaf_19_clk),
    .D(_00249_),
    .Q(\cpuregs.regs[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17076_ (.CLK(clknet_leaf_112_clk),
    .D(_00250_),
    .Q(\cpuregs.regs[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17077_ (.CLK(clknet_leaf_116_clk),
    .D(_00251_),
    .Q(\cpuregs.regs[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17078_ (.CLK(clknet_leaf_127_clk),
    .D(_00252_),
    .Q(\cpuregs.regs[22][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17079_ (.CLK(clknet_leaf_177_clk),
    .D(_00253_),
    .Q(\cpuregs.regs[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17080_ (.CLK(clknet_leaf_176_clk),
    .D(_00254_),
    .Q(\cpuregs.regs[22][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17081_ (.CLK(clknet_leaf_13_clk),
    .D(_00255_),
    .Q(\cpuregs.regs[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17082_ (.CLK(clknet_leaf_189_clk),
    .D(_00256_),
    .Q(\cpuregs.regs[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17083_ (.CLK(clknet_leaf_3_clk),
    .D(_00257_),
    .Q(\cpuregs.regs[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17084_ (.CLK(clknet_leaf_3_clk),
    .D(_00258_),
    .Q(\cpuregs.regs[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17085_ (.CLK(clknet_leaf_1_clk),
    .D(_00259_),
    .Q(\cpuregs.regs[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17086_ (.CLK(clknet_leaf_172_clk),
    .D(_00260_),
    .Q(\cpuregs.regs[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17087_ (.CLK(clknet_leaf_181_clk),
    .D(_00261_),
    .Q(\cpuregs.regs[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17088_ (.CLK(clknet_leaf_186_clk),
    .D(_00262_),
    .Q(\cpuregs.regs[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17089_ (.CLK(clknet_leaf_183_clk),
    .D(_00263_),
    .Q(\cpuregs.regs[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17090_ (.CLK(clknet_leaf_181_clk),
    .D(_00264_),
    .Q(\cpuregs.regs[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17091_ (.CLK(clknet_leaf_143_clk),
    .D(_00265_),
    .Q(\cpuregs.regs[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17092_ (.CLK(clknet_leaf_157_clk),
    .D(_00266_),
    .Q(\cpuregs.regs[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17093_ (.CLK(clknet_leaf_156_clk),
    .D(_00267_),
    .Q(\cpuregs.regs[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17094_ (.CLK(clknet_leaf_139_clk),
    .D(_00268_),
    .Q(\cpuregs.regs[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17095_ (.CLK(clknet_leaf_147_clk),
    .D(_00269_),
    .Q(\cpuregs.regs[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17096_ (.CLK(clknet_leaf_142_clk),
    .D(_00270_),
    .Q(\cpuregs.regs[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17097_ (.CLK(clknet_leaf_142_clk),
    .D(_00271_),
    .Q(\cpuregs.regs[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17098_ (.CLK(clknet_leaf_139_clk),
    .D(_00272_),
    .Q(\cpuregs.regs[23][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17099_ (.CLK(clknet_leaf_177_clk),
    .D(_00273_),
    .Q(\cpuregs.regs[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17100_ (.CLK(clknet_leaf_180_clk),
    .D(_00274_),
    .Q(\cpuregs.regs[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17101_ (.CLK(clknet_leaf_120_clk),
    .D(_00275_),
    .Q(\cpuregs.regs[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17102_ (.CLK(clknet_leaf_122_clk),
    .D(_00276_),
    .Q(\cpuregs.regs[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17103_ (.CLK(clknet_leaf_124_clk),
    .D(_00277_),
    .Q(\cpuregs.regs[23][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17104_ (.CLK(clknet_leaf_164_clk),
    .D(_00278_),
    .Q(\cpuregs.regs[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17105_ (.CLK(clknet_leaf_162_clk),
    .D(_00279_),
    .Q(\cpuregs.regs[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17106_ (.CLK(clknet_leaf_111_clk),
    .D(_00280_),
    .Q(\cpuregs.regs[23][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17107_ (.CLK(clknet_leaf_19_clk),
    .D(_00281_),
    .Q(\cpuregs.regs[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17108_ (.CLK(clknet_leaf_112_clk),
    .D(_00282_),
    .Q(\cpuregs.regs[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17109_ (.CLK(clknet_leaf_116_clk),
    .D(_00283_),
    .Q(\cpuregs.regs[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17110_ (.CLK(clknet_leaf_127_clk),
    .D(_00284_),
    .Q(\cpuregs.regs[23][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17111_ (.CLK(clknet_leaf_177_clk),
    .D(_00285_),
    .Q(\cpuregs.regs[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17112_ (.CLK(clknet_leaf_176_clk),
    .D(_00286_),
    .Q(\cpuregs.regs[23][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17113_ (.CLK(clknet_leaf_171_clk),
    .D(_00287_),
    .Q(\cpuregs.regs[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17114_ (.CLK(clknet_leaf_187_clk),
    .D(_00288_),
    .Q(\cpuregs.regs[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17115_ (.CLK(clknet_leaf_12_clk),
    .D(_00289_),
    .Q(\cpuregs.regs[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17116_ (.CLK(clknet_leaf_12_clk),
    .D(_00290_),
    .Q(\cpuregs.regs[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17117_ (.CLK(clknet_leaf_13_clk),
    .D(_00291_),
    .Q(\cpuregs.regs[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17118_ (.CLK(clknet_leaf_167_clk),
    .D(_00292_),
    .Q(\cpuregs.regs[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17119_ (.CLK(clknet_leaf_179_clk),
    .D(_00293_),
    .Q(\cpuregs.regs[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17120_ (.CLK(clknet_leaf_174_clk),
    .D(_00294_),
    .Q(\cpuregs.regs[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17121_ (.CLK(clknet_leaf_184_clk),
    .D(_00295_),
    .Q(\cpuregs.regs[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17122_ (.CLK(clknet_leaf_185_clk),
    .D(_00296_),
    .Q(\cpuregs.regs[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17123_ (.CLK(clknet_leaf_134_clk),
    .D(_00297_),
    .Q(\cpuregs.regs[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17124_ (.CLK(clknet_leaf_143_clk),
    .D(_00298_),
    .Q(\cpuregs.regs[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17125_ (.CLK(clknet_leaf_148_clk),
    .D(_00299_),
    .Q(\cpuregs.regs[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17126_ (.CLK(clknet_leaf_137_clk),
    .D(_00300_),
    .Q(\cpuregs.regs[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17127_ (.CLK(clknet_leaf_142_clk),
    .D(_00301_),
    .Q(\cpuregs.regs[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17128_ (.CLK(clknet_leaf_134_clk),
    .D(_00302_),
    .Q(\cpuregs.regs[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17129_ (.CLK(clknet_leaf_134_clk),
    .D(_00303_),
    .Q(\cpuregs.regs[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17130_ (.CLK(clknet_leaf_147_clk),
    .D(_00304_),
    .Q(\cpuregs.regs[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17131_ (.CLK(clknet_leaf_149_clk),
    .D(_00305_),
    .Q(\cpuregs.regs[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17132_ (.CLK(clknet_leaf_149_clk),
    .D(_00306_),
    .Q(\cpuregs.regs[24][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17133_ (.CLK(clknet_leaf_123_clk),
    .D(_00307_),
    .Q(\cpuregs.regs[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17134_ (.CLK(clknet_leaf_123_clk),
    .D(_00308_),
    .Q(\cpuregs.regs[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17135_ (.CLK(clknet_leaf_124_clk),
    .D(_00309_),
    .Q(\cpuregs.regs[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17136_ (.CLK(clknet_leaf_110_clk),
    .D(_00310_),
    .Q(\cpuregs.regs[24][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17137_ (.CLK(clknet_leaf_115_clk),
    .D(_00311_),
    .Q(\cpuregs.regs[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17138_ (.CLK(clknet_leaf_113_clk),
    .D(_00312_),
    .Q(\cpuregs.regs[24][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17139_ (.CLK(clknet_leaf_109_clk),
    .D(_00313_),
    .Q(\cpuregs.regs[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17140_ (.CLK(clknet_leaf_120_clk),
    .D(_00314_),
    .Q(\cpuregs.regs[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17141_ (.CLK(clknet_leaf_116_clk),
    .D(_00315_),
    .Q(\cpuregs.regs[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17142_ (.CLK(clknet_leaf_126_clk),
    .D(_00316_),
    .Q(\cpuregs.regs[24][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17143_ (.CLK(clknet_leaf_156_clk),
    .D(_00317_),
    .Q(\cpuregs.regs[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17144_ (.CLK(clknet_leaf_176_clk),
    .D(_00318_),
    .Q(\cpuregs.regs[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17145_ (.CLK(clknet_leaf_15_clk),
    .D(_00319_),
    .Q(\cpuregs.regs[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17146_ (.CLK(clknet_leaf_187_clk),
    .D(_00320_),
    .Q(\cpuregs.regs[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17147_ (.CLK(clknet_leaf_12_clk),
    .D(_00321_),
    .Q(\cpuregs.regs[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17148_ (.CLK(clknet_leaf_12_clk),
    .D(_00322_),
    .Q(\cpuregs.regs[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17149_ (.CLK(clknet_leaf_2_clk),
    .D(_00323_),
    .Q(\cpuregs.regs[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17150_ (.CLK(clknet_leaf_167_clk),
    .D(_00324_),
    .Q(\cpuregs.regs[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17151_ (.CLK(clknet_leaf_179_clk),
    .D(_00325_),
    .Q(\cpuregs.regs[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17152_ (.CLK(clknet_leaf_174_clk),
    .D(_00326_),
    .Q(\cpuregs.regs[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17153_ (.CLK(clknet_leaf_184_clk),
    .D(_00327_),
    .Q(\cpuregs.regs[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17154_ (.CLK(clknet_leaf_185_clk),
    .D(_00328_),
    .Q(\cpuregs.regs[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17155_ (.CLK(clknet_leaf_134_clk),
    .D(_00329_),
    .Q(\cpuregs.regs[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17156_ (.CLK(clknet_leaf_143_clk),
    .D(_00330_),
    .Q(\cpuregs.regs[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17157_ (.CLK(clknet_leaf_148_clk),
    .D(_00331_),
    .Q(\cpuregs.regs[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17158_ (.CLK(clknet_leaf_137_clk),
    .D(_00332_),
    .Q(\cpuregs.regs[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17159_ (.CLK(clknet_leaf_144_clk),
    .D(_00333_),
    .Q(\cpuregs.regs[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17160_ (.CLK(clknet_leaf_133_clk),
    .D(_00334_),
    .Q(\cpuregs.regs[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17161_ (.CLK(clknet_leaf_134_clk),
    .D(_00335_),
    .Q(\cpuregs.regs[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17162_ (.CLK(clknet_leaf_147_clk),
    .D(_00336_),
    .Q(\cpuregs.regs[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17163_ (.CLK(clknet_leaf_150_clk),
    .D(_00337_),
    .Q(\cpuregs.regs[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17164_ (.CLK(clknet_leaf_149_clk),
    .D(_00338_),
    .Q(\cpuregs.regs[25][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17165_ (.CLK(clknet_leaf_123_clk),
    .D(_00339_),
    .Q(\cpuregs.regs[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17166_ (.CLK(clknet_leaf_123_clk),
    .D(_00340_),
    .Q(\cpuregs.regs[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17167_ (.CLK(clknet_leaf_124_clk),
    .D(_00341_),
    .Q(\cpuregs.regs[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17168_ (.CLK(clknet_leaf_110_clk),
    .D(_00342_),
    .Q(\cpuregs.regs[25][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17169_ (.CLK(clknet_leaf_115_clk),
    .D(_00343_),
    .Q(\cpuregs.regs[25][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17170_ (.CLK(clknet_leaf_114_clk),
    .D(_00344_),
    .Q(\cpuregs.regs[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17171_ (.CLK(clknet_leaf_109_clk),
    .D(_00345_),
    .Q(\cpuregs.regs[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17172_ (.CLK(clknet_leaf_120_clk),
    .D(_00346_),
    .Q(\cpuregs.regs[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17173_ (.CLK(clknet_leaf_116_clk),
    .D(_00347_),
    .Q(\cpuregs.regs[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17174_ (.CLK(clknet_leaf_126_clk),
    .D(_00348_),
    .Q(\cpuregs.regs[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17175_ (.CLK(clknet_leaf_156_clk),
    .D(_00349_),
    .Q(\cpuregs.regs[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17176_ (.CLK(clknet_leaf_176_clk),
    .D(_00350_),
    .Q(\cpuregs.regs[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17177_ (.CLK(clknet_leaf_14_clk),
    .D(_00351_),
    .Q(\cpuregs.regs[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17178_ (.CLK(clknet_leaf_188_clk),
    .D(_00352_),
    .Q(\cpuregs.regs[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17179_ (.CLK(clknet_leaf_12_clk),
    .D(_00353_),
    .Q(\cpuregs.regs[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17180_ (.CLK(clknet_leaf_12_clk),
    .D(_00354_),
    .Q(\cpuregs.regs[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17181_ (.CLK(clknet_leaf_2_clk),
    .D(_00355_),
    .Q(\cpuregs.regs[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17182_ (.CLK(clknet_leaf_167_clk),
    .D(_00356_),
    .Q(\cpuregs.regs[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17183_ (.CLK(clknet_leaf_179_clk),
    .D(_00357_),
    .Q(\cpuregs.regs[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17184_ (.CLK(clknet_leaf_174_clk),
    .D(_00358_),
    .Q(\cpuregs.regs[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17185_ (.CLK(clknet_leaf_189_clk),
    .D(_00359_),
    .Q(\cpuregs.regs[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17186_ (.CLK(clknet_leaf_185_clk),
    .D(_00360_),
    .Q(\cpuregs.regs[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17187_ (.CLK(clknet_leaf_133_clk),
    .D(_00361_),
    .Q(\cpuregs.regs[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17188_ (.CLK(clknet_leaf_159_clk),
    .D(_00362_),
    .Q(\cpuregs.regs[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17189_ (.CLK(clknet_leaf_148_clk),
    .D(_00363_),
    .Q(\cpuregs.regs[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17190_ (.CLK(clknet_leaf_137_clk),
    .D(_00364_),
    .Q(\cpuregs.regs[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17191_ (.CLK(clknet_leaf_144_clk),
    .D(_00365_),
    .Q(\cpuregs.regs[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17192_ (.CLK(clknet_leaf_133_clk),
    .D(_00366_),
    .Q(\cpuregs.regs[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17193_ (.CLK(clknet_leaf_135_clk),
    .D(_00367_),
    .Q(\cpuregs.regs[26][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17194_ (.CLK(clknet_leaf_147_clk),
    .D(_00368_),
    .Q(\cpuregs.regs[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17195_ (.CLK(clknet_leaf_150_clk),
    .D(_00369_),
    .Q(\cpuregs.regs[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17196_ (.CLK(clknet_leaf_151_clk),
    .D(_00370_),
    .Q(\cpuregs.regs[26][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17197_ (.CLK(clknet_leaf_121_clk),
    .D(_00371_),
    .Q(\cpuregs.regs[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17198_ (.CLK(clknet_leaf_123_clk),
    .D(_00372_),
    .Q(\cpuregs.regs[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17199_ (.CLK(clknet_leaf_124_clk),
    .D(_00373_),
    .Q(\cpuregs.regs[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17200_ (.CLK(clknet_leaf_110_clk),
    .D(_00374_),
    .Q(\cpuregs.regs[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17201_ (.CLK(clknet_leaf_160_clk),
    .D(_00375_),
    .Q(\cpuregs.regs[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17202_ (.CLK(clknet_leaf_111_clk),
    .D(_00376_),
    .Q(\cpuregs.regs[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17203_ (.CLK(clknet_leaf_109_clk),
    .D(_00377_),
    .Q(\cpuregs.regs[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17204_ (.CLK(clknet_leaf_113_clk),
    .D(_00378_),
    .Q(\cpuregs.regs[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17205_ (.CLK(clknet_leaf_115_clk),
    .D(_00379_),
    .Q(\cpuregs.regs[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17206_ (.CLK(clknet_leaf_125_clk),
    .D(_00380_),
    .Q(\cpuregs.regs[26][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17207_ (.CLK(clknet_leaf_155_clk),
    .D(_00381_),
    .Q(\cpuregs.regs[26][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17208_ (.CLK(clknet_leaf_176_clk),
    .D(_00382_),
    .Q(\cpuregs.regs[26][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17209_ (.CLK(clknet_leaf_14_clk),
    .D(_00383_),
    .Q(\cpuregs.regs[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17210_ (.CLK(clknet_leaf_188_clk),
    .D(_00384_),
    .Q(\cpuregs.regs[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17211_ (.CLK(clknet_leaf_12_clk),
    .D(_00385_),
    .Q(\cpuregs.regs[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17212_ (.CLK(clknet_leaf_12_clk),
    .D(_00386_),
    .Q(\cpuregs.regs[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17213_ (.CLK(clknet_leaf_2_clk),
    .D(_00387_),
    .Q(\cpuregs.regs[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17214_ (.CLK(clknet_leaf_167_clk),
    .D(_00388_),
    .Q(\cpuregs.regs[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17215_ (.CLK(clknet_leaf_179_clk),
    .D(_00389_),
    .Q(\cpuregs.regs[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17216_ (.CLK(clknet_leaf_174_clk),
    .D(_00390_),
    .Q(\cpuregs.regs[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17217_ (.CLK(clknet_leaf_189_clk),
    .D(_00391_),
    .Q(\cpuregs.regs[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17218_ (.CLK(clknet_leaf_185_clk),
    .D(_00392_),
    .Q(\cpuregs.regs[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17219_ (.CLK(clknet_leaf_133_clk),
    .D(_00393_),
    .Q(\cpuregs.regs[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17220_ (.CLK(clknet_leaf_159_clk),
    .D(_00394_),
    .Q(\cpuregs.regs[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17221_ (.CLK(clknet_leaf_148_clk),
    .D(_00395_),
    .Q(\cpuregs.regs[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17222_ (.CLK(clknet_leaf_137_clk),
    .D(_00396_),
    .Q(\cpuregs.regs[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17223_ (.CLK(clknet_leaf_144_clk),
    .D(_00397_),
    .Q(\cpuregs.regs[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17224_ (.CLK(clknet_leaf_133_clk),
    .D(_00398_),
    .Q(\cpuregs.regs[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17225_ (.CLK(clknet_leaf_135_clk),
    .D(_00399_),
    .Q(\cpuregs.regs[27][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17226_ (.CLK(clknet_leaf_147_clk),
    .D(_00400_),
    .Q(\cpuregs.regs[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17227_ (.CLK(clknet_leaf_150_clk),
    .D(_00401_),
    .Q(\cpuregs.regs[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17228_ (.CLK(clknet_leaf_151_clk),
    .D(_00402_),
    .Q(\cpuregs.regs[27][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17229_ (.CLK(clknet_leaf_121_clk),
    .D(_00403_),
    .Q(\cpuregs.regs[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17230_ (.CLK(clknet_leaf_123_clk),
    .D(_00404_),
    .Q(\cpuregs.regs[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17231_ (.CLK(clknet_leaf_124_clk),
    .D(_00405_),
    .Q(\cpuregs.regs[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17232_ (.CLK(clknet_leaf_110_clk),
    .D(_00406_),
    .Q(\cpuregs.regs[27][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17233_ (.CLK(clknet_leaf_160_clk),
    .D(_00407_),
    .Q(\cpuregs.regs[27][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17234_ (.CLK(clknet_leaf_114_clk),
    .D(_00408_),
    .Q(\cpuregs.regs[27][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17235_ (.CLK(clknet_leaf_109_clk),
    .D(_00409_),
    .Q(\cpuregs.regs[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17236_ (.CLK(clknet_leaf_120_clk),
    .D(_00410_),
    .Q(\cpuregs.regs[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17237_ (.CLK(clknet_leaf_115_clk),
    .D(_00411_),
    .Q(\cpuregs.regs[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17238_ (.CLK(clknet_leaf_125_clk),
    .D(_00412_),
    .Q(\cpuregs.regs[27][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17239_ (.CLK(clknet_leaf_155_clk),
    .D(_00413_),
    .Q(\cpuregs.regs[27][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17240_ (.CLK(clknet_leaf_176_clk),
    .D(_00414_),
    .Q(\cpuregs.regs[27][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17241_ (.CLK(clknet_leaf_15_clk),
    .D(_00415_),
    .Q(\cpuregs.regs[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17242_ (.CLK(clknet_leaf_186_clk),
    .D(_00416_),
    .Q(\cpuregs.regs[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17243_ (.CLK(clknet_leaf_13_clk),
    .D(_00417_),
    .Q(\cpuregs.regs[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17244_ (.CLK(clknet_leaf_13_clk),
    .D(_00418_),
    .Q(\cpuregs.regs[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17245_ (.CLK(clknet_leaf_187_clk),
    .D(_00419_),
    .Q(\cpuregs.regs[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17246_ (.CLK(clknet_leaf_166_clk),
    .D(_00420_),
    .Q(\cpuregs.regs[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17247_ (.CLK(clknet_leaf_181_clk),
    .D(_00421_),
    .Q(\cpuregs.regs[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17248_ (.CLK(clknet_leaf_175_clk),
    .D(_00422_),
    .Q(\cpuregs.regs[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17249_ (.CLK(clknet_leaf_183_clk),
    .D(_00423_),
    .Q(\cpuregs.regs[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17250_ (.CLK(clknet_leaf_183_clk),
    .D(_00424_),
    .Q(\cpuregs.regs[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17251_ (.CLK(clknet_leaf_132_clk),
    .D(_00425_),
    .Q(\cpuregs.regs[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17252_ (.CLK(clknet_leaf_143_clk),
    .D(_00426_),
    .Q(\cpuregs.regs[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17253_ (.CLK(clknet_leaf_148_clk),
    .D(_00427_),
    .Q(\cpuregs.regs[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17254_ (.CLK(clknet_leaf_137_clk),
    .D(_00428_),
    .Q(\cpuregs.regs[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17255_ (.CLK(clknet_leaf_142_clk),
    .D(_00429_),
    .Q(\cpuregs.regs[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17256_ (.CLK(clknet_leaf_132_clk),
    .D(_00430_),
    .Q(\cpuregs.regs[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17257_ (.CLK(clknet_leaf_135_clk),
    .D(_00431_),
    .Q(\cpuregs.regs[28][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17258_ (.CLK(clknet_leaf_140_clk),
    .D(_00432_),
    .Q(\cpuregs.regs[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17259_ (.CLK(clknet_leaf_150_clk),
    .D(_00433_),
    .Q(\cpuregs.regs[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17260_ (.CLK(clknet_leaf_151_clk),
    .D(_00434_),
    .Q(\cpuregs.regs[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17261_ (.CLK(clknet_leaf_97_clk),
    .D(_00435_),
    .Q(\cpuregs.regs[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17262_ (.CLK(clknet_leaf_97_clk),
    .D(_00436_),
    .Q(\cpuregs.regs[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17263_ (.CLK(clknet_leaf_122_clk),
    .D(_00437_),
    .Q(\cpuregs.regs[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17264_ (.CLK(clknet_leaf_110_clk),
    .D(_00438_),
    .Q(\cpuregs.regs[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17265_ (.CLK(clknet_leaf_160_clk),
    .D(_00439_),
    .Q(\cpuregs.regs[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17266_ (.CLK(clknet_leaf_113_clk),
    .D(_00440_),
    .Q(\cpuregs.regs[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17267_ (.CLK(clknet_leaf_165_clk),
    .D(_00441_),
    .Q(\cpuregs.regs[28][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17268_ (.CLK(clknet_leaf_113_clk),
    .D(_00442_),
    .Q(\cpuregs.regs[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17269_ (.CLK(clknet_leaf_115_clk),
    .D(_00443_),
    .Q(\cpuregs.regs[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17270_ (.CLK(clknet_leaf_125_clk),
    .D(_00444_),
    .Q(\cpuregs.regs[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17271_ (.CLK(clknet_leaf_155_clk),
    .D(_00445_),
    .Q(\cpuregs.regs[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17272_ (.CLK(clknet_leaf_177_clk),
    .D(_00446_),
    .Q(\cpuregs.regs[28][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17273_ (.CLK(clknet_leaf_17_clk),
    .D(_00447_),
    .Q(\cpuregs.regs[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17274_ (.CLK(clknet_leaf_188_clk),
    .D(_00448_),
    .Q(\cpuregs.regs[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17275_ (.CLK(clknet_leaf_16_clk),
    .D(_00449_),
    .Q(\cpuregs.regs[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17276_ (.CLK(clknet_leaf_7_clk),
    .D(_00450_),
    .Q(\cpuregs.regs[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17277_ (.CLK(clknet_leaf_2_clk),
    .D(_00451_),
    .Q(\cpuregs.regs[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17278_ (.CLK(clknet_leaf_17_clk),
    .D(_00452_),
    .Q(\cpuregs.regs[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17279_ (.CLK(clknet_leaf_176_clk),
    .D(_00453_),
    .Q(\cpuregs.regs[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17280_ (.CLK(clknet_leaf_13_clk),
    .D(_00454_),
    .Q(\cpuregs.regs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17281_ (.CLK(clknet_leaf_186_clk),
    .D(_00455_),
    .Q(\cpuregs.regs[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17282_ (.CLK(clknet_leaf_175_clk),
    .D(_00456_),
    .Q(\cpuregs.regs[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17283_ (.CLK(clknet_leaf_126_clk),
    .D(_00457_),
    .Q(\cpuregs.regs[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17284_ (.CLK(clknet_leaf_160_clk),
    .D(_00458_),
    .Q(\cpuregs.regs[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17285_ (.CLK(clknet_leaf_153_clk),
    .D(_00459_),
    .Q(\cpuregs.regs[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17286_ (.CLK(clknet_leaf_136_clk),
    .D(_00460_),
    .Q(\cpuregs.regs[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17287_ (.CLK(clknet_leaf_157_clk),
    .D(_00461_),
    .Q(\cpuregs.regs[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17288_ (.CLK(clknet_leaf_115_clk),
    .D(_00462_),
    .Q(\cpuregs.regs[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17289_ (.CLK(clknet_leaf_135_clk),
    .D(_00463_),
    .Q(\cpuregs.regs[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17290_ (.CLK(clknet_leaf_144_clk),
    .D(_00464_),
    .Q(\cpuregs.regs[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17291_ (.CLK(clknet_leaf_154_clk),
    .D(_00465_),
    .Q(\cpuregs.regs[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17292_ (.CLK(clknet_leaf_152_clk),
    .D(_00466_),
    .Q(\cpuregs.regs[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17293_ (.CLK(clknet_leaf_100_clk),
    .D(_00467_),
    .Q(\cpuregs.regs[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17294_ (.CLK(clknet_leaf_98_clk),
    .D(_00468_),
    .Q(\cpuregs.regs[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17295_ (.CLK(clknet_leaf_119_clk),
    .D(_00469_),
    .Q(\cpuregs.regs[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17296_ (.CLK(clknet_leaf_165_clk),
    .D(_00470_),
    .Q(\cpuregs.regs[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17297_ (.CLK(clknet_leaf_114_clk),
    .D(_00471_),
    .Q(\cpuregs.regs[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17298_ (.CLK(clknet_leaf_109_clk),
    .D(_00472_),
    .Q(\cpuregs.regs[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17299_ (.CLK(clknet_leaf_166_clk),
    .D(_00473_),
    .Q(\cpuregs.regs[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17300_ (.CLK(clknet_leaf_105_clk),
    .D(_00474_),
    .Q(\cpuregs.regs[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17301_ (.CLK(clknet_leaf_113_clk),
    .D(_00475_),
    .Q(\cpuregs.regs[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17302_ (.CLK(clknet_leaf_128_clk),
    .D(_00476_),
    .Q(\cpuregs.regs[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17303_ (.CLK(clknet_leaf_162_clk),
    .D(_00477_),
    .Q(\cpuregs.regs[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17304_ (.CLK(clknet_leaf_170_clk),
    .D(_00478_),
    .Q(\cpuregs.regs[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17305_ (.CLK(clknet_leaf_15_clk),
    .D(_00479_),
    .Q(\cpuregs.regs[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17306_ (.CLK(clknet_leaf_188_clk),
    .D(_00480_),
    .Q(\cpuregs.regs[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17307_ (.CLK(clknet_leaf_13_clk),
    .D(_00481_),
    .Q(\cpuregs.regs[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17308_ (.CLK(clknet_leaf_12_clk),
    .D(_00482_),
    .Q(\cpuregs.regs[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17309_ (.CLK(clknet_leaf_2_clk),
    .D(_00483_),
    .Q(\cpuregs.regs[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17310_ (.CLK(clknet_leaf_166_clk),
    .D(_00484_),
    .Q(\cpuregs.regs[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17311_ (.CLK(clknet_leaf_181_clk),
    .D(_00485_),
    .Q(\cpuregs.regs[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17312_ (.CLK(clknet_leaf_175_clk),
    .D(_00486_),
    .Q(\cpuregs.regs[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17313_ (.CLK(clknet_leaf_184_clk),
    .D(_00487_),
    .Q(\cpuregs.regs[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17314_ (.CLK(clknet_leaf_183_clk),
    .D(_00488_),
    .Q(\cpuregs.regs[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17315_ (.CLK(clknet_leaf_131_clk),
    .D(_00489_),
    .Q(\cpuregs.regs[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17316_ (.CLK(clknet_leaf_159_clk),
    .D(_00490_),
    .Q(\cpuregs.regs[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17317_ (.CLK(clknet_leaf_148_clk),
    .D(_00491_),
    .Q(\cpuregs.regs[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17318_ (.CLK(clknet_leaf_138_clk),
    .D(_00492_),
    .Q(\cpuregs.regs[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17319_ (.CLK(clknet_leaf_145_clk),
    .D(_00493_),
    .Q(\cpuregs.regs[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17320_ (.CLK(clknet_leaf_132_clk),
    .D(_00494_),
    .Q(\cpuregs.regs[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17321_ (.CLK(clknet_leaf_132_clk),
    .D(_00495_),
    .Q(\cpuregs.regs[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17322_ (.CLK(clknet_leaf_139_clk),
    .D(_00496_),
    .Q(\cpuregs.regs[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17323_ (.CLK(clknet_leaf_151_clk),
    .D(_00497_),
    .Q(\cpuregs.regs[30][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17324_ (.CLK(clknet_leaf_151_clk),
    .D(_00498_),
    .Q(\cpuregs.regs[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17325_ (.CLK(clknet_leaf_98_clk),
    .D(_00499_),
    .Q(\cpuregs.regs[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17326_ (.CLK(clknet_leaf_97_clk),
    .D(_00500_),
    .Q(\cpuregs.regs[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17327_ (.CLK(clknet_leaf_121_clk),
    .D(_00501_),
    .Q(\cpuregs.regs[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17328_ (.CLK(clknet_leaf_164_clk),
    .D(_00502_),
    .Q(\cpuregs.regs[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17329_ (.CLK(clknet_leaf_161_clk),
    .D(_00503_),
    .Q(\cpuregs.regs[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17330_ (.CLK(clknet_leaf_111_clk),
    .D(_00504_),
    .Q(\cpuregs.regs[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17331_ (.CLK(clknet_leaf_165_clk),
    .D(_00505_),
    .Q(\cpuregs.regs[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17332_ (.CLK(clknet_leaf_112_clk),
    .D(_00506_),
    .Q(\cpuregs.regs[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17333_ (.CLK(clknet_leaf_115_clk),
    .D(_00507_),
    .Q(\cpuregs.regs[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17334_ (.CLK(clknet_leaf_128_clk),
    .D(_00508_),
    .Q(\cpuregs.regs[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17335_ (.CLK(clknet_leaf_177_clk),
    .D(_00509_),
    .Q(\cpuregs.regs[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17336_ (.CLK(clknet_leaf_176_clk),
    .D(_00510_),
    .Q(\cpuregs.regs[30][31] ));
 sky130_fd_sc_hd__dfxtp_2 _17337_ (.CLK(clknet_leaf_17_clk),
    .D(_00084_),
    .Q(_00064_));
 sky130_fd_sc_hd__dfxtp_2 _17338_ (.CLK(clknet_leaf_17_clk),
    .D(_00085_),
    .Q(_00065_));
 sky130_fd_sc_hd__dfxtp_1 _17339_ (.CLK(clknet_leaf_17_clk),
    .D(_00086_),
    .Q(_00066_));
 sky130_fd_sc_hd__dfxtp_4 _17340_ (.CLK(clknet_leaf_16_clk),
    .D(_00087_),
    .Q(_00067_));
 sky130_fd_sc_hd__dfxtp_4 _17341_ (.CLK(clknet_leaf_16_clk),
    .D(_00088_),
    .Q(_00068_));
 sky130_fd_sc_hd__dfxtp_1 _17342_ (.CLK(clknet_leaf_18_clk),
    .D(_00511_),
    .Q(\cpuregs.regs[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17343_ (.CLK(clknet_leaf_189_clk),
    .D(_00512_),
    .Q(\cpuregs.regs[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17344_ (.CLK(clknet_leaf_10_clk),
    .D(_00513_),
    .Q(\cpuregs.regs[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17345_ (.CLK(clknet_leaf_10_clk),
    .D(_00514_),
    .Q(\cpuregs.regs[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17346_ (.CLK(clknet_leaf_187_clk),
    .D(_00515_),
    .Q(\cpuregs.regs[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17347_ (.CLK(clknet_leaf_18_clk),
    .D(_00516_),
    .Q(\cpuregs.regs[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17348_ (.CLK(clknet_leaf_180_clk),
    .D(_00517_),
    .Q(\cpuregs.regs[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17349_ (.CLK(clknet_leaf_174_clk),
    .D(_00518_),
    .Q(\cpuregs.regs[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17350_ (.CLK(clknet_leaf_185_clk),
    .D(_00519_),
    .Q(\cpuregs.regs[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17351_ (.CLK(clknet_leaf_182_clk),
    .D(_00520_),
    .Q(\cpuregs.regs[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17352_ (.CLK(clknet_leaf_133_clk),
    .D(_00521_),
    .Q(\cpuregs.regs[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17353_ (.CLK(clknet_leaf_159_clk),
    .D(_00522_),
    .Q(\cpuregs.regs[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17354_ (.CLK(clknet_leaf_148_clk),
    .D(_00523_),
    .Q(\cpuregs.regs[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17355_ (.CLK(clknet_leaf_139_clk),
    .D(_00524_),
    .Q(\cpuregs.regs[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17356_ (.CLK(clknet_leaf_147_clk),
    .D(_00525_),
    .Q(\cpuregs.regs[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17357_ (.CLK(clknet_leaf_127_clk),
    .D(_00526_),
    .Q(\cpuregs.regs[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17358_ (.CLK(clknet_leaf_132_clk),
    .D(_00527_),
    .Q(\cpuregs.regs[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17359_ (.CLK(clknet_leaf_139_clk),
    .D(_00528_),
    .Q(\cpuregs.regs[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17360_ (.CLK(clknet_leaf_154_clk),
    .D(_00529_),
    .Q(\cpuregs.regs[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17361_ (.CLK(clknet_leaf_151_clk),
    .D(_00530_),
    .Q(\cpuregs.regs[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17362_ (.CLK(clknet_leaf_99_clk),
    .D(_00531_),
    .Q(\cpuregs.regs[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17363_ (.CLK(clknet_leaf_98_clk),
    .D(_00532_),
    .Q(\cpuregs.regs[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17364_ (.CLK(clknet_leaf_122_clk),
    .D(_00533_),
    .Q(\cpuregs.regs[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17365_ (.CLK(clknet_leaf_164_clk),
    .D(_00534_),
    .Q(\cpuregs.regs[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17366_ (.CLK(clknet_leaf_114_clk),
    .D(_00535_),
    .Q(\cpuregs.regs[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17367_ (.CLK(clknet_leaf_111_clk),
    .D(_00536_),
    .Q(\cpuregs.regs[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17368_ (.CLK(clknet_leaf_164_clk),
    .D(_00537_),
    .Q(\cpuregs.regs[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17369_ (.CLK(clknet_leaf_100_clk),
    .D(_00538_),
    .Q(\cpuregs.regs[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17370_ (.CLK(clknet_leaf_119_clk),
    .D(_00539_),
    .Q(\cpuregs.regs[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17371_ (.CLK(clknet_leaf_128_clk),
    .D(_00540_),
    .Q(\cpuregs.regs[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17372_ (.CLK(clknet_leaf_163_clk),
    .D(_00541_),
    .Q(\cpuregs.regs[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17373_ (.CLK(clknet_leaf_163_clk),
    .D(_00542_),
    .Q(\cpuregs.regs[12][31] ));
 sky130_fd_sc_hd__dfxtp_4 _17374_ (.CLK(clknet_leaf_20_clk),
    .D(_00543_),
    .Q(\cpuregs.waddr[0] ));
 sky130_fd_sc_hd__dfxtp_4 _17375_ (.CLK(clknet_leaf_21_clk),
    .D(_00544_),
    .Q(\cpuregs.waddr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _17376_ (.CLK(clknet_leaf_21_clk),
    .D(_00545_),
    .Q(\cpuregs.waddr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _17377_ (.CLK(clknet_leaf_17_clk),
    .D(_00546_),
    .Q(\cpuregs.regs[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17378_ (.CLK(clknet_leaf_189_clk),
    .D(_00547_),
    .Q(\cpuregs.regs[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17379_ (.CLK(clknet_leaf_14_clk),
    .D(_00548_),
    .Q(\cpuregs.regs[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17380_ (.CLK(clknet_leaf_16_clk),
    .D(_00549_),
    .Q(\cpuregs.regs[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17381_ (.CLK(clknet_leaf_187_clk),
    .D(_00550_),
    .Q(\cpuregs.regs[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17382_ (.CLK(clknet_leaf_19_clk),
    .D(_00551_),
    .Q(\cpuregs.regs[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17383_ (.CLK(clknet_leaf_180_clk),
    .D(_00552_),
    .Q(\cpuregs.regs[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17384_ (.CLK(clknet_leaf_172_clk),
    .D(_00553_),
    .Q(\cpuregs.regs[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17385_ (.CLK(clknet_leaf_183_clk),
    .D(_00554_),
    .Q(\cpuregs.regs[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17386_ (.CLK(clknet_leaf_182_clk),
    .D(_00555_),
    .Q(\cpuregs.regs[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17387_ (.CLK(clknet_leaf_130_clk),
    .D(_00556_),
    .Q(\cpuregs.regs[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17388_ (.CLK(clknet_leaf_116_clk),
    .D(_00557_),
    .Q(\cpuregs.regs[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17389_ (.CLK(clknet_leaf_153_clk),
    .D(_00558_),
    .Q(\cpuregs.regs[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17390_ (.CLK(clknet_leaf_140_clk),
    .D(_00559_),
    .Q(\cpuregs.regs[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17391_ (.CLK(clknet_leaf_146_clk),
    .D(_00560_),
    .Q(\cpuregs.regs[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17392_ (.CLK(clknet_leaf_130_clk),
    .D(_00561_),
    .Q(\cpuregs.regs[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17393_ (.CLK(clknet_leaf_141_clk),
    .D(_00562_),
    .Q(\cpuregs.regs[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17394_ (.CLK(clknet_leaf_140_clk),
    .D(_00563_),
    .Q(\cpuregs.regs[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17395_ (.CLK(clknet_leaf_153_clk),
    .D(_00564_),
    .Q(\cpuregs.regs[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17396_ (.CLK(clknet_leaf_179_clk),
    .D(_00565_),
    .Q(\cpuregs.regs[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17397_ (.CLK(clknet_leaf_101_clk),
    .D(_00566_),
    .Q(\cpuregs.regs[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17398_ (.CLK(clknet_leaf_98_clk),
    .D(_00567_),
    .Q(\cpuregs.regs[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17399_ (.CLK(clknet_leaf_121_clk),
    .D(_00568_),
    .Q(\cpuregs.regs[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17400_ (.CLK(clknet_leaf_164_clk),
    .D(_00569_),
    .Q(\cpuregs.regs[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17401_ (.CLK(clknet_leaf_161_clk),
    .D(_00570_),
    .Q(\cpuregs.regs[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17402_ (.CLK(clknet_leaf_111_clk),
    .D(_00571_),
    .Q(\cpuregs.regs[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17403_ (.CLK(clknet_leaf_166_clk),
    .D(_00572_),
    .Q(\cpuregs.regs[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17404_ (.CLK(clknet_leaf_100_clk),
    .D(_00573_),
    .Q(\cpuregs.regs[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17405_ (.CLK(clknet_leaf_119_clk),
    .D(_00574_),
    .Q(\cpuregs.regs[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17406_ (.CLK(clknet_leaf_128_clk),
    .D(_00575_),
    .Q(\cpuregs.regs[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17407_ (.CLK(clknet_leaf_163_clk),
    .D(_00576_),
    .Q(\cpuregs.regs[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17408_ (.CLK(clknet_leaf_169_clk),
    .D(_00577_),
    .Q(\cpuregs.regs[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17409_ (.CLK(clknet_leaf_15_clk),
    .D(_00578_),
    .Q(\cpuregs.regs[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17410_ (.CLK(clknet_leaf_188_clk),
    .D(_00579_),
    .Q(\cpuregs.regs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17411_ (.CLK(clknet_leaf_11_clk),
    .D(_00580_),
    .Q(\cpuregs.regs[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17412_ (.CLK(clknet_leaf_7_clk),
    .D(_00581_),
    .Q(\cpuregs.regs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17413_ (.CLK(clknet_leaf_1_clk),
    .D(_00582_),
    .Q(\cpuregs.regs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17414_ (.CLK(clknet_leaf_18_clk),
    .D(_00583_),
    .Q(\cpuregs.regs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17415_ (.CLK(clknet_leaf_178_clk),
    .D(_00584_),
    .Q(\cpuregs.regs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17416_ (.CLK(clknet_leaf_173_clk),
    .D(_00585_),
    .Q(\cpuregs.regs[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17417_ (.CLK(clknet_leaf_186_clk),
    .D(_00586_),
    .Q(\cpuregs.regs[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17418_ (.CLK(clknet_leaf_185_clk),
    .D(_00587_),
    .Q(\cpuregs.regs[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17419_ (.CLK(clknet_leaf_127_clk),
    .D(_00588_),
    .Q(\cpuregs.regs[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17420_ (.CLK(clknet_leaf_162_clk),
    .D(_00589_),
    .Q(\cpuregs.regs[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17421_ (.CLK(clknet_leaf_149_clk),
    .D(_00590_),
    .Q(\cpuregs.regs[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17422_ (.CLK(clknet_leaf_137_clk),
    .D(_00591_),
    .Q(\cpuregs.regs[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17423_ (.CLK(clknet_leaf_145_clk),
    .D(_00592_),
    .Q(\cpuregs.regs[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17424_ (.CLK(clknet_leaf_159_clk),
    .D(_00593_),
    .Q(\cpuregs.regs[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17425_ (.CLK(clknet_leaf_136_clk),
    .D(_00594_),
    .Q(\cpuregs.regs[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17426_ (.CLK(clknet_leaf_140_clk),
    .D(_00595_),
    .Q(\cpuregs.regs[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17427_ (.CLK(clknet_leaf_178_clk),
    .D(_00596_),
    .Q(\cpuregs.regs[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17428_ (.CLK(clknet_leaf_179_clk),
    .D(_00597_),
    .Q(\cpuregs.regs[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17429_ (.CLK(clknet_leaf_106_clk),
    .D(_00598_),
    .Q(\cpuregs.regs[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17430_ (.CLK(clknet_leaf_97_clk),
    .D(_00599_),
    .Q(\cpuregs.regs[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17431_ (.CLK(clknet_leaf_118_clk),
    .D(_00600_),
    .Q(\cpuregs.regs[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17432_ (.CLK(clknet_leaf_165_clk),
    .D(_00601_),
    .Q(\cpuregs.regs[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17433_ (.CLK(clknet_leaf_114_clk),
    .D(_00602_),
    .Q(\cpuregs.regs[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17434_ (.CLK(clknet_leaf_112_clk),
    .D(_00603_),
    .Q(\cpuregs.regs[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17435_ (.CLK(clknet_leaf_166_clk),
    .D(_00604_),
    .Q(\cpuregs.regs[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17436_ (.CLK(clknet_leaf_106_clk),
    .D(_00605_),
    .Q(\cpuregs.regs[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17437_ (.CLK(clknet_leaf_114_clk),
    .D(_00606_),
    .Q(\cpuregs.regs[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17438_ (.CLK(clknet_leaf_125_clk),
    .D(_00607_),
    .Q(\cpuregs.regs[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17439_ (.CLK(clknet_leaf_169_clk),
    .D(_00608_),
    .Q(\cpuregs.regs[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17440_ (.CLK(clknet_leaf_170_clk),
    .D(_00609_),
    .Q(\cpuregs.regs[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17441_ (.CLK(clknet_leaf_15_clk),
    .D(_00610_),
    .Q(\cpuregs.regs[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17442_ (.CLK(clknet_leaf_188_clk),
    .D(_00611_),
    .Q(\cpuregs.regs[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17443_ (.CLK(clknet_leaf_14_clk),
    .D(_00612_),
    .Q(\cpuregs.regs[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17444_ (.CLK(clknet_leaf_12_clk),
    .D(_00613_),
    .Q(\cpuregs.regs[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17445_ (.CLK(clknet_leaf_2_clk),
    .D(_00614_),
    .Q(\cpuregs.regs[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17446_ (.CLK(clknet_leaf_167_clk),
    .D(_00615_),
    .Q(\cpuregs.regs[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17447_ (.CLK(clknet_leaf_181_clk),
    .D(_00616_),
    .Q(\cpuregs.regs[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17448_ (.CLK(clknet_leaf_175_clk),
    .D(_00617_),
    .Q(\cpuregs.regs[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17449_ (.CLK(clknet_leaf_184_clk),
    .D(_00618_),
    .Q(\cpuregs.regs[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17450_ (.CLK(clknet_leaf_183_clk),
    .D(_00619_),
    .Q(\cpuregs.regs[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17451_ (.CLK(clknet_leaf_131_clk),
    .D(_00620_),
    .Q(\cpuregs.regs[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17452_ (.CLK(clknet_leaf_159_clk),
    .D(_00621_),
    .Q(\cpuregs.regs[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17453_ (.CLK(clknet_leaf_148_clk),
    .D(_00622_),
    .Q(\cpuregs.regs[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17454_ (.CLK(clknet_leaf_137_clk),
    .D(_00623_),
    .Q(\cpuregs.regs[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17455_ (.CLK(clknet_leaf_144_clk),
    .D(_00624_),
    .Q(\cpuregs.regs[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17456_ (.CLK(clknet_leaf_133_clk),
    .D(_00625_),
    .Q(\cpuregs.regs[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17457_ (.CLK(clknet_leaf_132_clk),
    .D(_00626_),
    .Q(\cpuregs.regs[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17458_ (.CLK(clknet_leaf_147_clk),
    .D(_00627_),
    .Q(\cpuregs.regs[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17459_ (.CLK(clknet_leaf_151_clk),
    .D(_00628_),
    .Q(\cpuregs.regs[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17460_ (.CLK(clknet_leaf_151_clk),
    .D(_00629_),
    .Q(\cpuregs.regs[31][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17461_ (.CLK(clknet_leaf_98_clk),
    .D(_00630_),
    .Q(\cpuregs.regs[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17462_ (.CLK(clknet_leaf_97_clk),
    .D(_00631_),
    .Q(\cpuregs.regs[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17463_ (.CLK(clknet_leaf_122_clk),
    .D(_00632_),
    .Q(\cpuregs.regs[31][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17464_ (.CLK(clknet_leaf_164_clk),
    .D(_00633_),
    .Q(\cpuregs.regs[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17465_ (.CLK(clknet_leaf_160_clk),
    .D(_00634_),
    .Q(\cpuregs.regs[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17466_ (.CLK(clknet_leaf_112_clk),
    .D(_00635_),
    .Q(\cpuregs.regs[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17467_ (.CLK(clknet_leaf_109_clk),
    .D(_00636_),
    .Q(\cpuregs.regs[31][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17468_ (.CLK(clknet_leaf_112_clk),
    .D(_00637_),
    .Q(\cpuregs.regs[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17469_ (.CLK(clknet_leaf_114_clk),
    .D(_00638_),
    .Q(\cpuregs.regs[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17470_ (.CLK(clknet_leaf_128_clk),
    .D(_00639_),
    .Q(\cpuregs.regs[31][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17471_ (.CLK(clknet_leaf_177_clk),
    .D(_00640_),
    .Q(\cpuregs.regs[31][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17472_ (.CLK(clknet_leaf_176_clk),
    .D(_00641_),
    .Q(\cpuregs.regs[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17473_ (.CLK(clknet_leaf_17_clk),
    .D(_00642_),
    .Q(\cpuregs.regs[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17474_ (.CLK(clknet_leaf_1_clk),
    .D(_00643_),
    .Q(\cpuregs.regs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17475_ (.CLK(clknet_leaf_16_clk),
    .D(_00644_),
    .Q(\cpuregs.regs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17476_ (.CLK(clknet_leaf_7_clk),
    .D(_00645_),
    .Q(\cpuregs.regs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17477_ (.CLK(clknet_leaf_2_clk),
    .D(_00646_),
    .Q(\cpuregs.regs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17478_ (.CLK(clknet_leaf_17_clk),
    .D(_00647_),
    .Q(\cpuregs.regs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17479_ (.CLK(clknet_leaf_178_clk),
    .D(_00648_),
    .Q(\cpuregs.regs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17480_ (.CLK(clknet_leaf_13_clk),
    .D(_00649_),
    .Q(\cpuregs.regs[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17481_ (.CLK(clknet_leaf_186_clk),
    .D(_00650_),
    .Q(\cpuregs.regs[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17482_ (.CLK(clknet_leaf_175_clk),
    .D(_00651_),
    .Q(\cpuregs.regs[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17483_ (.CLK(clknet_leaf_126_clk),
    .D(_00652_),
    .Q(\cpuregs.regs[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17484_ (.CLK(clknet_leaf_160_clk),
    .D(_00653_),
    .Q(\cpuregs.regs[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17485_ (.CLK(clknet_leaf_153_clk),
    .D(_00654_),
    .Q(\cpuregs.regs[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17486_ (.CLK(clknet_leaf_136_clk),
    .D(_00655_),
    .Q(\cpuregs.regs[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17487_ (.CLK(clknet_leaf_144_clk),
    .D(_00656_),
    .Q(\cpuregs.regs[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17488_ (.CLK(clknet_leaf_116_clk),
    .D(_00657_),
    .Q(\cpuregs.regs[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17489_ (.CLK(clknet_leaf_134_clk),
    .D(_00658_),
    .Q(\cpuregs.regs[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17490_ (.CLK(clknet_leaf_142_clk),
    .D(_00659_),
    .Q(\cpuregs.regs[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17491_ (.CLK(clknet_leaf_156_clk),
    .D(_00660_),
    .Q(\cpuregs.regs[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17492_ (.CLK(clknet_leaf_152_clk),
    .D(_00661_),
    .Q(\cpuregs.regs[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17493_ (.CLK(clknet_leaf_100_clk),
    .D(_00662_),
    .Q(\cpuregs.regs[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17494_ (.CLK(clknet_leaf_98_clk),
    .D(_00663_),
    .Q(\cpuregs.regs[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17495_ (.CLK(clknet_leaf_119_clk),
    .D(_00664_),
    .Q(\cpuregs.regs[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17496_ (.CLK(clknet_leaf_165_clk),
    .D(_00665_),
    .Q(\cpuregs.regs[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17497_ (.CLK(clknet_leaf_114_clk),
    .D(_00666_),
    .Q(\cpuregs.regs[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17498_ (.CLK(clknet_leaf_109_clk),
    .D(_00667_),
    .Q(\cpuregs.regs[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17499_ (.CLK(clknet_leaf_20_clk),
    .D(_00668_),
    .Q(\cpuregs.regs[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17500_ (.CLK(clknet_leaf_105_clk),
    .D(_00669_),
    .Q(\cpuregs.regs[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17501_ (.CLK(clknet_leaf_119_clk),
    .D(_00670_),
    .Q(\cpuregs.regs[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17502_ (.CLK(clknet_leaf_118_clk),
    .D(_00671_),
    .Q(\cpuregs.regs[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17503_ (.CLK(clknet_leaf_162_clk),
    .D(_00672_),
    .Q(\cpuregs.regs[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17504_ (.CLK(clknet_leaf_170_clk),
    .D(_00673_),
    .Q(\cpuregs.regs[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17505_ (.CLK(clknet_leaf_15_clk),
    .D(_00674_),
    .Q(\cpuregs.regs[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17506_ (.CLK(clknet_leaf_188_clk),
    .D(_00675_),
    .Q(\cpuregs.regs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17507_ (.CLK(clknet_leaf_11_clk),
    .D(_00676_),
    .Q(\cpuregs.regs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17508_ (.CLK(clknet_leaf_7_clk),
    .D(_00677_),
    .Q(\cpuregs.regs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17509_ (.CLK(clknet_leaf_1_clk),
    .D(_00678_),
    .Q(\cpuregs.regs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17510_ (.CLK(clknet_leaf_18_clk),
    .D(_00679_),
    .Q(\cpuregs.regs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17511_ (.CLK(clknet_leaf_178_clk),
    .D(_00680_),
    .Q(\cpuregs.regs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17512_ (.CLK(clknet_leaf_173_clk),
    .D(_00681_),
    .Q(\cpuregs.regs[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17513_ (.CLK(clknet_leaf_186_clk),
    .D(_00682_),
    .Q(\cpuregs.regs[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17514_ (.CLK(clknet_leaf_175_clk),
    .D(_00683_),
    .Q(\cpuregs.regs[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17515_ (.CLK(clknet_leaf_127_clk),
    .D(_00684_),
    .Q(\cpuregs.regs[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17516_ (.CLK(clknet_leaf_162_clk),
    .D(_00685_),
    .Q(\cpuregs.regs[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17517_ (.CLK(clknet_leaf_148_clk),
    .D(_00686_),
    .Q(\cpuregs.regs[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17518_ (.CLK(clknet_leaf_137_clk),
    .D(_00687_),
    .Q(\cpuregs.regs[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17519_ (.CLK(clknet_leaf_145_clk),
    .D(_00688_),
    .Q(\cpuregs.regs[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17520_ (.CLK(clknet_leaf_130_clk),
    .D(_00689_),
    .Q(\cpuregs.regs[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17521_ (.CLK(clknet_leaf_136_clk),
    .D(_00690_),
    .Q(\cpuregs.regs[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17522_ (.CLK(clknet_leaf_146_clk),
    .D(_00691_),
    .Q(\cpuregs.regs[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17523_ (.CLK(clknet_leaf_154_clk),
    .D(_00692_),
    .Q(\cpuregs.regs[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17524_ (.CLK(clknet_leaf_152_clk),
    .D(_00693_),
    .Q(\cpuregs.regs[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17525_ (.CLK(clknet_leaf_105_clk),
    .D(_00694_),
    .Q(\cpuregs.regs[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17526_ (.CLK(clknet_leaf_97_clk),
    .D(_00695_),
    .Q(\cpuregs.regs[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17527_ (.CLK(clknet_leaf_117_clk),
    .D(_00696_),
    .Q(\cpuregs.regs[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17528_ (.CLK(clknet_leaf_165_clk),
    .D(_00697_),
    .Q(\cpuregs.regs[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17529_ (.CLK(clknet_leaf_114_clk),
    .D(_00698_),
    .Q(\cpuregs.regs[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17530_ (.CLK(clknet_leaf_106_clk),
    .D(_00699_),
    .Q(\cpuregs.regs[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17531_ (.CLK(clknet_leaf_166_clk),
    .D(_00700_),
    .Q(\cpuregs.regs[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17532_ (.CLK(clknet_leaf_107_clk),
    .D(_00701_),
    .Q(\cpuregs.regs[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17533_ (.CLK(clknet_leaf_114_clk),
    .D(_00702_),
    .Q(\cpuregs.regs[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17534_ (.CLK(clknet_leaf_125_clk),
    .D(_00703_),
    .Q(\cpuregs.regs[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17535_ (.CLK(clknet_leaf_163_clk),
    .D(_00704_),
    .Q(\cpuregs.regs[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17536_ (.CLK(clknet_leaf_172_clk),
    .D(_00705_),
    .Q(\cpuregs.regs[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17537_ (.CLK(clknet_leaf_15_clk),
    .D(_00706_),
    .Q(\cpuregs.regs[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17538_ (.CLK(clknet_leaf_188_clk),
    .D(_00707_),
    .Q(\cpuregs.regs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17539_ (.CLK(clknet_leaf_11_clk),
    .D(_00708_),
    .Q(\cpuregs.regs[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17540_ (.CLK(clknet_leaf_10_clk),
    .D(_00709_),
    .Q(\cpuregs.regs[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17541_ (.CLK(clknet_leaf_1_clk),
    .D(_00710_),
    .Q(\cpuregs.regs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17542_ (.CLK(clknet_leaf_166_clk),
    .D(_00711_),
    .Q(\cpuregs.regs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17543_ (.CLK(clknet_leaf_178_clk),
    .D(_00712_),
    .Q(\cpuregs.regs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17544_ (.CLK(clknet_leaf_173_clk),
    .D(_00713_),
    .Q(\cpuregs.regs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17545_ (.CLK(clknet_leaf_185_clk),
    .D(_00714_),
    .Q(\cpuregs.regs[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17546_ (.CLK(clknet_leaf_182_clk),
    .D(_00715_),
    .Q(\cpuregs.regs[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17547_ (.CLK(clknet_leaf_127_clk),
    .D(_00716_),
    .Q(\cpuregs.regs[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17548_ (.CLK(clknet_leaf_158_clk),
    .D(_00717_),
    .Q(\cpuregs.regs[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17549_ (.CLK(clknet_leaf_145_clk),
    .D(_00718_),
    .Q(\cpuregs.regs[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17550_ (.CLK(clknet_leaf_136_clk),
    .D(_00719_),
    .Q(\cpuregs.regs[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17551_ (.CLK(clknet_leaf_145_clk),
    .D(_00720_),
    .Q(\cpuregs.regs[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17552_ (.CLK(clknet_leaf_130_clk),
    .D(_00721_),
    .Q(\cpuregs.regs[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17553_ (.CLK(clknet_leaf_136_clk),
    .D(_00722_),
    .Q(\cpuregs.regs[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17554_ (.CLK(clknet_leaf_140_clk),
    .D(_00723_),
    .Q(\cpuregs.regs[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17555_ (.CLK(clknet_leaf_154_clk),
    .D(_00724_),
    .Q(\cpuregs.regs[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17556_ (.CLK(clknet_leaf_152_clk),
    .D(_00725_),
    .Q(\cpuregs.regs[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17557_ (.CLK(clknet_leaf_100_clk),
    .D(_00726_),
    .Q(\cpuregs.regs[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17558_ (.CLK(clknet_leaf_97_clk),
    .D(_00727_),
    .Q(\cpuregs.regs[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17559_ (.CLK(clknet_leaf_118_clk),
    .D(_00728_),
    .Q(\cpuregs.regs[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17560_ (.CLK(clknet_leaf_109_clk),
    .D(_00729_),
    .Q(\cpuregs.regs[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17561_ (.CLK(clknet_leaf_114_clk),
    .D(_00730_),
    .Q(\cpuregs.regs[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17562_ (.CLK(clknet_leaf_106_clk),
    .D(_00731_),
    .Q(\cpuregs.regs[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17563_ (.CLK(clknet_leaf_165_clk),
    .D(_00732_),
    .Q(\cpuregs.regs[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17564_ (.CLK(clknet_leaf_105_clk),
    .D(_00733_),
    .Q(\cpuregs.regs[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17565_ (.CLK(clknet_leaf_113_clk),
    .D(_00734_),
    .Q(\cpuregs.regs[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17566_ (.CLK(clknet_leaf_125_clk),
    .D(_00735_),
    .Q(\cpuregs.regs[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17567_ (.CLK(clknet_leaf_162_clk),
    .D(_00736_),
    .Q(\cpuregs.regs[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17568_ (.CLK(clknet_leaf_170_clk),
    .D(_00737_),
    .Q(\cpuregs.regs[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17569_ (.CLK(clknet_leaf_17_clk),
    .D(_00738_),
    .Q(\cpuregs.regs[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17570_ (.CLK(clknet_leaf_189_clk),
    .D(_00739_),
    .Q(\cpuregs.regs[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17571_ (.CLK(clknet_leaf_15_clk),
    .D(_00740_),
    .Q(\cpuregs.regs[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17572_ (.CLK(clknet_leaf_16_clk),
    .D(_00741_),
    .Q(\cpuregs.regs[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17573_ (.CLK(clknet_leaf_187_clk),
    .D(_00742_),
    .Q(\cpuregs.regs[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17574_ (.CLK(clknet_leaf_19_clk),
    .D(_00743_),
    .Q(\cpuregs.regs[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17575_ (.CLK(clknet_leaf_180_clk),
    .D(_00744_),
    .Q(\cpuregs.regs[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17576_ (.CLK(clknet_leaf_172_clk),
    .D(_00745_),
    .Q(\cpuregs.regs[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17577_ (.CLK(clknet_leaf_183_clk),
    .D(_00746_),
    .Q(\cpuregs.regs[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17578_ (.CLK(clknet_leaf_182_clk),
    .D(_00747_),
    .Q(\cpuregs.regs[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17579_ (.CLK(clknet_leaf_131_clk),
    .D(_00748_),
    .Q(\cpuregs.regs[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17580_ (.CLK(clknet_leaf_115_clk),
    .D(_00749_),
    .Q(\cpuregs.regs[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17581_ (.CLK(clknet_leaf_149_clk),
    .D(_00750_),
    .Q(\cpuregs.regs[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17582_ (.CLK(clknet_leaf_138_clk),
    .D(_00751_),
    .Q(\cpuregs.regs[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17583_ (.CLK(clknet_leaf_146_clk),
    .D(_00752_),
    .Q(\cpuregs.regs[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17584_ (.CLK(clknet_leaf_129_clk),
    .D(_00753_),
    .Q(\cpuregs.regs[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17585_ (.CLK(clknet_leaf_131_clk),
    .D(_00754_),
    .Q(\cpuregs.regs[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17586_ (.CLK(clknet_leaf_141_clk),
    .D(_00755_),
    .Q(\cpuregs.regs[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17587_ (.CLK(clknet_leaf_153_clk),
    .D(_00756_),
    .Q(\cpuregs.regs[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17588_ (.CLK(clknet_leaf_152_clk),
    .D(_00757_),
    .Q(\cpuregs.regs[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17589_ (.CLK(clknet_leaf_98_clk),
    .D(_00758_),
    .Q(\cpuregs.regs[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17590_ (.CLK(clknet_leaf_98_clk),
    .D(_00759_),
    .Q(\cpuregs.regs[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17591_ (.CLK(clknet_leaf_121_clk),
    .D(_00760_),
    .Q(\cpuregs.regs[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17592_ (.CLK(clknet_leaf_161_clk),
    .D(_00761_),
    .Q(\cpuregs.regs[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17593_ (.CLK(clknet_leaf_161_clk),
    .D(_00762_),
    .Q(\cpuregs.regs[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17594_ (.CLK(clknet_leaf_111_clk),
    .D(_00763_),
    .Q(\cpuregs.regs[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17595_ (.CLK(clknet_leaf_166_clk),
    .D(_00764_),
    .Q(\cpuregs.regs[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17596_ (.CLK(clknet_leaf_105_clk),
    .D(_00765_),
    .Q(\cpuregs.regs[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17597_ (.CLK(clknet_leaf_119_clk),
    .D(_00766_),
    .Q(\cpuregs.regs[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17598_ (.CLK(clknet_leaf_129_clk),
    .D(_00767_),
    .Q(\cpuregs.regs[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17599_ (.CLK(clknet_leaf_163_clk),
    .D(_00768_),
    .Q(\cpuregs.regs[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17600_ (.CLK(clknet_leaf_169_clk),
    .D(_00769_),
    .Q(\cpuregs.regs[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17601_ (.CLK(clknet_leaf_16_clk),
    .D(_00770_),
    .Q(\cpuregs.regs[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17602_ (.CLK(clknet_leaf_188_clk),
    .D(_00771_),
    .Q(\cpuregs.regs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17603_ (.CLK(clknet_leaf_7_clk),
    .D(_00772_),
    .Q(\cpuregs.regs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17604_ (.CLK(clknet_leaf_7_clk),
    .D(_00773_),
    .Q(\cpuregs.regs[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17605_ (.CLK(clknet_leaf_2_clk),
    .D(_00774_),
    .Q(\cpuregs.regs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17606_ (.CLK(clknet_leaf_18_clk),
    .D(_00775_),
    .Q(\cpuregs.regs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17607_ (.CLK(clknet_leaf_178_clk),
    .D(_00776_),
    .Q(\cpuregs.regs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17608_ (.CLK(clknet_leaf_173_clk),
    .D(_00777_),
    .Q(\cpuregs.regs[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17609_ (.CLK(clknet_leaf_186_clk),
    .D(_00778_),
    .Q(\cpuregs.regs[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17610_ (.CLK(clknet_leaf_175_clk),
    .D(_00779_),
    .Q(\cpuregs.regs[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17611_ (.CLK(clknet_leaf_127_clk),
    .D(_00780_),
    .Q(\cpuregs.regs[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17612_ (.CLK(clknet_leaf_160_clk),
    .D(_00781_),
    .Q(\cpuregs.regs[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17613_ (.CLK(clknet_leaf_145_clk),
    .D(_00782_),
    .Q(\cpuregs.regs[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17614_ (.CLK(clknet_leaf_136_clk),
    .D(_00783_),
    .Q(\cpuregs.regs[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17615_ (.CLK(clknet_leaf_145_clk),
    .D(_00784_),
    .Q(\cpuregs.regs[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17616_ (.CLK(clknet_leaf_130_clk),
    .D(_00785_),
    .Q(\cpuregs.regs[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17617_ (.CLK(clknet_leaf_136_clk),
    .D(_00786_),
    .Q(\cpuregs.regs[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17618_ (.CLK(clknet_leaf_140_clk),
    .D(_00787_),
    .Q(\cpuregs.regs[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17619_ (.CLK(clknet_leaf_154_clk),
    .D(_00788_),
    .Q(\cpuregs.regs[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17620_ (.CLK(clknet_leaf_152_clk),
    .D(_00789_),
    .Q(\cpuregs.regs[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17621_ (.CLK(clknet_leaf_100_clk),
    .D(_00790_),
    .Q(\cpuregs.regs[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17622_ (.CLK(clknet_leaf_97_clk),
    .D(_00791_),
    .Q(\cpuregs.regs[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17623_ (.CLK(clknet_leaf_118_clk),
    .D(_00792_),
    .Q(\cpuregs.regs[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17624_ (.CLK(clknet_leaf_109_clk),
    .D(_00793_),
    .Q(\cpuregs.regs[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17625_ (.CLK(clknet_leaf_114_clk),
    .D(_00794_),
    .Q(\cpuregs.regs[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17626_ (.CLK(clknet_leaf_106_clk),
    .D(_00795_),
    .Q(\cpuregs.regs[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17627_ (.CLK(clknet_leaf_166_clk),
    .D(_00796_),
    .Q(\cpuregs.regs[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17628_ (.CLK(clknet_leaf_106_clk),
    .D(_00797_),
    .Q(\cpuregs.regs[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17629_ (.CLK(clknet_leaf_113_clk),
    .D(_00798_),
    .Q(\cpuregs.regs[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17630_ (.CLK(clknet_leaf_124_clk),
    .D(_00799_),
    .Q(\cpuregs.regs[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17631_ (.CLK(clknet_leaf_163_clk),
    .D(_00800_),
    .Q(\cpuregs.regs[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17632_ (.CLK(clknet_leaf_172_clk),
    .D(_00801_),
    .Q(\cpuregs.regs[5][31] ));
 sky130_fd_sc_hd__dfxtp_4 _17633_ (.CLK(clknet_leaf_50_clk),
    .D(_00802_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_4 _17634_ (.CLK(clknet_leaf_52_clk),
    .D(_00803_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_4 _17635_ (.CLK(clknet_leaf_51_clk),
    .D(_00804_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_4 _17636_ (.CLK(clknet_leaf_51_clk),
    .D(_00805_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_4 _17637_ (.CLK(clknet_leaf_50_clk),
    .D(_00806_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_2 _17638_ (.CLK(clknet_leaf_51_clk),
    .D(_00807_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_4 _17639_ (.CLK(clknet_leaf_51_clk),
    .D(_00808_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_2 _17640_ (.CLK(clknet_leaf_51_clk),
    .D(_00809_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _17641_ (.CLK(clknet_leaf_46_clk),
    .D(_00810_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_4 _17642_ (.CLK(clknet_leaf_46_clk),
    .D(_00811_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_4 _17643_ (.CLK(clknet_leaf_47_clk),
    .D(_00812_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_4 _17644_ (.CLK(clknet_leaf_47_clk),
    .D(_00813_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_4 _17645_ (.CLK(clknet_leaf_47_clk),
    .D(_00814_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_4 _17646_ (.CLK(clknet_leaf_47_clk),
    .D(_00815_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_4 _17647_ (.CLK(clknet_leaf_47_clk),
    .D(_00816_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_4 _17648_ (.CLK(clknet_leaf_49_clk),
    .D(_00817_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_4 _17649_ (.CLK(clknet_leaf_47_clk),
    .D(_00818_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_2 _17650_ (.CLK(clknet_leaf_47_clk),
    .D(_00819_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_2 _17651_ (.CLK(clknet_leaf_49_clk),
    .D(_00820_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_2 _17652_ (.CLK(clknet_leaf_49_clk),
    .D(_00821_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_2 _17653_ (.CLK(clknet_leaf_48_clk),
    .D(_00822_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_2 _17654_ (.CLK(clknet_leaf_47_clk),
    .D(_00823_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_4 _17655_ (.CLK(clknet_leaf_72_clk),
    .D(_00824_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_2 _17656_ (.CLK(clknet_leaf_48_clk),
    .D(_00825_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_2 _17657_ (.CLK(clknet_leaf_71_clk),
    .D(_00826_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_2 _17658_ (.CLK(clknet_leaf_71_clk),
    .D(_00827_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_2 _17659_ (.CLK(clknet_leaf_72_clk),
    .D(_00828_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_4 _17660_ (.CLK(clknet_leaf_49_clk),
    .D(_00829_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_4 _17661_ (.CLK(clknet_leaf_72_clk),
    .D(_00830_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_4 _17662_ (.CLK(clknet_leaf_72_clk),
    .D(_00831_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_4 _17663_ (.CLK(clknet_leaf_70_clk),
    .D(_00832_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_1 _17664_ (.CLK(clknet_leaf_17_clk),
    .D(_00833_),
    .Q(\cpuregs.regs[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17665_ (.CLK(clknet_leaf_188_clk),
    .D(_00834_),
    .Q(\cpuregs.regs[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17666_ (.CLK(clknet_leaf_16_clk),
    .D(_00835_),
    .Q(\cpuregs.regs[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17667_ (.CLK(clknet_leaf_8_clk),
    .D(_00836_),
    .Q(\cpuregs.regs[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17668_ (.CLK(clknet_leaf_2_clk),
    .D(_00837_),
    .Q(\cpuregs.regs[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17669_ (.CLK(clknet_leaf_19_clk),
    .D(_00838_),
    .Q(\cpuregs.regs[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17670_ (.CLK(clknet_leaf_177_clk),
    .D(_00839_),
    .Q(\cpuregs.regs[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17671_ (.CLK(clknet_leaf_172_clk),
    .D(_00840_),
    .Q(\cpuregs.regs[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17672_ (.CLK(clknet_leaf_185_clk),
    .D(_00841_),
    .Q(\cpuregs.regs[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17673_ (.CLK(clknet_leaf_176_clk),
    .D(_00842_),
    .Q(\cpuregs.regs[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17674_ (.CLK(clknet_leaf_126_clk),
    .D(_00843_),
    .Q(\cpuregs.regs[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17675_ (.CLK(clknet_leaf_160_clk),
    .D(_00844_),
    .Q(\cpuregs.regs[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17676_ (.CLK(clknet_leaf_150_clk),
    .D(_00845_),
    .Q(\cpuregs.regs[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17677_ (.CLK(clknet_leaf_136_clk),
    .D(_00846_),
    .Q(\cpuregs.regs[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17678_ (.CLK(clknet_leaf_144_clk),
    .D(_00847_),
    .Q(\cpuregs.regs[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17679_ (.CLK(clknet_leaf_116_clk),
    .D(_00848_),
    .Q(\cpuregs.regs[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17680_ (.CLK(clknet_leaf_134_clk),
    .D(_00849_),
    .Q(\cpuregs.regs[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17681_ (.CLK(clknet_leaf_142_clk),
    .D(_00850_),
    .Q(\cpuregs.regs[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17682_ (.CLK(clknet_leaf_156_clk),
    .D(_00851_),
    .Q(\cpuregs.regs[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17683_ (.CLK(clknet_leaf_152_clk),
    .D(_00852_),
    .Q(\cpuregs.regs[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17684_ (.CLK(clknet_leaf_100_clk),
    .D(_00853_),
    .Q(\cpuregs.regs[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17685_ (.CLK(clknet_leaf_97_clk),
    .D(_00854_),
    .Q(\cpuregs.regs[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17686_ (.CLK(clknet_leaf_119_clk),
    .D(_00855_),
    .Q(\cpuregs.regs[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17687_ (.CLK(clknet_leaf_164_clk),
    .D(_00856_),
    .Q(\cpuregs.regs[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17688_ (.CLK(clknet_leaf_115_clk),
    .D(_00857_),
    .Q(\cpuregs.regs[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17689_ (.CLK(clknet_leaf_108_clk),
    .D(_00858_),
    .Q(\cpuregs.regs[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17690_ (.CLK(clknet_leaf_20_clk),
    .D(_00859_),
    .Q(\cpuregs.regs[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17691_ (.CLK(clknet_leaf_105_clk),
    .D(_00860_),
    .Q(\cpuregs.regs[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17692_ (.CLK(clknet_leaf_119_clk),
    .D(_00861_),
    .Q(\cpuregs.regs[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17693_ (.CLK(clknet_leaf_125_clk),
    .D(_00862_),
    .Q(\cpuregs.regs[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17694_ (.CLK(clknet_leaf_162_clk),
    .D(_00863_),
    .Q(\cpuregs.regs[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17695_ (.CLK(clknet_leaf_169_clk),
    .D(_00864_),
    .Q(\cpuregs.regs[0][31] ));
 sky130_fd_sc_hd__dfxtp_2 _17696_ (.CLK(clknet_leaf_39_clk),
    .D(_00865_),
    .Q(net299));
 sky130_fd_sc_hd__dfxtp_1 _17697_ (.CLK(clknet_leaf_75_clk),
    .D(_00866_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_1 _17698_ (.CLK(clknet_leaf_75_clk),
    .D(_00867_),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_1 _17699_ (.CLK(clknet_leaf_75_clk),
    .D(_00868_),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_1 _17700_ (.CLK(clknet_leaf_75_clk),
    .D(_00869_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 _17701_ (.CLK(clknet_leaf_75_clk),
    .D(_00870_),
    .Q(net157));
 sky130_fd_sc_hd__dfxtp_1 _17702_ (.CLK(clknet_leaf_75_clk),
    .D(_00871_),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_1 _17703_ (.CLK(clknet_leaf_75_clk),
    .D(_00872_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_1 _17704_ (.CLK(clknet_leaf_75_clk),
    .D(_00873_),
    .Q(net160));
 sky130_fd_sc_hd__dfxtp_1 _17705_ (.CLK(clknet_leaf_75_clk),
    .D(_00874_),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_1 _17706_ (.CLK(clknet_leaf_75_clk),
    .D(_00875_),
    .Q(net162));
 sky130_fd_sc_hd__dfxtp_1 _17707_ (.CLK(clknet_leaf_75_clk),
    .D(_00876_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_1 _17708_ (.CLK(clknet_leaf_76_clk),
    .D(_00877_),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_1 _17709_ (.CLK(clknet_leaf_75_clk),
    .D(_00878_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_1 _17710_ (.CLK(clknet_leaf_75_clk),
    .D(_00879_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_1 _17711_ (.CLK(clknet_leaf_76_clk),
    .D(_00880_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_1 _17712_ (.CLK(clknet_leaf_83_clk),
    .D(_00881_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_1 _17713_ (.CLK(clknet_leaf_76_clk),
    .D(_00882_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 _17714_ (.CLK(clknet_leaf_76_clk),
    .D(_00883_),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_1 _17715_ (.CLK(clknet_leaf_76_clk),
    .D(_00884_),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_1 _17716_ (.CLK(clknet_leaf_76_clk),
    .D(_00885_),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_1 _17717_ (.CLK(clknet_leaf_76_clk),
    .D(_00886_),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_1 _17718_ (.CLK(clknet_leaf_76_clk),
    .D(_00887_),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_1 _17719_ (.CLK(clknet_leaf_83_clk),
    .D(_00888_),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_1 _17720_ (.CLK(clknet_leaf_77_clk),
    .D(_00889_),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_1 _17721_ (.CLK(clknet_leaf_83_clk),
    .D(_00890_),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_1 _17722_ (.CLK(clknet_leaf_77_clk),
    .D(_00891_),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_1 _17723_ (.CLK(clknet_leaf_76_clk),
    .D(_00892_),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_1 _17724_ (.CLK(clknet_leaf_82_clk),
    .D(_00893_),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_1 _17725_ (.CLK(clknet_leaf_83_clk),
    .D(_00894_),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_1 _17726_ (.CLK(clknet_leaf_82_clk),
    .D(_00895_),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_1 _17727_ (.CLK(clknet_leaf_74_clk),
    .D(_00896_),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_1 _17728_ (.CLK(clknet_leaf_74_clk),
    .D(_00897_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 _17729_ (.CLK(clknet_leaf_101_clk),
    .D(_00898_),
    .Q(\count_instr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _17730_ (.CLK(clknet_leaf_101_clk),
    .D(_00899_),
    .Q(\count_instr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _17731_ (.CLK(clknet_leaf_101_clk),
    .D(_00900_),
    .Q(\count_instr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _17732_ (.CLK(clknet_leaf_101_clk),
    .D(_00901_),
    .Q(\count_instr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _17733_ (.CLK(clknet_leaf_93_clk),
    .D(_00902_),
    .Q(\count_instr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _17734_ (.CLK(clknet_leaf_96_clk),
    .D(_00903_),
    .Q(\count_instr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _17735_ (.CLK(clknet_leaf_96_clk),
    .D(_00904_),
    .Q(\count_instr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _17736_ (.CLK(clknet_leaf_96_clk),
    .D(_00905_),
    .Q(\count_instr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _17737_ (.CLK(clknet_leaf_96_clk),
    .D(_00906_),
    .Q(\count_instr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _17738_ (.CLK(clknet_leaf_96_clk),
    .D(_00907_),
    .Q(\count_instr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _17739_ (.CLK(clknet_leaf_96_clk),
    .D(_00908_),
    .Q(\count_instr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _17740_ (.CLK(clknet_leaf_95_clk),
    .D(_00909_),
    .Q(\count_instr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _17741_ (.CLK(clknet_leaf_94_clk),
    .D(_00910_),
    .Q(\count_instr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _17742_ (.CLK(clknet_leaf_95_clk),
    .D(_00911_),
    .Q(\count_instr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _17743_ (.CLK(clknet_leaf_94_clk),
    .D(_00912_),
    .Q(\count_instr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _17744_ (.CLK(clknet_leaf_87_clk),
    .D(_00913_),
    .Q(\count_instr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _17745_ (.CLK(clknet_leaf_87_clk),
    .D(_00914_),
    .Q(\count_instr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _17746_ (.CLK(clknet_leaf_86_clk),
    .D(_00915_),
    .Q(\count_instr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _17747_ (.CLK(clknet_leaf_86_clk),
    .D(_00916_),
    .Q(\count_instr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _17748_ (.CLK(clknet_leaf_86_clk),
    .D(_00917_),
    .Q(\count_instr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _17749_ (.CLK(clknet_leaf_86_clk),
    .D(_00918_),
    .Q(\count_instr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _17750_ (.CLK(clknet_leaf_86_clk),
    .D(_00919_),
    .Q(\count_instr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _17751_ (.CLK(clknet_leaf_85_clk),
    .D(_00920_),
    .Q(\count_instr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _17752_ (.CLK(clknet_leaf_85_clk),
    .D(_00921_),
    .Q(\count_instr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _17753_ (.CLK(clknet_leaf_85_clk),
    .D(_00922_),
    .Q(\count_instr[24] ));
 sky130_fd_sc_hd__dfxtp_1 _17754_ (.CLK(clknet_leaf_85_clk),
    .D(_00923_),
    .Q(\count_instr[25] ));
 sky130_fd_sc_hd__dfxtp_1 _17755_ (.CLK(clknet_leaf_89_clk),
    .D(_00924_),
    .Q(\count_instr[26] ));
 sky130_fd_sc_hd__dfxtp_1 _17756_ (.CLK(clknet_leaf_82_clk),
    .D(_00925_),
    .Q(\count_instr[27] ));
 sky130_fd_sc_hd__dfxtp_1 _17757_ (.CLK(clknet_leaf_82_clk),
    .D(_00926_),
    .Q(\count_instr[28] ));
 sky130_fd_sc_hd__dfxtp_1 _17758_ (.CLK(clknet_leaf_89_clk),
    .D(_00927_),
    .Q(\count_instr[29] ));
 sky130_fd_sc_hd__dfxtp_1 _17759_ (.CLK(clknet_leaf_90_clk),
    .D(_00928_),
    .Q(\count_instr[30] ));
 sky130_fd_sc_hd__dfxtp_1 _17760_ (.CLK(clknet_leaf_90_clk),
    .D(_00929_),
    .Q(\count_instr[31] ));
 sky130_fd_sc_hd__dfxtp_1 _17761_ (.CLK(clknet_leaf_90_clk),
    .D(_00930_),
    .Q(\count_instr[32] ));
 sky130_fd_sc_hd__dfxtp_1 _17762_ (.CLK(clknet_leaf_90_clk),
    .D(_00931_),
    .Q(\count_instr[33] ));
 sky130_fd_sc_hd__dfxtp_1 _17763_ (.CLK(clknet_leaf_90_clk),
    .D(_00932_),
    .Q(\count_instr[34] ));
 sky130_fd_sc_hd__dfxtp_1 _17764_ (.CLK(clknet_leaf_92_clk),
    .D(_00933_),
    .Q(\count_instr[35] ));
 sky130_fd_sc_hd__dfxtp_1 _17765_ (.CLK(clknet_leaf_92_clk),
    .D(_00934_),
    .Q(\count_instr[36] ));
 sky130_fd_sc_hd__dfxtp_1 _17766_ (.CLK(clknet_leaf_94_clk),
    .D(_00935_),
    .Q(\count_instr[37] ));
 sky130_fd_sc_hd__dfxtp_1 _17767_ (.CLK(clknet_leaf_94_clk),
    .D(_00936_),
    .Q(\count_instr[38] ));
 sky130_fd_sc_hd__dfxtp_1 _17768_ (.CLK(clknet_leaf_94_clk),
    .D(_00937_),
    .Q(\count_instr[39] ));
 sky130_fd_sc_hd__dfxtp_1 _17769_ (.CLK(clknet_leaf_95_clk),
    .D(_00938_),
    .Q(\count_instr[40] ));
 sky130_fd_sc_hd__dfxtp_1 _17770_ (.CLK(clknet_leaf_95_clk),
    .D(_00939_),
    .Q(\count_instr[41] ));
 sky130_fd_sc_hd__dfxtp_1 _17771_ (.CLK(clknet_leaf_95_clk),
    .D(_00940_),
    .Q(\count_instr[42] ));
 sky130_fd_sc_hd__dfxtp_1 _17772_ (.CLK(clknet_leaf_95_clk),
    .D(_00941_),
    .Q(\count_instr[43] ));
 sky130_fd_sc_hd__dfxtp_1 _17773_ (.CLK(clknet_leaf_95_clk),
    .D(_00942_),
    .Q(\count_instr[44] ));
 sky130_fd_sc_hd__dfxtp_1 _17774_ (.CLK(clknet_leaf_95_clk),
    .D(_00943_),
    .Q(\count_instr[45] ));
 sky130_fd_sc_hd__dfxtp_1 _17775_ (.CLK(clknet_leaf_87_clk),
    .D(_00944_),
    .Q(\count_instr[46] ));
 sky130_fd_sc_hd__dfxtp_1 _17776_ (.CLK(clknet_leaf_87_clk),
    .D(_00945_),
    .Q(\count_instr[47] ));
 sky130_fd_sc_hd__dfxtp_1 _17777_ (.CLK(clknet_leaf_86_clk),
    .D(_00946_),
    .Q(\count_instr[48] ));
 sky130_fd_sc_hd__dfxtp_1 _17778_ (.CLK(clknet_leaf_86_clk),
    .D(_00947_),
    .Q(\count_instr[49] ));
 sky130_fd_sc_hd__dfxtp_1 _17779_ (.CLK(clknet_leaf_86_clk),
    .D(_00948_),
    .Q(\count_instr[50] ));
 sky130_fd_sc_hd__dfxtp_1 _17780_ (.CLK(clknet_leaf_86_clk),
    .D(_00949_),
    .Q(\count_instr[51] ));
 sky130_fd_sc_hd__dfxtp_1 _17781_ (.CLK(clknet_leaf_86_clk),
    .D(_00950_),
    .Q(\count_instr[52] ));
 sky130_fd_sc_hd__dfxtp_1 _17782_ (.CLK(clknet_leaf_85_clk),
    .D(_00951_),
    .Q(\count_instr[53] ));
 sky130_fd_sc_hd__dfxtp_1 _17783_ (.CLK(clknet_leaf_85_clk),
    .D(_00952_),
    .Q(\count_instr[54] ));
 sky130_fd_sc_hd__dfxtp_1 _17784_ (.CLK(clknet_leaf_85_clk),
    .D(_00953_),
    .Q(\count_instr[55] ));
 sky130_fd_sc_hd__dfxtp_1 _17785_ (.CLK(clknet_leaf_85_clk),
    .D(_00954_),
    .Q(\count_instr[56] ));
 sky130_fd_sc_hd__dfxtp_1 _17786_ (.CLK(clknet_leaf_84_clk),
    .D(_00955_),
    .Q(\count_instr[57] ));
 sky130_fd_sc_hd__dfxtp_1 _17787_ (.CLK(clknet_leaf_84_clk),
    .D(_00956_),
    .Q(\count_instr[58] ));
 sky130_fd_sc_hd__dfxtp_1 _17788_ (.CLK(clknet_leaf_84_clk),
    .D(_00957_),
    .Q(\count_instr[59] ));
 sky130_fd_sc_hd__dfxtp_1 _17789_ (.CLK(clknet_leaf_84_clk),
    .D(_00958_),
    .Q(\count_instr[60] ));
 sky130_fd_sc_hd__dfxtp_1 _17790_ (.CLK(clknet_leaf_84_clk),
    .D(_00959_),
    .Q(\count_instr[61] ));
 sky130_fd_sc_hd__dfxtp_1 _17791_ (.CLK(clknet_leaf_82_clk),
    .D(_00960_),
    .Q(\count_instr[62] ));
 sky130_fd_sc_hd__dfxtp_1 _17792_ (.CLK(clknet_leaf_82_clk),
    .D(_00961_),
    .Q(\count_instr[63] ));
 sky130_fd_sc_hd__dfxtp_1 _17793_ (.CLK(clknet_leaf_22_clk),
    .D(_00962_),
    .Q(\reg_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _17794_ (.CLK(clknet_leaf_22_clk),
    .D(_00963_),
    .Q(\reg_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _17795_ (.CLK(clknet_leaf_57_clk),
    .D(_00964_),
    .Q(\reg_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _17796_ (.CLK(clknet_leaf_57_clk),
    .D(_00965_),
    .Q(\reg_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _17797_ (.CLK(clknet_leaf_57_clk),
    .D(_00966_),
    .Q(\reg_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _17798_ (.CLK(clknet_leaf_56_clk),
    .D(_00967_),
    .Q(\reg_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _17799_ (.CLK(clknet_leaf_57_clk),
    .D(_00968_),
    .Q(\reg_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _17800_ (.CLK(clknet_leaf_57_clk),
    .D(_00969_),
    .Q(\reg_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _17801_ (.CLK(clknet_leaf_55_clk),
    .D(_00970_),
    .Q(\reg_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _17802_ (.CLK(clknet_leaf_55_clk),
    .D(_00971_),
    .Q(\reg_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _17803_ (.CLK(clknet_leaf_56_clk),
    .D(_00972_),
    .Q(\reg_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _17804_ (.CLK(clknet_leaf_56_clk),
    .D(_00973_),
    .Q(\reg_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _17805_ (.CLK(clknet_leaf_62_clk),
    .D(_00974_),
    .Q(\reg_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _17806_ (.CLK(clknet_leaf_62_clk),
    .D(_00975_),
    .Q(\reg_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _17807_ (.CLK(clknet_leaf_61_clk),
    .D(_00976_),
    .Q(\reg_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _17808_ (.CLK(clknet_leaf_62_clk),
    .D(_00977_),
    .Q(\reg_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _17809_ (.CLK(clknet_leaf_62_clk),
    .D(_00978_),
    .Q(\reg_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _17810_ (.CLK(clknet_leaf_61_clk),
    .D(_00979_),
    .Q(\reg_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _17811_ (.CLK(clknet_leaf_62_clk),
    .D(_00980_),
    .Q(\reg_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _17812_ (.CLK(clknet_leaf_62_clk),
    .D(_00981_),
    .Q(\reg_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _17813_ (.CLK(clknet_leaf_63_clk),
    .D(_00982_),
    .Q(\reg_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _17814_ (.CLK(clknet_leaf_63_clk),
    .D(_00983_),
    .Q(\reg_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _17815_ (.CLK(clknet_leaf_63_clk),
    .D(_00984_),
    .Q(\reg_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 _17816_ (.CLK(clknet_leaf_68_clk),
    .D(_00985_),
    .Q(\reg_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _17817_ (.CLK(clknet_leaf_64_clk),
    .D(_00986_),
    .Q(\reg_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _17818_ (.CLK(clknet_leaf_66_clk),
    .D(_00987_),
    .Q(\reg_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _17819_ (.CLK(clknet_leaf_66_clk),
    .D(_00988_),
    .Q(\reg_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _17820_ (.CLK(clknet_leaf_67_clk),
    .D(_00989_),
    .Q(\reg_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _17821_ (.CLK(clknet_leaf_67_clk),
    .D(_00990_),
    .Q(\reg_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 _17822_ (.CLK(clknet_leaf_67_clk),
    .D(_00991_),
    .Q(\reg_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _17823_ (.CLK(clknet_leaf_68_clk),
    .D(_00992_),
    .Q(\reg_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _17824_ (.CLK(clknet_leaf_22_clk),
    .D(_00993_),
    .Q(\reg_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _17825_ (.CLK(clknet_leaf_22_clk),
    .D(_00994_),
    .Q(\reg_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _17826_ (.CLK(clknet_leaf_21_clk),
    .D(_00995_),
    .Q(\reg_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _17827_ (.CLK(clknet_leaf_57_clk),
    .D(_00996_),
    .Q(\reg_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _17828_ (.CLK(clknet_leaf_57_clk),
    .D(_00997_),
    .Q(\reg_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _17829_ (.CLK(clknet_leaf_57_clk),
    .D(_00998_),
    .Q(\reg_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _17830_ (.CLK(clknet_leaf_57_clk),
    .D(_00999_),
    .Q(\reg_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _17831_ (.CLK(clknet_leaf_58_clk),
    .D(_01000_),
    .Q(\reg_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _17832_ (.CLK(clknet_leaf_57_clk),
    .D(_01001_),
    .Q(\reg_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _17833_ (.CLK(clknet_leaf_57_clk),
    .D(_01002_),
    .Q(\reg_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _17834_ (.CLK(clknet_leaf_58_clk),
    .D(_01003_),
    .Q(\reg_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _17835_ (.CLK(clknet_leaf_57_clk),
    .D(_01004_),
    .Q(\reg_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _17836_ (.CLK(clknet_leaf_59_clk),
    .D(_01005_),
    .Q(\reg_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _17837_ (.CLK(clknet_leaf_60_clk),
    .D(_01006_),
    .Q(\reg_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _17838_ (.CLK(clknet_leaf_61_clk),
    .D(_01007_),
    .Q(\reg_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _17839_ (.CLK(clknet_leaf_61_clk),
    .D(_01008_),
    .Q(\reg_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _17840_ (.CLK(clknet_leaf_61_clk),
    .D(_01009_),
    .Q(\reg_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _17841_ (.CLK(clknet_leaf_60_clk),
    .D(_01010_),
    .Q(\reg_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _17842_ (.CLK(clknet_leaf_60_clk),
    .D(_01011_),
    .Q(\reg_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _17843_ (.CLK(clknet_leaf_60_clk),
    .D(_01012_),
    .Q(\reg_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _17844_ (.CLK(clknet_leaf_108_clk),
    .D(_01013_),
    .Q(\reg_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _17845_ (.CLK(clknet_leaf_60_clk),
    .D(_01014_),
    .Q(\reg_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _17846_ (.CLK(clknet_leaf_63_clk),
    .D(_01015_),
    .Q(\reg_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _17847_ (.CLK(clknet_leaf_60_clk),
    .D(_01016_),
    .Q(\reg_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _17848_ (.CLK(clknet_leaf_64_clk),
    .D(_01017_),
    .Q(\reg_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _17849_ (.CLK(clknet_leaf_108_clk),
    .D(_01018_),
    .Q(\reg_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _17850_ (.CLK(clknet_leaf_107_clk),
    .D(_01019_),
    .Q(\reg_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _17851_ (.CLK(clknet_leaf_104_clk),
    .D(_01020_),
    .Q(\reg_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _17852_ (.CLK(clknet_leaf_104_clk),
    .D(_01021_),
    .Q(\reg_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _17853_ (.CLK(clknet_leaf_104_clk),
    .D(_01022_),
    .Q(\reg_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 _17854_ (.CLK(clknet_leaf_64_clk),
    .D(_01023_),
    .Q(\reg_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _17855_ (.CLK(clknet_leaf_102_clk),
    .D(_01024_),
    .Q(\count_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _17856_ (.CLK(clknet_leaf_101_clk),
    .D(_01025_),
    .Q(\count_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _17857_ (.CLK(clknet_leaf_101_clk),
    .D(_01026_),
    .Q(\count_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _17858_ (.CLK(clknet_leaf_93_clk),
    .D(_01027_),
    .Q(\count_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _17859_ (.CLK(clknet_leaf_93_clk),
    .D(_01028_),
    .Q(\count_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _17860_ (.CLK(clknet_leaf_93_clk),
    .D(_01029_),
    .Q(\count_cycle[5] ));
 sky130_fd_sc_hd__dfxtp_1 _17861_ (.CLK(clknet_leaf_93_clk),
    .D(_01030_),
    .Q(\count_cycle[6] ));
 sky130_fd_sc_hd__dfxtp_1 _17862_ (.CLK(clknet_leaf_93_clk),
    .D(_01031_),
    .Q(\count_cycle[7] ));
 sky130_fd_sc_hd__dfxtp_1 _17863_ (.CLK(clknet_leaf_96_clk),
    .D(_01032_),
    .Q(\count_cycle[8] ));
 sky130_fd_sc_hd__dfxtp_1 _17864_ (.CLK(clknet_leaf_96_clk),
    .D(_01033_),
    .Q(\count_cycle[9] ));
 sky130_fd_sc_hd__dfxtp_1 _17865_ (.CLK(clknet_leaf_93_clk),
    .D(_01034_),
    .Q(\count_cycle[10] ));
 sky130_fd_sc_hd__dfxtp_1 _17866_ (.CLK(clknet_leaf_94_clk),
    .D(_01035_),
    .Q(\count_cycle[11] ));
 sky130_fd_sc_hd__dfxtp_1 _17867_ (.CLK(clknet_leaf_94_clk),
    .D(_01036_),
    .Q(\count_cycle[12] ));
 sky130_fd_sc_hd__dfxtp_1 _17868_ (.CLK(clknet_leaf_94_clk),
    .D(_01037_),
    .Q(\count_cycle[13] ));
 sky130_fd_sc_hd__dfxtp_1 _17869_ (.CLK(clknet_leaf_94_clk),
    .D(_01038_),
    .Q(\count_cycle[14] ));
 sky130_fd_sc_hd__dfxtp_1 _17870_ (.CLK(clknet_leaf_88_clk),
    .D(_01039_),
    .Q(\count_cycle[15] ));
 sky130_fd_sc_hd__dfxtp_1 _17871_ (.CLK(clknet_leaf_88_clk),
    .D(_01040_),
    .Q(\count_cycle[16] ));
 sky130_fd_sc_hd__dfxtp_1 _17872_ (.CLK(clknet_leaf_90_clk),
    .D(_01041_),
    .Q(\count_cycle[17] ));
 sky130_fd_sc_hd__dfxtp_1 _17873_ (.CLK(clknet_leaf_88_clk),
    .D(_01042_),
    .Q(\count_cycle[18] ));
 sky130_fd_sc_hd__dfxtp_1 _17874_ (.CLK(clknet_leaf_88_clk),
    .D(_01043_),
    .Q(\count_cycle[19] ));
 sky130_fd_sc_hd__dfxtp_1 _17875_ (.CLK(clknet_leaf_88_clk),
    .D(_01044_),
    .Q(\count_cycle[20] ));
 sky130_fd_sc_hd__dfxtp_1 _17876_ (.CLK(clknet_leaf_88_clk),
    .D(_01045_),
    .Q(\count_cycle[21] ));
 sky130_fd_sc_hd__dfxtp_1 _17877_ (.CLK(clknet_leaf_88_clk),
    .D(_01046_),
    .Q(\count_cycle[22] ));
 sky130_fd_sc_hd__dfxtp_1 _17878_ (.CLK(clknet_leaf_85_clk),
    .D(_01047_),
    .Q(\count_cycle[23] ));
 sky130_fd_sc_hd__dfxtp_1 _17879_ (.CLK(clknet_leaf_88_clk),
    .D(_01048_),
    .Q(\count_cycle[24] ));
 sky130_fd_sc_hd__dfxtp_1 _17880_ (.CLK(clknet_leaf_88_clk),
    .D(_01049_),
    .Q(\count_cycle[25] ));
 sky130_fd_sc_hd__dfxtp_1 _17881_ (.CLK(clknet_leaf_89_clk),
    .D(_01050_),
    .Q(\count_cycle[26] ));
 sky130_fd_sc_hd__dfxtp_1 _17882_ (.CLK(clknet_leaf_89_clk),
    .D(_01051_),
    .Q(\count_cycle[27] ));
 sky130_fd_sc_hd__dfxtp_1 _17883_ (.CLK(clknet_leaf_89_clk),
    .D(_01052_),
    .Q(\count_cycle[28] ));
 sky130_fd_sc_hd__dfxtp_1 _17884_ (.CLK(clknet_leaf_81_clk),
    .D(_01053_),
    .Q(\count_cycle[29] ));
 sky130_fd_sc_hd__dfxtp_1 _17885_ (.CLK(clknet_leaf_89_clk),
    .D(_01054_),
    .Q(\count_cycle[30] ));
 sky130_fd_sc_hd__dfxtp_1 _17886_ (.CLK(clknet_leaf_90_clk),
    .D(_01055_),
    .Q(\count_cycle[31] ));
 sky130_fd_sc_hd__dfxtp_1 _17887_ (.CLK(clknet_leaf_90_clk),
    .D(_01056_),
    .Q(\count_cycle[32] ));
 sky130_fd_sc_hd__dfxtp_1 _17888_ (.CLK(clknet_leaf_90_clk),
    .D(_01057_),
    .Q(\count_cycle[33] ));
 sky130_fd_sc_hd__dfxtp_1 _17889_ (.CLK(clknet_leaf_92_clk),
    .D(_01058_),
    .Q(\count_cycle[34] ));
 sky130_fd_sc_hd__dfxtp_1 _17890_ (.CLK(clknet_leaf_92_clk),
    .D(_01059_),
    .Q(\count_cycle[35] ));
 sky130_fd_sc_hd__dfxtp_1 _17891_ (.CLK(clknet_leaf_92_clk),
    .D(_01060_),
    .Q(\count_cycle[36] ));
 sky130_fd_sc_hd__dfxtp_1 _17892_ (.CLK(clknet_leaf_92_clk),
    .D(_01061_),
    .Q(\count_cycle[37] ));
 sky130_fd_sc_hd__dfxtp_1 _17893_ (.CLK(clknet_leaf_93_clk),
    .D(_01062_),
    .Q(\count_cycle[38] ));
 sky130_fd_sc_hd__dfxtp_1 _17894_ (.CLK(clknet_leaf_93_clk),
    .D(_01063_),
    .Q(\count_cycle[39] ));
 sky130_fd_sc_hd__dfxtp_1 _17895_ (.CLK(clknet_leaf_96_clk),
    .D(_01064_),
    .Q(\count_cycle[40] ));
 sky130_fd_sc_hd__dfxtp_1 _17896_ (.CLK(clknet_leaf_95_clk),
    .D(_01065_),
    .Q(\count_cycle[41] ));
 sky130_fd_sc_hd__dfxtp_1 _17897_ (.CLK(clknet_leaf_95_clk),
    .D(_01066_),
    .Q(\count_cycle[42] ));
 sky130_fd_sc_hd__dfxtp_1 _17898_ (.CLK(clknet_leaf_94_clk),
    .D(_01067_),
    .Q(\count_cycle[43] ));
 sky130_fd_sc_hd__dfxtp_1 _17899_ (.CLK(clknet_leaf_95_clk),
    .D(_01068_),
    .Q(\count_cycle[44] ));
 sky130_fd_sc_hd__dfxtp_1 _17900_ (.CLK(clknet_leaf_94_clk),
    .D(_01069_),
    .Q(\count_cycle[45] ));
 sky130_fd_sc_hd__dfxtp_1 _17901_ (.CLK(clknet_leaf_94_clk),
    .D(_01070_),
    .Q(\count_cycle[46] ));
 sky130_fd_sc_hd__dfxtp_1 _17902_ (.CLK(clknet_leaf_87_clk),
    .D(_01071_),
    .Q(\count_cycle[47] ));
 sky130_fd_sc_hd__dfxtp_1 _17903_ (.CLK(clknet_leaf_87_clk),
    .D(_01072_),
    .Q(\count_cycle[48] ));
 sky130_fd_sc_hd__dfxtp_1 _17904_ (.CLK(clknet_leaf_87_clk),
    .D(_01073_),
    .Q(\count_cycle[49] ));
 sky130_fd_sc_hd__dfxtp_1 _17905_ (.CLK(clknet_leaf_88_clk),
    .D(_01074_),
    .Q(\count_cycle[50] ));
 sky130_fd_sc_hd__dfxtp_1 _17906_ (.CLK(clknet_leaf_87_clk),
    .D(_01075_),
    .Q(\count_cycle[51] ));
 sky130_fd_sc_hd__dfxtp_1 _17907_ (.CLK(clknet_leaf_85_clk),
    .D(_01076_),
    .Q(\count_cycle[52] ));
 sky130_fd_sc_hd__dfxtp_1 _17908_ (.CLK(clknet_leaf_85_clk),
    .D(_01077_),
    .Q(\count_cycle[53] ));
 sky130_fd_sc_hd__dfxtp_1 _17909_ (.CLK(clknet_leaf_85_clk),
    .D(_01078_),
    .Q(\count_cycle[54] ));
 sky130_fd_sc_hd__dfxtp_1 _17910_ (.CLK(clknet_leaf_85_clk),
    .D(_01079_),
    .Q(\count_cycle[55] ));
 sky130_fd_sc_hd__dfxtp_1 _17911_ (.CLK(clknet_leaf_85_clk),
    .D(_01080_),
    .Q(\count_cycle[56] ));
 sky130_fd_sc_hd__dfxtp_1 _17912_ (.CLK(clknet_leaf_84_clk),
    .D(_01081_),
    .Q(\count_cycle[57] ));
 sky130_fd_sc_hd__dfxtp_1 _17913_ (.CLK(clknet_leaf_84_clk),
    .D(_01082_),
    .Q(\count_cycle[58] ));
 sky130_fd_sc_hd__dfxtp_1 _17914_ (.CLK(clknet_leaf_84_clk),
    .D(_01083_),
    .Q(\count_cycle[59] ));
 sky130_fd_sc_hd__dfxtp_1 _17915_ (.CLK(clknet_leaf_82_clk),
    .D(_01084_),
    .Q(\count_cycle[60] ));
 sky130_fd_sc_hd__dfxtp_1 _17916_ (.CLK(clknet_leaf_82_clk),
    .D(_01085_),
    .Q(\count_cycle[61] ));
 sky130_fd_sc_hd__dfxtp_1 _17917_ (.CLK(clknet_leaf_82_clk),
    .D(_01086_),
    .Q(\count_cycle[62] ));
 sky130_fd_sc_hd__dfxtp_1 _17918_ (.CLK(clknet_leaf_81_clk),
    .D(_01087_),
    .Q(\count_cycle[63] ));
 sky130_fd_sc_hd__dfxtp_2 _17919_ (.CLK(clknet_leaf_69_clk),
    .D(_01088_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_1 _17920_ (.CLK(clknet_leaf_64_clk),
    .D(_08369_),
    .Q(\reg_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _17921_ (.CLK(clknet_leaf_54_clk),
    .D(_08380_),
    .Q(\reg_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _17922_ (.CLK(clknet_leaf_26_clk),
    .D(_08391_),
    .Q(\reg_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _17923_ (.CLK(clknet_leaf_54_clk),
    .D(_08394_),
    .Q(\reg_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _17924_ (.CLK(clknet_leaf_56_clk),
    .D(_08395_),
    .Q(\reg_out[4] ));
 sky130_fd_sc_hd__dfxtp_1 _17925_ (.CLK(clknet_leaf_61_clk),
    .D(_08396_),
    .Q(\reg_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _17926_ (.CLK(clknet_leaf_54_clk),
    .D(_08397_),
    .Q(\reg_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _17927_ (.CLK(clknet_leaf_55_clk),
    .D(_08398_),
    .Q(\reg_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _17928_ (.CLK(clknet_leaf_55_clk),
    .D(_08399_),
    .Q(\reg_out[8] ));
 sky130_fd_sc_hd__dfxtp_1 _17929_ (.CLK(clknet_leaf_65_clk),
    .D(_08400_),
    .Q(\reg_out[9] ));
 sky130_fd_sc_hd__dfxtp_1 _17930_ (.CLK(clknet_leaf_62_clk),
    .D(_08370_),
    .Q(\reg_out[10] ));
 sky130_fd_sc_hd__dfxtp_1 _17931_ (.CLK(clknet_leaf_55_clk),
    .D(_08371_),
    .Q(\reg_out[11] ));
 sky130_fd_sc_hd__dfxtp_1 _17932_ (.CLK(clknet_leaf_50_clk),
    .D(_08372_),
    .Q(\reg_out[12] ));
 sky130_fd_sc_hd__dfxtp_1 _17933_ (.CLK(clknet_leaf_66_clk),
    .D(_08373_),
    .Q(\reg_out[13] ));
 sky130_fd_sc_hd__dfxtp_1 _17934_ (.CLK(clknet_leaf_69_clk),
    .D(_08374_),
    .Q(\reg_out[14] ));
 sky130_fd_sc_hd__dfxtp_1 _17935_ (.CLK(clknet_leaf_68_clk),
    .D(_08375_),
    .Q(\reg_out[15] ));
 sky130_fd_sc_hd__dfxtp_1 _17936_ (.CLK(clknet_leaf_50_clk),
    .D(_08376_),
    .Q(\reg_out[16] ));
 sky130_fd_sc_hd__dfxtp_1 _17937_ (.CLK(clknet_leaf_66_clk),
    .D(_08377_),
    .Q(\reg_out[17] ));
 sky130_fd_sc_hd__dfxtp_1 _17938_ (.CLK(clknet_leaf_69_clk),
    .D(_08378_),
    .Q(\reg_out[18] ));
 sky130_fd_sc_hd__dfxtp_1 _17939_ (.CLK(clknet_leaf_68_clk),
    .D(_08379_),
    .Q(\reg_out[19] ));
 sky130_fd_sc_hd__dfxtp_1 _17940_ (.CLK(clknet_leaf_67_clk),
    .D(_08381_),
    .Q(\reg_out[20] ));
 sky130_fd_sc_hd__dfxtp_1 _17941_ (.CLK(clknet_leaf_67_clk),
    .D(_08382_),
    .Q(\reg_out[21] ));
 sky130_fd_sc_hd__dfxtp_1 _17942_ (.CLK(clknet_leaf_67_clk),
    .D(_08383_),
    .Q(\reg_out[22] ));
 sky130_fd_sc_hd__dfxtp_1 _17943_ (.CLK(clknet_leaf_67_clk),
    .D(_08384_),
    .Q(\reg_out[23] ));
 sky130_fd_sc_hd__dfxtp_1 _17944_ (.CLK(clknet_leaf_70_clk),
    .D(_08385_),
    .Q(\reg_out[24] ));
 sky130_fd_sc_hd__dfxtp_1 _17945_ (.CLK(clknet_leaf_78_clk),
    .D(_08386_),
    .Q(\reg_out[25] ));
 sky130_fd_sc_hd__dfxtp_1 _17946_ (.CLK(clknet_leaf_78_clk),
    .D(_08387_),
    .Q(\reg_out[26] ));
 sky130_fd_sc_hd__dfxtp_1 _17947_ (.CLK(clknet_leaf_74_clk),
    .D(_08388_),
    .Q(\reg_out[27] ));
 sky130_fd_sc_hd__dfxtp_1 _17948_ (.CLK(clknet_leaf_70_clk),
    .D(_08389_),
    .Q(\reg_out[28] ));
 sky130_fd_sc_hd__dfxtp_1 _17949_ (.CLK(clknet_leaf_77_clk),
    .D(_08390_),
    .Q(\reg_out[29] ));
 sky130_fd_sc_hd__dfxtp_1 _17950_ (.CLK(clknet_leaf_70_clk),
    .D(_08392_),
    .Q(\reg_out[30] ));
 sky130_fd_sc_hd__dfxtp_1 _17951_ (.CLK(clknet_leaf_70_clk),
    .D(_08393_),
    .Q(\reg_out[31] ));
 sky130_fd_sc_hd__dfxtp_1 _17952_ (.CLK(clknet_leaf_191_clk),
    .D(_01089_),
    .Q(net183));
 sky130_fd_sc_hd__dfxtp_1 _17953_ (.CLK(clknet_leaf_191_clk),
    .D(_01090_),
    .Q(net186));
 sky130_fd_sc_hd__dfxtp_1 _17954_ (.CLK(clknet_leaf_191_clk),
    .D(_01091_),
    .Q(net187));
 sky130_fd_sc_hd__dfxtp_1 _17955_ (.CLK(clknet_leaf_191_clk),
    .D(_01092_),
    .Q(net188));
 sky130_fd_sc_hd__dfxtp_1 _17956_ (.CLK(clknet_leaf_191_clk),
    .D(_01093_),
    .Q(net189));
 sky130_fd_sc_hd__dfxtp_1 _17957_ (.CLK(clknet_leaf_191_clk),
    .D(_01094_),
    .Q(net190));
 sky130_fd_sc_hd__dfxtp_1 _17958_ (.CLK(clknet_leaf_191_clk),
    .D(_01095_),
    .Q(net191));
 sky130_fd_sc_hd__dfxtp_1 _17959_ (.CLK(clknet_leaf_191_clk),
    .D(_01096_),
    .Q(net192));
 sky130_fd_sc_hd__dfxtp_1 _17960_ (.CLK(clknet_leaf_191_clk),
    .D(_01097_),
    .Q(net163));
 sky130_fd_sc_hd__dfxtp_1 _17961_ (.CLK(clknet_leaf_191_clk),
    .D(_01098_),
    .Q(net164));
 sky130_fd_sc_hd__dfxtp_1 _17962_ (.CLK(clknet_leaf_191_clk),
    .D(_01099_),
    .Q(net165));
 sky130_fd_sc_hd__dfxtp_1 _17963_ (.CLK(clknet_leaf_191_clk),
    .D(_01100_),
    .Q(net166));
 sky130_fd_sc_hd__dfxtp_1 _17964_ (.CLK(clknet_leaf_191_clk),
    .D(_01101_),
    .Q(net167));
 sky130_fd_sc_hd__dfxtp_1 _17965_ (.CLK(clknet_leaf_0_clk),
    .D(_01102_),
    .Q(net168));
 sky130_fd_sc_hd__dfxtp_1 _17966_ (.CLK(clknet_leaf_0_clk),
    .D(_01103_),
    .Q(net169));
 sky130_fd_sc_hd__dfxtp_1 _17967_ (.CLK(clknet_leaf_0_clk),
    .D(_01104_),
    .Q(net170));
 sky130_fd_sc_hd__dfxtp_1 _17968_ (.CLK(clknet_leaf_4_clk),
    .D(_01105_),
    .Q(net171));
 sky130_fd_sc_hd__dfxtp_1 _17969_ (.CLK(clknet_leaf_4_clk),
    .D(_01106_),
    .Q(net172));
 sky130_fd_sc_hd__dfxtp_1 _17970_ (.CLK(clknet_leaf_4_clk),
    .D(_01107_),
    .Q(net173));
 sky130_fd_sc_hd__dfxtp_1 _17971_ (.CLK(clknet_leaf_4_clk),
    .D(_01108_),
    .Q(net174));
 sky130_fd_sc_hd__dfxtp_2 _17972_ (.CLK(clknet_leaf_44_clk),
    .D(_01109_),
    .Q(net175));
 sky130_fd_sc_hd__dfxtp_2 _17973_ (.CLK(clknet_leaf_44_clk),
    .D(_01110_),
    .Q(net176));
 sky130_fd_sc_hd__dfxtp_2 _17974_ (.CLK(clknet_leaf_43_clk),
    .D(_01111_),
    .Q(net177));
 sky130_fd_sc_hd__dfxtp_2 _17975_ (.CLK(clknet_leaf_44_clk),
    .D(_01112_),
    .Q(net178));
 sky130_fd_sc_hd__dfxtp_2 _17976_ (.CLK(clknet_leaf_44_clk),
    .D(_01113_),
    .Q(net179));
 sky130_fd_sc_hd__dfxtp_2 _17977_ (.CLK(clknet_leaf_44_clk),
    .D(_01114_),
    .Q(net180));
 sky130_fd_sc_hd__dfxtp_2 _17978_ (.CLK(clknet_leaf_44_clk),
    .D(_01115_),
    .Q(net181));
 sky130_fd_sc_hd__dfxtp_2 _17979_ (.CLK(clknet_leaf_43_clk),
    .D(_01116_),
    .Q(net182));
 sky130_fd_sc_hd__dfxtp_2 _17980_ (.CLK(clknet_leaf_44_clk),
    .D(_01117_),
    .Q(net184));
 sky130_fd_sc_hd__dfxtp_2 _17981_ (.CLK(clknet_leaf_43_clk),
    .D(_01118_),
    .Q(net185));
 sky130_fd_sc_hd__dfxtp_1 _17982_ (.CLK(clknet_leaf_63_clk),
    .D(_01119_),
    .Q(irq_delay));
 sky130_fd_sc_hd__dfxtp_4 _17983_ (.CLK(clknet_leaf_63_clk),
    .D(_01120_),
    .Q(irq_active));
 sky130_fd_sc_hd__dfxtp_1 _17984_ (.CLK(clknet_leaf_103_clk),
    .D(_01121_),
    .Q(\irq_mask[0] ));
 sky130_fd_sc_hd__dfxtp_2 _17985_ (.CLK(clknet_leaf_103_clk),
    .D(_01122_),
    .Q(\irq_mask[1] ));
 sky130_fd_sc_hd__dfxtp_4 _17986_ (.CLK(clknet_leaf_103_clk),
    .D(_01123_),
    .Q(\irq_mask[2] ));
 sky130_fd_sc_hd__dfxtp_1 _17987_ (.CLK(clknet_leaf_105_clk),
    .D(_01124_),
    .Q(\irq_mask[3] ));
 sky130_fd_sc_hd__dfxtp_1 _17988_ (.CLK(clknet_leaf_105_clk),
    .D(_01125_),
    .Q(\irq_mask[4] ));
 sky130_fd_sc_hd__dfxtp_1 _17989_ (.CLK(clknet_leaf_105_clk),
    .D(_01126_),
    .Q(\irq_mask[5] ));
 sky130_fd_sc_hd__dfxtp_1 _17990_ (.CLK(clknet_leaf_105_clk),
    .D(_01127_),
    .Q(\irq_mask[6] ));
 sky130_fd_sc_hd__dfxtp_1 _17991_ (.CLK(clknet_leaf_104_clk),
    .D(_01128_),
    .Q(\irq_mask[7] ));
 sky130_fd_sc_hd__dfxtp_1 _17992_ (.CLK(clknet_leaf_104_clk),
    .D(_01129_),
    .Q(\irq_mask[8] ));
 sky130_fd_sc_hd__dfxtp_1 _17993_ (.CLK(clknet_leaf_103_clk),
    .D(_01130_),
    .Q(\irq_mask[9] ));
 sky130_fd_sc_hd__dfxtp_1 _17994_ (.CLK(clknet_leaf_103_clk),
    .D(_01131_),
    .Q(\irq_mask[10] ));
 sky130_fd_sc_hd__dfxtp_1 _17995_ (.CLK(clknet_leaf_65_clk),
    .D(_01132_),
    .Q(\irq_mask[11] ));
 sky130_fd_sc_hd__dfxtp_1 _17996_ (.CLK(clknet_leaf_65_clk),
    .D(_01133_),
    .Q(\irq_mask[12] ));
 sky130_fd_sc_hd__dfxtp_1 _17997_ (.CLK(clknet_leaf_103_clk),
    .D(_01134_),
    .Q(\irq_mask[13] ));
 sky130_fd_sc_hd__dfxtp_1 _17998_ (.CLK(clknet_leaf_103_clk),
    .D(_01135_),
    .Q(\irq_mask[14] ));
 sky130_fd_sc_hd__dfxtp_1 _17999_ (.CLK(clknet_leaf_80_clk),
    .D(_01136_),
    .Q(\irq_mask[15] ));
 sky130_fd_sc_hd__dfxtp_1 _18000_ (.CLK(clknet_leaf_79_clk),
    .D(_01137_),
    .Q(\irq_mask[16] ));
 sky130_fd_sc_hd__dfxtp_1 _18001_ (.CLK(clknet_leaf_66_clk),
    .D(_01138_),
    .Q(\irq_mask[17] ));
 sky130_fd_sc_hd__dfxtp_1 _18002_ (.CLK(clknet_leaf_66_clk),
    .D(_01139_),
    .Q(\irq_mask[18] ));
 sky130_fd_sc_hd__dfxtp_1 _18003_ (.CLK(clknet_leaf_66_clk),
    .D(_01140_),
    .Q(\irq_mask[19] ));
 sky130_fd_sc_hd__dfxtp_1 _18004_ (.CLK(clknet_leaf_66_clk),
    .D(_01141_),
    .Q(\irq_mask[20] ));
 sky130_fd_sc_hd__dfxtp_1 _18005_ (.CLK(clknet_leaf_79_clk),
    .D(_01142_),
    .Q(\irq_mask[21] ));
 sky130_fd_sc_hd__dfxtp_1 _18006_ (.CLK(clknet_leaf_80_clk),
    .D(_01143_),
    .Q(\irq_mask[22] ));
 sky130_fd_sc_hd__dfxtp_1 _18007_ (.CLK(clknet_leaf_78_clk),
    .D(_01144_),
    .Q(\irq_mask[23] ));
 sky130_fd_sc_hd__dfxtp_1 _18008_ (.CLK(clknet_leaf_78_clk),
    .D(_01145_),
    .Q(\irq_mask[24] ));
 sky130_fd_sc_hd__dfxtp_1 _18009_ (.CLK(clknet_leaf_78_clk),
    .D(_01146_),
    .Q(\irq_mask[25] ));
 sky130_fd_sc_hd__dfxtp_1 _18010_ (.CLK(clknet_leaf_78_clk),
    .D(_01147_),
    .Q(\irq_mask[26] ));
 sky130_fd_sc_hd__dfxtp_1 _18011_ (.CLK(clknet_leaf_79_clk),
    .D(_01148_),
    .Q(\irq_mask[27] ));
 sky130_fd_sc_hd__dfxtp_1 _18012_ (.CLK(clknet_leaf_76_clk),
    .D(_01149_),
    .Q(\irq_mask[28] ));
 sky130_fd_sc_hd__dfxtp_1 _18013_ (.CLK(clknet_leaf_76_clk),
    .D(_01150_),
    .Q(\irq_mask[29] ));
 sky130_fd_sc_hd__dfxtp_1 _18014_ (.CLK(clknet_leaf_77_clk),
    .D(_01151_),
    .Q(\irq_mask[30] ));
 sky130_fd_sc_hd__dfxtp_1 _18015_ (.CLK(clknet_leaf_76_clk),
    .D(_01152_),
    .Q(\irq_mask[31] ));
 sky130_fd_sc_hd__dfxtp_1 _18016_ (.CLK(clknet_leaf_104_clk),
    .D(_00001_),
    .Q(\irq_pending[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18017_ (.CLK(clknet_leaf_64_clk),
    .D(_00012_),
    .Q(\irq_pending[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18018_ (.CLK(clknet_leaf_64_clk),
    .D(_00023_),
    .Q(\irq_pending[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18019_ (.CLK(clknet_leaf_104_clk),
    .D(_00026_),
    .Q(\irq_pending[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18020_ (.CLK(clknet_leaf_105_clk),
    .D(_00027_),
    .Q(\irq_pending[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18021_ (.CLK(clknet_leaf_104_clk),
    .D(_00028_),
    .Q(\irq_pending[5] ));
 sky130_fd_sc_hd__dfxtp_2 _18022_ (.CLK(clknet_leaf_105_clk),
    .D(_00029_),
    .Q(\irq_pending[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18023_ (.CLK(clknet_leaf_104_clk),
    .D(_00030_),
    .Q(\irq_pending[7] ));
 sky130_fd_sc_hd__dfxtp_1 _18024_ (.CLK(clknet_leaf_104_clk),
    .D(_00031_),
    .Q(\irq_pending[8] ));
 sky130_fd_sc_hd__dfxtp_1 _18025_ (.CLK(clknet_leaf_64_clk),
    .D(_00032_),
    .Q(\irq_pending[9] ));
 sky130_fd_sc_hd__dfxtp_1 _18026_ (.CLK(clknet_leaf_65_clk),
    .D(_00002_),
    .Q(\irq_pending[10] ));
 sky130_fd_sc_hd__dfxtp_1 _18027_ (.CLK(clknet_leaf_65_clk),
    .D(_00003_),
    .Q(\irq_pending[11] ));
 sky130_fd_sc_hd__dfxtp_1 _18028_ (.CLK(clknet_leaf_65_clk),
    .D(_00004_),
    .Q(\irq_pending[12] ));
 sky130_fd_sc_hd__dfxtp_1 _18029_ (.CLK(clknet_leaf_65_clk),
    .D(_00005_),
    .Q(\irq_pending[13] ));
 sky130_fd_sc_hd__dfxtp_1 _18030_ (.CLK(clknet_leaf_66_clk),
    .D(_00006_),
    .Q(\irq_pending[14] ));
 sky130_fd_sc_hd__dfxtp_1 _18031_ (.CLK(clknet_leaf_66_clk),
    .D(_00007_),
    .Q(\irq_pending[15] ));
 sky130_fd_sc_hd__dfxtp_1 _18032_ (.CLK(clknet_leaf_80_clk),
    .D(_00008_),
    .Q(\irq_pending[16] ));
 sky130_fd_sc_hd__dfxtp_1 _18033_ (.CLK(clknet_leaf_66_clk),
    .D(_00009_),
    .Q(\irq_pending[17] ));
 sky130_fd_sc_hd__dfxtp_1 _18034_ (.CLK(clknet_leaf_66_clk),
    .D(_00010_),
    .Q(\irq_pending[18] ));
 sky130_fd_sc_hd__dfxtp_1 _18035_ (.CLK(clknet_leaf_66_clk),
    .D(_00011_),
    .Q(\irq_pending[19] ));
 sky130_fd_sc_hd__dfxtp_1 _18036_ (.CLK(clknet_leaf_79_clk),
    .D(_00013_),
    .Q(\irq_pending[20] ));
 sky130_fd_sc_hd__dfxtp_1 _18037_ (.CLK(clknet_leaf_79_clk),
    .D(_00014_),
    .Q(\irq_pending[21] ));
 sky130_fd_sc_hd__dfxtp_1 _18038_ (.CLK(clknet_leaf_80_clk),
    .D(_00015_),
    .Q(\irq_pending[22] ));
 sky130_fd_sc_hd__dfxtp_1 _18039_ (.CLK(clknet_leaf_67_clk),
    .D(_00016_),
    .Q(\irq_pending[23] ));
 sky130_fd_sc_hd__dfxtp_1 _18040_ (.CLK(clknet_leaf_78_clk),
    .D(_00017_),
    .Q(\irq_pending[24] ));
 sky130_fd_sc_hd__dfxtp_1 _18041_ (.CLK(clknet_leaf_78_clk),
    .D(_00018_),
    .Q(\irq_pending[25] ));
 sky130_fd_sc_hd__dfxtp_1 _18042_ (.CLK(clknet_leaf_78_clk),
    .D(_00019_),
    .Q(\irq_pending[26] ));
 sky130_fd_sc_hd__dfxtp_1 _18043_ (.CLK(clknet_leaf_82_clk),
    .D(_00020_),
    .Q(\irq_pending[27] ));
 sky130_fd_sc_hd__dfxtp_1 _18044_ (.CLK(clknet_leaf_76_clk),
    .D(_00021_),
    .Q(\irq_pending[28] ));
 sky130_fd_sc_hd__dfxtp_1 _18045_ (.CLK(clknet_leaf_82_clk),
    .D(_00022_),
    .Q(\irq_pending[29] ));
 sky130_fd_sc_hd__dfxtp_1 _18046_ (.CLK(clknet_leaf_77_clk),
    .D(_00024_),
    .Q(\irq_pending[30] ));
 sky130_fd_sc_hd__dfxtp_1 _18047_ (.CLK(clknet_leaf_77_clk),
    .D(_00025_),
    .Q(\irq_pending[31] ));
 sky130_fd_sc_hd__dfxtp_4 _18048_ (.CLK(clknet_leaf_51_clk),
    .D(_01153_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_4 _18049_ (.CLK(clknet_leaf_45_clk),
    .D(_01154_),
    .Q(net110));
 sky130_fd_sc_hd__dfxtp_4 _18050_ (.CLK(clknet_leaf_45_clk),
    .D(_01155_),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_2 _18051_ (.CLK(clknet_leaf_45_clk),
    .D(_01156_),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_4 _18052_ (.CLK(clknet_leaf_52_clk),
    .D(_01157_),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_4 _18053_ (.CLK(clknet_leaf_20_clk),
    .D(_01158_),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_4 _18054_ (.CLK(clknet_leaf_20_clk),
    .D(_01159_),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_4 _18055_ (.CLK(clknet_leaf_59_clk),
    .D(_01160_),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_4 _18056_ (.CLK(clknet_leaf_47_clk),
    .D(_01161_),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_4 _18057_ (.CLK(clknet_leaf_71_clk),
    .D(_01162_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_4 _18058_ (.CLK(clknet_leaf_73_clk),
    .D(_01163_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_4 _18059_ (.CLK(clknet_leaf_73_clk),
    .D(_01164_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_4 _18060_ (.CLK(clknet_leaf_73_clk),
    .D(_01165_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_4 _18061_ (.CLK(clknet_leaf_73_clk),
    .D(_01166_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_4 _18062_ (.CLK(clknet_leaf_73_clk),
    .D(_01167_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_4 _18063_ (.CLK(clknet_leaf_73_clk),
    .D(_01168_),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_4 _18064_ (.CLK(clknet_leaf_73_clk),
    .D(_01169_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_4 _18065_ (.CLK(clknet_leaf_72_clk),
    .D(_01170_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_2 _18066_ (.CLK(clknet_leaf_72_clk),
    .D(_01171_),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_4 _18067_ (.CLK(clknet_leaf_72_clk),
    .D(_01172_),
    .Q(net109));
 sky130_fd_sc_hd__dfxtp_4 _18068_ (.CLK(clknet_leaf_73_clk),
    .D(_01173_),
    .Q(net111));
 sky130_fd_sc_hd__dfxtp_4 _18069_ (.CLK(clknet_leaf_73_clk),
    .D(_01174_),
    .Q(net112));
 sky130_fd_sc_hd__dfxtp_4 _18070_ (.CLK(clknet_leaf_73_clk),
    .D(_01175_),
    .Q(net113));
 sky130_fd_sc_hd__dfxtp_4 _18071_ (.CLK(clknet_leaf_72_clk),
    .D(_01176_),
    .Q(net114));
 sky130_fd_sc_hd__dfxtp_2 _18072_ (.CLK(clknet_leaf_73_clk),
    .D(_01177_),
    .Q(net115));
 sky130_fd_sc_hd__dfxtp_4 _18073_ (.CLK(clknet_leaf_74_clk),
    .D(_01178_),
    .Q(net116));
 sky130_fd_sc_hd__dfxtp_2 _18074_ (.CLK(clknet_leaf_48_clk),
    .D(_01179_),
    .Q(net117));
 sky130_fd_sc_hd__dfxtp_4 _18075_ (.CLK(clknet_leaf_75_clk),
    .D(_01180_),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_4 _18076_ (.CLK(clknet_leaf_75_clk),
    .D(_01181_),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_4 _18077_ (.CLK(clknet_leaf_73_clk),
    .D(_01182_),
    .Q(net120));
 sky130_fd_sc_hd__dfxtp_4 _18078_ (.CLK(clknet_leaf_73_clk),
    .D(_01183_),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_2 _18079_ (.CLK(clknet_leaf_47_clk),
    .D(_01184_),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_2 _18080_ (.CLK(clknet_leaf_26_clk),
    .D(_01185_),
    .Q(mem_do_prefetch));
 sky130_fd_sc_hd__dfxtp_1 _18081_ (.CLK(clknet_leaf_40_clk),
    .D(_01186_),
    .Q(mem_do_rinst));
 sky130_fd_sc_hd__dfxtp_1 _18082_ (.CLK(clknet_leaf_39_clk),
    .D(_01187_),
    .Q(mem_do_rdata));
 sky130_fd_sc_hd__dfxtp_2 _18083_ (.CLK(clknet_leaf_27_clk),
    .D(_01188_),
    .Q(mem_do_wdata));
 sky130_fd_sc_hd__dfxtp_4 _18084_ (.CLK(clknet_leaf_27_clk),
    .D(_00000_),
    .Q(decoder_trigger));
 sky130_fd_sc_hd__dfxtp_1 _18085_ (.CLK(clknet_leaf_102_clk),
    .D(_01189_),
    .Q(\timer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18086_ (.CLK(clknet_leaf_102_clk),
    .D(_01190_),
    .Q(\timer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18087_ (.CLK(clknet_leaf_102_clk),
    .D(_01191_),
    .Q(\timer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18088_ (.CLK(clknet_leaf_102_clk),
    .D(_01192_),
    .Q(\timer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18089_ (.CLK(clknet_leaf_101_clk),
    .D(_01193_),
    .Q(\timer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18090_ (.CLK(clknet_leaf_100_clk),
    .D(_01194_),
    .Q(\timer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18091_ (.CLK(clknet_leaf_102_clk),
    .D(_01195_),
    .Q(\timer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18092_ (.CLK(clknet_leaf_100_clk),
    .D(_01196_),
    .Q(\timer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _18093_ (.CLK(clknet_leaf_102_clk),
    .D(_01197_),
    .Q(\timer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _18094_ (.CLK(clknet_leaf_103_clk),
    .D(_01198_),
    .Q(\timer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _18095_ (.CLK(clknet_leaf_91_clk),
    .D(_01199_),
    .Q(\timer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _18096_ (.CLK(clknet_leaf_92_clk),
    .D(_01200_),
    .Q(\timer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _18097_ (.CLK(clknet_leaf_92_clk),
    .D(_01201_),
    .Q(\timer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _18098_ (.CLK(clknet_leaf_92_clk),
    .D(_01202_),
    .Q(\timer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _18099_ (.CLK(clknet_leaf_91_clk),
    .D(_01203_),
    .Q(\timer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _18100_ (.CLK(clknet_leaf_90_clk),
    .D(_01204_),
    .Q(\timer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _18101_ (.CLK(clknet_leaf_90_clk),
    .D(_01205_),
    .Q(\timer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _18102_ (.CLK(clknet_leaf_91_clk),
    .D(_01206_),
    .Q(\timer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _18103_ (.CLK(clknet_leaf_80_clk),
    .D(_01207_),
    .Q(\timer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _18104_ (.CLK(clknet_leaf_90_clk),
    .D(_01208_),
    .Q(\timer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _18105_ (.CLK(clknet_leaf_90_clk),
    .D(_01209_),
    .Q(\timer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _18106_ (.CLK(clknet_leaf_90_clk),
    .D(_01210_),
    .Q(\timer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _18107_ (.CLK(clknet_leaf_89_clk),
    .D(_01211_),
    .Q(\timer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _18108_ (.CLK(clknet_leaf_81_clk),
    .D(_01212_),
    .Q(\timer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _18109_ (.CLK(clknet_leaf_81_clk),
    .D(_01213_),
    .Q(\timer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _18110_ (.CLK(clknet_leaf_81_clk),
    .D(_01214_),
    .Q(\timer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _18111_ (.CLK(clknet_leaf_81_clk),
    .D(_01215_),
    .Q(\timer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _18112_ (.CLK(clknet_leaf_81_clk),
    .D(_01216_),
    .Q(\timer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _18113_ (.CLK(clknet_leaf_81_clk),
    .D(_01217_),
    .Q(\timer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _18114_ (.CLK(clknet_leaf_82_clk),
    .D(_01218_),
    .Q(\timer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _18115_ (.CLK(clknet_leaf_82_clk),
    .D(_01219_),
    .Q(\timer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _18116_ (.CLK(clknet_leaf_82_clk),
    .D(_01220_),
    .Q(\timer[31] ));
 sky130_fd_sc_hd__dfxtp_2 _18117_ (.CLK(clknet_leaf_63_clk),
    .D(_01221_),
    .Q(\irq_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _18118_ (.CLK(clknet_leaf_63_clk),
    .D(_01222_),
    .Q(\irq_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _18119_ (.CLK(clknet_leaf_53_clk),
    .D(_01223_),
    .Q(latched_store));
 sky130_fd_sc_hd__dfxtp_2 _18120_ (.CLK(clknet_leaf_54_clk),
    .D(_01224_),
    .Q(latched_stalu));
 sky130_fd_sc_hd__dfxtp_4 _18121_ (.CLK(clknet_leaf_55_clk),
    .D(_01225_),
    .Q(latched_branch));
 sky130_fd_sc_hd__dfxtp_1 _18122_ (.CLK(clknet_leaf_27_clk),
    .D(_01226_),
    .Q(decoder_pseudo_trigger));
 sky130_fd_sc_hd__dfxtp_1 _18123_ (.CLK(clknet_leaf_41_clk),
    .D(_01227_),
    .Q(latched_is_lh));
 sky130_fd_sc_hd__dfxtp_1 _18124_ (.CLK(clknet_leaf_40_clk),
    .D(_01228_),
    .Q(latched_is_lb));
 sky130_fd_sc_hd__dfxtp_2 _18125_ (.CLK(clknet_leaf_21_clk),
    .D(_01229_),
    .Q(latched_compr));
 sky130_fd_sc_hd__dfxtp_1 _18126_ (.CLK(clknet_leaf_42_clk),
    .D(\alu_out[0] ),
    .Q(\alu_out_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18127_ (.CLK(clknet_leaf_29_clk),
    .D(\alu_out[1] ),
    .Q(\alu_out_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18128_ (.CLK(clknet_leaf_26_clk),
    .D(\alu_out[2] ),
    .Q(\alu_out_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18129_ (.CLK(clknet_leaf_26_clk),
    .D(\alu_out[3] ),
    .Q(\alu_out_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18130_ (.CLK(clknet_leaf_27_clk),
    .D(\alu_out[4] ),
    .Q(\alu_out_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18131_ (.CLK(clknet_leaf_40_clk),
    .D(\alu_out[5] ),
    .Q(\alu_out_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18132_ (.CLK(clknet_leaf_28_clk),
    .D(\alu_out[6] ),
    .Q(\alu_out_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18133_ (.CLK(clknet_leaf_40_clk),
    .D(\alu_out[7] ),
    .Q(\alu_out_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _18134_ (.CLK(clknet_leaf_42_clk),
    .D(\alu_out[8] ),
    .Q(\alu_out_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _18135_ (.CLK(clknet_leaf_50_clk),
    .D(\alu_out[9] ),
    .Q(\alu_out_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _18136_ (.CLK(clknet_leaf_48_clk),
    .D(\alu_out[10] ),
    .Q(\alu_out_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _18137_ (.CLK(clknet_leaf_47_clk),
    .D(\alu_out[11] ),
    .Q(\alu_out_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _18138_ (.CLK(clknet_leaf_41_clk),
    .D(\alu_out[12] ),
    .Q(\alu_out_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _18139_ (.CLK(clknet_leaf_71_clk),
    .D(\alu_out[13] ),
    .Q(\alu_out_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _18140_ (.CLK(clknet_leaf_46_clk),
    .D(\alu_out[14] ),
    .Q(\alu_out_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _18141_ (.CLK(clknet_leaf_47_clk),
    .D(\alu_out[15] ),
    .Q(\alu_out_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _18142_ (.CLK(clknet_leaf_45_clk),
    .D(\alu_out[16] ),
    .Q(\alu_out_q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _18143_ (.CLK(clknet_leaf_46_clk),
    .D(\alu_out[17] ),
    .Q(\alu_out_q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _18144_ (.CLK(clknet_leaf_47_clk),
    .D(\alu_out[18] ),
    .Q(\alu_out_q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _18145_ (.CLK(clknet_leaf_49_clk),
    .D(\alu_out[19] ),
    .Q(\alu_out_q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _18146_ (.CLK(clknet_leaf_70_clk),
    .D(\alu_out[20] ),
    .Q(\alu_out_q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _18147_ (.CLK(clknet_leaf_46_clk),
    .D(\alu_out[21] ),
    .Q(\alu_out_q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _18148_ (.CLK(clknet_leaf_70_clk),
    .D(\alu_out[22] ),
    .Q(\alu_out_q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _18149_ (.CLK(clknet_leaf_70_clk),
    .D(\alu_out[23] ),
    .Q(\alu_out_q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _18150_ (.CLK(clknet_leaf_46_clk),
    .D(\alu_out[24] ),
    .Q(\alu_out_q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _18151_ (.CLK(clknet_leaf_51_clk),
    .D(\alu_out[25] ),
    .Q(\alu_out_q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _18152_ (.CLK(clknet_leaf_45_clk),
    .D(\alu_out[26] ),
    .Q(\alu_out_q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _18153_ (.CLK(clknet_leaf_45_clk),
    .D(\alu_out[27] ),
    .Q(\alu_out_q[27] ));
 sky130_fd_sc_hd__dfxtp_1 _18154_ (.CLK(clknet_leaf_73_clk),
    .D(\alu_out[28] ),
    .Q(\alu_out_q[28] ));
 sky130_fd_sc_hd__dfxtp_1 _18155_ (.CLK(clknet_leaf_46_clk),
    .D(\alu_out[29] ),
    .Q(\alu_out_q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _18156_ (.CLK(clknet_leaf_47_clk),
    .D(\alu_out[30] ),
    .Q(\alu_out_q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _18157_ (.CLK(clknet_leaf_72_clk),
    .D(\alu_out[31] ),
    .Q(\alu_out_q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _18158_ (.CLK(clknet_leaf_40_clk),
    .D(clear_prefetched_high_word),
    .Q(clear_prefetched_high_word_q));
 sky130_fd_sc_hd__dfxtp_1 _18159_ (.CLK(clknet_leaf_21_clk),
    .D(_01230_),
    .Q(do_waitirq));
 sky130_fd_sc_hd__dfxtp_2 _18160_ (.CLK(clknet_leaf_23_clk),
    .D(_01231_),
    .Q(\decoded_imm_j[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18161_ (.CLK(clknet_leaf_23_clk),
    .D(_01232_),
    .Q(\decoded_imm_j[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18162_ (.CLK(clknet_leaf_24_clk),
    .D(_01233_),
    .Q(\decoded_imm_j[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18163_ (.CLK(clknet_leaf_23_clk),
    .D(_01234_),
    .Q(\decoded_imm_j[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18164_ (.CLK(clknet_leaf_24_clk),
    .D(_01235_),
    .Q(\decoded_imm_j[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18165_ (.CLK(clknet_leaf_32_clk),
    .D(_01236_),
    .Q(\decoded_imm_j[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18166_ (.CLK(clknet_leaf_24_clk),
    .D(_01237_),
    .Q(\decoded_imm_j[7] ));
 sky130_fd_sc_hd__dfxtp_1 _18167_ (.CLK(clknet_leaf_32_clk),
    .D(_01238_),
    .Q(\decoded_imm_j[8] ));
 sky130_fd_sc_hd__dfxtp_1 _18168_ (.CLK(clknet_leaf_23_clk),
    .D(_01239_),
    .Q(\decoded_imm_j[9] ));
 sky130_fd_sc_hd__dfxtp_2 _18169_ (.CLK(clknet_leaf_23_clk),
    .D(_01240_),
    .Q(\decoded_imm_j[10] ));
 sky130_fd_sc_hd__dfxtp_1 _18170_ (.CLK(clknet_leaf_24_clk),
    .D(_01241_),
    .Q(\decoded_imm_j[11] ));
 sky130_fd_sc_hd__dfxtp_2 _18171_ (.CLK(clknet_leaf_24_clk),
    .D(_01242_),
    .Q(\decoded_imm_j[12] ));
 sky130_fd_sc_hd__dfxtp_2 _18172_ (.CLK(clknet_leaf_24_clk),
    .D(_01243_),
    .Q(\decoded_imm_j[13] ));
 sky130_fd_sc_hd__dfxtp_2 _18173_ (.CLK(clknet_leaf_24_clk),
    .D(_01244_),
    .Q(\decoded_imm_j[14] ));
 sky130_fd_sc_hd__dfxtp_2 _18174_ (.CLK(clknet_leaf_31_clk),
    .D(_01245_),
    .Q(\decoded_imm_j[15] ));
 sky130_fd_sc_hd__dfxtp_2 _18175_ (.CLK(clknet_leaf_24_clk),
    .D(_01246_),
    .Q(\decoded_imm_j[16] ));
 sky130_fd_sc_hd__dfxtp_2 _18176_ (.CLK(clknet_leaf_31_clk),
    .D(_01247_),
    .Q(\decoded_imm_j[17] ));
 sky130_fd_sc_hd__dfxtp_2 _18177_ (.CLK(clknet_leaf_31_clk),
    .D(_01248_),
    .Q(\decoded_imm_j[18] ));
 sky130_fd_sc_hd__dfxtp_2 _18178_ (.CLK(clknet_leaf_31_clk),
    .D(_01249_),
    .Q(\decoded_imm_j[19] ));
 sky130_fd_sc_hd__dfxtp_1 _18179_ (.CLK(clknet_leaf_22_clk),
    .D(_01250_),
    .Q(\decoded_imm_j[20] ));
 sky130_fd_sc_hd__dfxtp_1 _18180_ (.CLK(clknet_leaf_32_clk),
    .D(_01251_),
    .Q(instr_lui));
 sky130_fd_sc_hd__dfxtp_1 _18181_ (.CLK(clknet_leaf_31_clk),
    .D(_01252_),
    .Q(instr_auipc));
 sky130_fd_sc_hd__dfxtp_4 _18182_ (.CLK(clknet_leaf_32_clk),
    .D(_01253_),
    .Q(instr_jal));
 sky130_fd_sc_hd__dfxtp_1 _18183_ (.CLK(clknet_leaf_41_clk),
    .D(_01254_),
    .Q(instr_beq));
 sky130_fd_sc_hd__dfxtp_1 _18184_ (.CLK(clknet_leaf_43_clk),
    .D(_01255_),
    .Q(instr_bne));
 sky130_fd_sc_hd__dfxtp_1 _18185_ (.CLK(clknet_leaf_43_clk),
    .D(_01256_),
    .Q(instr_blt));
 sky130_fd_sc_hd__dfxtp_1 _18186_ (.CLK(clknet_leaf_43_clk),
    .D(_01257_),
    .Q(instr_bge));
 sky130_fd_sc_hd__dfxtp_1 _18187_ (.CLK(clknet_leaf_43_clk),
    .D(_01258_),
    .Q(instr_bltu));
 sky130_fd_sc_hd__dfxtp_1 _18188_ (.CLK(clknet_leaf_43_clk),
    .D(_01259_),
    .Q(instr_bgeu));
 sky130_fd_sc_hd__dfxtp_2 _18189_ (.CLK(clknet_leaf_31_clk),
    .D(_01260_),
    .Q(instr_jalr));
 sky130_fd_sc_hd__dfxtp_1 _18190_ (.CLK(clknet_leaf_41_clk),
    .D(_01261_),
    .Q(instr_lb));
 sky130_fd_sc_hd__dfxtp_1 _18191_ (.CLK(clknet_leaf_29_clk),
    .D(_01262_),
    .Q(instr_lh));
 sky130_fd_sc_hd__dfxtp_1 _18192_ (.CLK(clknet_leaf_29_clk),
    .D(_01263_),
    .Q(instr_lw));
 sky130_fd_sc_hd__dfxtp_1 _18193_ (.CLK(clknet_leaf_40_clk),
    .D(_01264_),
    .Q(instr_lbu));
 sky130_fd_sc_hd__dfxtp_1 _18194_ (.CLK(clknet_leaf_28_clk),
    .D(_01265_),
    .Q(instr_lhu));
 sky130_fd_sc_hd__dfxtp_1 _18195_ (.CLK(clknet_leaf_41_clk),
    .D(_01266_),
    .Q(instr_sb));
 sky130_fd_sc_hd__dfxtp_1 _18196_ (.CLK(clknet_leaf_29_clk),
    .D(_01267_),
    .Q(instr_sh));
 sky130_fd_sc_hd__dfxtp_1 _18197_ (.CLK(clknet_leaf_41_clk),
    .D(_01268_),
    .Q(instr_addi));
 sky130_fd_sc_hd__dfxtp_1 _18198_ (.CLK(clknet_leaf_43_clk),
    .D(_01269_),
    .Q(instr_slti));
 sky130_fd_sc_hd__dfxtp_1 _18199_ (.CLK(clknet_leaf_43_clk),
    .D(_01270_),
    .Q(instr_sltiu));
 sky130_fd_sc_hd__dfxtp_1 _18200_ (.CLK(clknet_leaf_42_clk),
    .D(_01271_),
    .Q(instr_xori));
 sky130_fd_sc_hd__dfxtp_1 _18201_ (.CLK(clknet_leaf_43_clk),
    .D(_01272_),
    .Q(instr_ori));
 sky130_fd_sc_hd__dfxtp_1 _18202_ (.CLK(clknet_leaf_43_clk),
    .D(_01273_),
    .Q(instr_andi));
 sky130_fd_sc_hd__dfxtp_1 _18203_ (.CLK(clknet_leaf_29_clk),
    .D(_01274_),
    .Q(instr_sw));
 sky130_fd_sc_hd__dfxtp_2 _18204_ (.CLK(clknet_leaf_28_clk),
    .D(_01275_),
    .Q(instr_slli));
 sky130_fd_sc_hd__dfxtp_1 _18205_ (.CLK(clknet_leaf_41_clk),
    .D(_01276_),
    .Q(instr_srli));
 sky130_fd_sc_hd__dfxtp_1 _18206_ (.CLK(clknet_leaf_42_clk),
    .D(_01277_),
    .Q(instr_add));
 sky130_fd_sc_hd__dfxtp_2 _18207_ (.CLK(clknet_leaf_41_clk),
    .D(_01278_),
    .Q(instr_sub));
 sky130_fd_sc_hd__dfxtp_2 _18208_ (.CLK(clknet_leaf_41_clk),
    .D(_01279_),
    .Q(instr_sll));
 sky130_fd_sc_hd__dfxtp_1 _18209_ (.CLK(clknet_leaf_39_clk),
    .D(_01280_),
    .Q(instr_slt));
 sky130_fd_sc_hd__dfxtp_1 _18210_ (.CLK(clknet_leaf_43_clk),
    .D(_01281_),
    .Q(instr_sltu));
 sky130_fd_sc_hd__dfxtp_1 _18211_ (.CLK(clknet_leaf_42_clk),
    .D(_01282_),
    .Q(instr_xor));
 sky130_fd_sc_hd__dfxtp_1 _18212_ (.CLK(clknet_leaf_41_clk),
    .D(_01283_),
    .Q(instr_srl));
 sky130_fd_sc_hd__dfxtp_2 _18213_ (.CLK(clknet_leaf_41_clk),
    .D(_01284_),
    .Q(instr_sra));
 sky130_fd_sc_hd__dfxtp_2 _18214_ (.CLK(clknet_leaf_43_clk),
    .D(_01285_),
    .Q(instr_or));
 sky130_fd_sc_hd__dfxtp_2 _18215_ (.CLK(clknet_leaf_39_clk),
    .D(_01286_),
    .Q(instr_and));
 sky130_fd_sc_hd__dfxtp_2 _18216_ (.CLK(clknet_leaf_28_clk),
    .D(_01287_),
    .Q(instr_srai));
 sky130_fd_sc_hd__dfxtp_1 _18217_ (.CLK(clknet_leaf_102_clk),
    .D(_01288_),
    .Q(instr_rdcycle));
 sky130_fd_sc_hd__dfxtp_4 _18218_ (.CLK(clknet_leaf_92_clk),
    .D(_01289_),
    .Q(instr_rdcycleh));
 sky130_fd_sc_hd__dfxtp_4 _18219_ (.CLK(clknet_leaf_92_clk),
    .D(_01290_),
    .Q(instr_rdinstr));
 sky130_fd_sc_hd__dfxtp_2 _18220_ (.CLK(clknet_leaf_92_clk),
    .D(_01291_),
    .Q(instr_rdinstrh));
 sky130_fd_sc_hd__dfxtp_1 _18221_ (.CLK(clknet_leaf_41_clk),
    .D(_01292_),
    .Q(instr_fence));
 sky130_fd_sc_hd__dfxtp_4 _18222_ (.CLK(clknet_leaf_38_clk),
    .D(_01293_),
    .Q(net262));
 sky130_fd_sc_hd__dfxtp_4 _18223_ (.CLK(clknet_leaf_25_clk),
    .D(_01294_),
    .Q(instr_retirq));
 sky130_fd_sc_hd__dfxtp_2 _18224_ (.CLK(clknet_leaf_65_clk),
    .D(_01295_),
    .Q(instr_maskirq));
 sky130_fd_sc_hd__dfxtp_2 _18225_ (.CLK(clknet_leaf_29_clk),
    .D(_01296_),
    .Q(instr_waitirq));
 sky130_fd_sc_hd__dfxtp_4 _18226_ (.CLK(clknet_leaf_104_clk),
    .D(_01297_),
    .Q(instr_timer));
 sky130_fd_sc_hd__dfxtp_1 _18227_ (.CLK(clknet_leaf_32_clk),
    .D(_01298_),
    .Q(\decoded_rd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18228_ (.CLK(clknet_leaf_32_clk),
    .D(_01299_),
    .Q(\decoded_rd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18229_ (.CLK(clknet_leaf_23_clk),
    .D(_01300_),
    .Q(\decoded_rd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18230_ (.CLK(clknet_leaf_9_clk),
    .D(_01301_),
    .Q(\decoded_rd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18231_ (.CLK(clknet_leaf_16_clk),
    .D(_01302_),
    .Q(\decoded_rd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18232_ (.CLK(clknet_leaf_9_clk),
    .D(_01303_),
    .Q(\cpuregs.raddr1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18233_ (.CLK(clknet_leaf_9_clk),
    .D(_01304_),
    .Q(\cpuregs.raddr1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18234_ (.CLK(clknet_leaf_9_clk),
    .D(_01305_),
    .Q(\cpuregs.raddr1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18235_ (.CLK(clknet_leaf_9_clk),
    .D(_01306_),
    .Q(\cpuregs.raddr1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18236_ (.CLK(clknet_leaf_8_clk),
    .D(_01307_),
    .Q(\cpuregs.raddr1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18237_ (.CLK(clknet_leaf_23_clk),
    .D(_01308_),
    .Q(\cpuregs.raddr2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18238_ (.CLK(clknet_leaf_23_clk),
    .D(_01309_),
    .Q(\cpuregs.raddr2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18239_ (.CLK(clknet_leaf_23_clk),
    .D(_01310_),
    .Q(\cpuregs.raddr2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18240_ (.CLK(clknet_leaf_24_clk),
    .D(_01311_),
    .Q(\cpuregs.raddr2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18241_ (.CLK(clknet_leaf_16_clk),
    .D(_01312_),
    .Q(\cpuregs.raddr2[4] ));
 sky130_fd_sc_hd__dfxtp_2 _18242_ (.CLK(clknet_leaf_22_clk),
    .D(_01313_),
    .Q(\decoded_imm[0] ));
 sky130_fd_sc_hd__dfxtp_2 _18243_ (.CLK(clknet_leaf_22_clk),
    .D(_01314_),
    .Q(\decoded_imm[1] ));
 sky130_fd_sc_hd__dfxtp_2 _18244_ (.CLK(clknet_leaf_25_clk),
    .D(_01315_),
    .Q(\decoded_imm[2] ));
 sky130_fd_sc_hd__dfxtp_2 _18245_ (.CLK(clknet_leaf_25_clk),
    .D(_01316_),
    .Q(\decoded_imm[3] ));
 sky130_fd_sc_hd__dfxtp_2 _18246_ (.CLK(clknet_leaf_25_clk),
    .D(_01317_),
    .Q(\decoded_imm[4] ));
 sky130_fd_sc_hd__dfxtp_2 _18247_ (.CLK(clknet_leaf_23_clk),
    .D(_01318_),
    .Q(\decoded_imm[5] ));
 sky130_fd_sc_hd__dfxtp_2 _18248_ (.CLK(clknet_leaf_23_clk),
    .D(_01319_),
    .Q(\decoded_imm[6] ));
 sky130_fd_sc_hd__dfxtp_2 _18249_ (.CLK(clknet_leaf_23_clk),
    .D(_01320_),
    .Q(\decoded_imm[7] ));
 sky130_fd_sc_hd__dfxtp_4 _18250_ (.CLK(clknet_leaf_22_clk),
    .D(_01321_),
    .Q(\decoded_imm[8] ));
 sky130_fd_sc_hd__dfxtp_4 _18251_ (.CLK(clknet_leaf_22_clk),
    .D(_01322_),
    .Q(\decoded_imm[9] ));
 sky130_fd_sc_hd__dfxtp_4 _18252_ (.CLK(clknet_leaf_22_clk),
    .D(_01323_),
    .Q(\decoded_imm[10] ));
 sky130_fd_sc_hd__dfxtp_4 _18253_ (.CLK(clknet_leaf_24_clk),
    .D(_01324_),
    .Q(\decoded_imm[11] ));
 sky130_fd_sc_hd__dfxtp_4 _18254_ (.CLK(clknet_leaf_26_clk),
    .D(_01325_),
    .Q(\decoded_imm[12] ));
 sky130_fd_sc_hd__dfxtp_4 _18255_ (.CLK(clknet_leaf_26_clk),
    .D(_01326_),
    .Q(\decoded_imm[13] ));
 sky130_fd_sc_hd__dfxtp_4 _18256_ (.CLK(clknet_leaf_25_clk),
    .D(_01327_),
    .Q(\decoded_imm[14] ));
 sky130_fd_sc_hd__dfxtp_4 _18257_ (.CLK(clknet_leaf_31_clk),
    .D(_01328_),
    .Q(\decoded_imm[15] ));
 sky130_fd_sc_hd__dfxtp_4 _18258_ (.CLK(clknet_leaf_24_clk),
    .D(_01329_),
    .Q(\decoded_imm[16] ));
 sky130_fd_sc_hd__dfxtp_4 _18259_ (.CLK(clknet_leaf_28_clk),
    .D(_01330_),
    .Q(\decoded_imm[17] ));
 sky130_fd_sc_hd__dfxtp_4 _18260_ (.CLK(clknet_leaf_31_clk),
    .D(_01331_),
    .Q(\decoded_imm[18] ));
 sky130_fd_sc_hd__dfxtp_4 _18261_ (.CLK(clknet_leaf_29_clk),
    .D(_01332_),
    .Q(\decoded_imm[19] ));
 sky130_fd_sc_hd__dfxtp_4 _18262_ (.CLK(clknet_leaf_26_clk),
    .D(_01333_),
    .Q(\decoded_imm[20] ));
 sky130_fd_sc_hd__dfxtp_4 _18263_ (.CLK(clknet_leaf_26_clk),
    .D(_01334_),
    .Q(\decoded_imm[21] ));
 sky130_fd_sc_hd__dfxtp_4 _18264_ (.CLK(clknet_leaf_26_clk),
    .D(_01335_),
    .Q(\decoded_imm[22] ));
 sky130_fd_sc_hd__dfxtp_4 _18265_ (.CLK(clknet_leaf_25_clk),
    .D(_01336_),
    .Q(\decoded_imm[23] ));
 sky130_fd_sc_hd__dfxtp_4 _18266_ (.CLK(clknet_leaf_26_clk),
    .D(_01337_),
    .Q(\decoded_imm[24] ));
 sky130_fd_sc_hd__dfxtp_4 _18267_ (.CLK(clknet_leaf_26_clk),
    .D(_01338_),
    .Q(\decoded_imm[25] ));
 sky130_fd_sc_hd__dfxtp_4 _18268_ (.CLK(clknet_leaf_25_clk),
    .D(_01339_),
    .Q(\decoded_imm[26] ));
 sky130_fd_sc_hd__dfxtp_4 _18269_ (.CLK(clknet_leaf_26_clk),
    .D(_01340_),
    .Q(\decoded_imm[27] ));
 sky130_fd_sc_hd__dfxtp_4 _18270_ (.CLK(clknet_leaf_26_clk),
    .D(_01341_),
    .Q(\decoded_imm[28] ));
 sky130_fd_sc_hd__dfxtp_2 _18271_ (.CLK(clknet_leaf_25_clk),
    .D(_01342_),
    .Q(\decoded_imm[29] ));
 sky130_fd_sc_hd__dfxtp_4 _18272_ (.CLK(clknet_leaf_25_clk),
    .D(_01343_),
    .Q(\decoded_imm[30] ));
 sky130_fd_sc_hd__dfxtp_2 _18273_ (.CLK(clknet_leaf_25_clk),
    .D(_01344_),
    .Q(\decoded_imm[31] ));
 sky130_fd_sc_hd__dfxtp_1 _18274_ (.CLK(clknet_leaf_25_clk),
    .D(_00033_),
    .Q(is_lui_auipc_jal));
 sky130_fd_sc_hd__dfxtp_1 _18275_ (.CLK(clknet_leaf_23_clk),
    .D(_01345_),
    .Q(compressed_instr));
 sky130_fd_sc_hd__dfxtp_2 _18276_ (.CLK(clknet_leaf_29_clk),
    .D(_01346_),
    .Q(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__dfxtp_2 _18277_ (.CLK(clknet_leaf_28_clk),
    .D(_01347_),
    .Q(is_slli_srli_srai));
 sky130_fd_sc_hd__dfxtp_1 _18278_ (.CLK(clknet_leaf_29_clk),
    .D(_01348_),
    .Q(is_jalr_addi_slti_sltiu_xori_ori_andi));
 sky130_fd_sc_hd__dfxtp_4 _18279_ (.CLK(clknet_leaf_31_clk),
    .D(_01349_),
    .Q(is_sb_sh_sw));
 sky130_fd_sc_hd__dfxtp_1 _18280_ (.CLK(clknet_leaf_43_clk),
    .D(_00034_),
    .Q(is_slti_blt_slt));
 sky130_fd_sc_hd__dfxtp_1 _18281_ (.CLK(clknet_leaf_43_clk),
    .D(_00035_),
    .Q(is_sltiu_bltu_sltu));
 sky130_fd_sc_hd__dfxtp_1 _18282_ (.CLK(clknet_leaf_24_clk),
    .D(_01350_),
    .Q(is_beq_bne_blt_bge_bltu_bgeu));
 sky130_fd_sc_hd__dfxtp_2 _18283_ (.CLK(clknet_leaf_32_clk),
    .D(_01351_),
    .Q(is_alu_reg_imm));
 sky130_fd_sc_hd__dfxtp_1 _18284_ (.CLK(clknet_leaf_8_clk),
    .D(_01352_),
    .Q(is_alu_reg_reg));
 sky130_fd_sc_hd__dfxtp_1 _18285_ (.CLK(clknet_leaf_42_clk),
    .D(_01353_),
    .Q(is_compare));
 sky130_fd_sc_hd__dfxtp_2 _18286_ (.CLK(clknet_leaf_38_clk),
    .D(_01354_),
    .Q(net193));
 sky130_fd_sc_hd__dfxtp_1 _18287_ (.CLK(clknet_leaf_38_clk),
    .D(_01355_),
    .Q(\mem_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18288_ (.CLK(clknet_leaf_39_clk),
    .D(_01356_),
    .Q(\mem_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18289_ (.CLK(clknet_leaf_37_clk),
    .D(_01357_),
    .Q(net263));
 sky130_fd_sc_hd__dfxtp_1 _18290_ (.CLK(clknet_leaf_5_clk),
    .D(_01358_),
    .Q(net274));
 sky130_fd_sc_hd__dfxtp_1 _18291_ (.CLK(clknet_leaf_5_clk),
    .D(_01359_),
    .Q(net285));
 sky130_fd_sc_hd__dfxtp_1 _18292_ (.CLK(clknet_leaf_38_clk),
    .D(_01360_),
    .Q(net288));
 sky130_fd_sc_hd__dfxtp_1 _18293_ (.CLK(clknet_leaf_5_clk),
    .D(_01361_),
    .Q(net289));
 sky130_fd_sc_hd__dfxtp_1 _18294_ (.CLK(clknet_leaf_5_clk),
    .D(_01362_),
    .Q(net290));
 sky130_fd_sc_hd__dfxtp_1 _18295_ (.CLK(clknet_leaf_5_clk),
    .D(_01363_),
    .Q(net291));
 sky130_fd_sc_hd__dfxtp_1 _18296_ (.CLK(clknet_leaf_5_clk),
    .D(_01364_),
    .Q(net292));
 sky130_fd_sc_hd__dfxtp_1 _18297_ (.CLK(clknet_leaf_5_clk),
    .D(_01365_),
    .Q(net293));
 sky130_fd_sc_hd__dfxtp_1 _18298_ (.CLK(clknet_leaf_5_clk),
    .D(_01366_),
    .Q(net294));
 sky130_fd_sc_hd__dfxtp_1 _18299_ (.CLK(clknet_leaf_5_clk),
    .D(_01367_),
    .Q(net264));
 sky130_fd_sc_hd__dfxtp_1 _18300_ (.CLK(clknet_leaf_5_clk),
    .D(_01368_),
    .Q(net265));
 sky130_fd_sc_hd__dfxtp_1 _18301_ (.CLK(clknet_leaf_5_clk),
    .D(_01369_),
    .Q(net266));
 sky130_fd_sc_hd__dfxtp_1 _18302_ (.CLK(clknet_leaf_6_clk),
    .D(_01370_),
    .Q(net267));
 sky130_fd_sc_hd__dfxtp_1 _18303_ (.CLK(clknet_leaf_6_clk),
    .D(_01371_),
    .Q(net268));
 sky130_fd_sc_hd__dfxtp_1 _18304_ (.CLK(clknet_leaf_6_clk),
    .D(_01372_),
    .Q(net269));
 sky130_fd_sc_hd__dfxtp_1 _18305_ (.CLK(clknet_leaf_35_clk),
    .D(_01373_),
    .Q(net270));
 sky130_fd_sc_hd__dfxtp_1 _18306_ (.CLK(clknet_leaf_35_clk),
    .D(_01374_),
    .Q(net271));
 sky130_fd_sc_hd__dfxtp_1 _18307_ (.CLK(clknet_leaf_35_clk),
    .D(_01375_),
    .Q(net272));
 sky130_fd_sc_hd__dfxtp_1 _18308_ (.CLK(clknet_leaf_35_clk),
    .D(_01376_),
    .Q(net273));
 sky130_fd_sc_hd__dfxtp_1 _18309_ (.CLK(clknet_leaf_35_clk),
    .D(_01377_),
    .Q(net275));
 sky130_fd_sc_hd__dfxtp_1 _18310_ (.CLK(clknet_leaf_35_clk),
    .D(_01378_),
    .Q(net276));
 sky130_fd_sc_hd__dfxtp_1 _18311_ (.CLK(clknet_leaf_35_clk),
    .D(_01379_),
    .Q(net277));
 sky130_fd_sc_hd__dfxtp_1 _18312_ (.CLK(clknet_leaf_35_clk),
    .D(_01380_),
    .Q(net278));
 sky130_fd_sc_hd__dfxtp_1 _18313_ (.CLK(clknet_leaf_35_clk),
    .D(_01381_),
    .Q(net279));
 sky130_fd_sc_hd__dfxtp_1 _18314_ (.CLK(clknet_leaf_36_clk),
    .D(_01382_),
    .Q(net280));
 sky130_fd_sc_hd__dfxtp_1 _18315_ (.CLK(clknet_leaf_36_clk),
    .D(_01383_),
    .Q(net281));
 sky130_fd_sc_hd__dfxtp_1 _18316_ (.CLK(clknet_leaf_36_clk),
    .D(_01384_),
    .Q(net282));
 sky130_fd_sc_hd__dfxtp_1 _18317_ (.CLK(clknet_leaf_38_clk),
    .D(_01385_),
    .Q(net283));
 sky130_fd_sc_hd__dfxtp_1 _18318_ (.CLK(clknet_leaf_38_clk),
    .D(_01386_),
    .Q(net284));
 sky130_fd_sc_hd__dfxtp_1 _18319_ (.CLK(clknet_leaf_37_clk),
    .D(_01387_),
    .Q(net286));
 sky130_fd_sc_hd__dfxtp_1 _18320_ (.CLK(clknet_leaf_37_clk),
    .D(_01388_),
    .Q(net287));
 sky130_fd_sc_hd__dfxtp_1 _18321_ (.CLK(clknet_leaf_38_clk),
    .D(_01389_),
    .Q(net295));
 sky130_fd_sc_hd__dfxtp_1 _18322_ (.CLK(clknet_leaf_38_clk),
    .D(_01390_),
    .Q(net296));
 sky130_fd_sc_hd__dfxtp_1 _18323_ (.CLK(clknet_leaf_38_clk),
    .D(_01391_),
    .Q(net297));
 sky130_fd_sc_hd__dfxtp_1 _18324_ (.CLK(clknet_leaf_38_clk),
    .D(_01392_),
    .Q(net298));
 sky130_fd_sc_hd__dfxtp_1 _18325_ (.CLK(clknet_leaf_39_clk),
    .D(_01393_),
    .Q(mem_la_secondword));
 sky130_fd_sc_hd__dfxtp_1 _18326_ (.CLK(clknet_leaf_39_clk),
    .D(_01394_),
    .Q(prefetched_high_word));
 sky130_fd_sc_hd__dfxtp_1 _18327_ (.CLK(clknet_leaf_19_clk),
    .D(_01395_),
    .Q(\cpuregs.waddr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18328_ (.CLK(clknet_leaf_19_clk),
    .D(_01396_),
    .Q(\cpuregs.waddr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18329_ (.CLK(clknet_leaf_37_clk),
    .D(_01397_),
    .Q(\mem_16bit_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18330_ (.CLK(clknet_leaf_38_clk),
    .D(_01398_),
    .Q(\mem_16bit_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18331_ (.CLK(clknet_leaf_36_clk),
    .D(_01399_),
    .Q(\mem_16bit_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18332_ (.CLK(clknet_leaf_36_clk),
    .D(_01400_),
    .Q(\mem_16bit_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18333_ (.CLK(clknet_leaf_35_clk),
    .D(_01401_),
    .Q(\mem_16bit_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18334_ (.CLK(clknet_leaf_36_clk),
    .D(_01402_),
    .Q(\mem_16bit_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18335_ (.CLK(clknet_leaf_35_clk),
    .D(_01403_),
    .Q(\mem_16bit_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18336_ (.CLK(clknet_leaf_37_clk),
    .D(_01404_),
    .Q(\mem_16bit_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _18337_ (.CLK(clknet_leaf_35_clk),
    .D(_01405_),
    .Q(\mem_16bit_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _18338_ (.CLK(clknet_leaf_37_clk),
    .D(_01406_),
    .Q(\mem_16bit_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _18339_ (.CLK(clknet_leaf_37_clk),
    .D(_01407_),
    .Q(\mem_16bit_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _18340_ (.CLK(clknet_leaf_38_clk),
    .D(_01408_),
    .Q(\mem_16bit_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _18341_ (.CLK(clknet_leaf_36_clk),
    .D(_01409_),
    .Q(\mem_16bit_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _18342_ (.CLK(clknet_leaf_37_clk),
    .D(_01410_),
    .Q(\mem_16bit_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _18343_ (.CLK(clknet_leaf_37_clk),
    .D(_01411_),
    .Q(\mem_16bit_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _18344_ (.CLK(clknet_leaf_36_clk),
    .D(_01412_),
    .Q(\mem_16bit_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _18345_ (.CLK(clknet_leaf_29_clk),
    .D(_01413_),
    .Q(\mem_rdata_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18346_ (.CLK(clknet_leaf_30_clk),
    .D(_01414_),
    .Q(\mem_rdata_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18347_ (.CLK(clknet_leaf_35_clk),
    .D(_01415_),
    .Q(\mem_rdata_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18348_ (.CLK(clknet_leaf_30_clk),
    .D(_01416_),
    .Q(\mem_rdata_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18349_ (.CLK(clknet_leaf_33_clk),
    .D(_01417_),
    .Q(\mem_rdata_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18350_ (.CLK(clknet_leaf_35_clk),
    .D(_01418_),
    .Q(\mem_rdata_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18351_ (.CLK(clknet_leaf_36_clk),
    .D(_01419_),
    .Q(\mem_rdata_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18352_ (.CLK(clknet_leaf_40_clk),
    .D(_01420_),
    .Q(mem_la_firstword_reg));
 sky130_fd_sc_hd__dfxtp_2 _18353_ (.CLK(clknet_leaf_50_clk),
    .D(_01421_),
    .Q(\reg_next_pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18354_ (.CLK(clknet_leaf_53_clk),
    .D(_00061_),
    .Q(\reg_sh[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18355_ (.CLK(clknet_leaf_52_clk),
    .D(_00062_),
    .Q(\reg_sh[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18356_ (.CLK(clknet_leaf_52_clk),
    .D(_00063_),
    .Q(\reg_sh[4] ));
 sky130_fd_sc_hd__dfxtp_1 _18357_ (.CLK(clknet_leaf_17_clk),
    .D(_01422_),
    .Q(\cpuregs.regs[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18358_ (.CLK(clknet_leaf_189_clk),
    .D(_01423_),
    .Q(\cpuregs.regs[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18359_ (.CLK(clknet_leaf_10_clk),
    .D(_01424_),
    .Q(\cpuregs.regs[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18360_ (.CLK(clknet_leaf_10_clk),
    .D(_01425_),
    .Q(\cpuregs.regs[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18361_ (.CLK(clknet_leaf_187_clk),
    .D(_01426_),
    .Q(\cpuregs.regs[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18362_ (.CLK(clknet_leaf_18_clk),
    .D(_01427_),
    .Q(\cpuregs.regs[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18363_ (.CLK(clknet_leaf_179_clk),
    .D(_01428_),
    .Q(\cpuregs.regs[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18364_ (.CLK(clknet_leaf_174_clk),
    .D(_01429_),
    .Q(\cpuregs.regs[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18365_ (.CLK(clknet_leaf_185_clk),
    .D(_01430_),
    .Q(\cpuregs.regs[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18366_ (.CLK(clknet_leaf_185_clk),
    .D(_01431_),
    .Q(\cpuregs.regs[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18367_ (.CLK(clknet_leaf_127_clk),
    .D(_01432_),
    .Q(\cpuregs.regs[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18368_ (.CLK(clknet_leaf_160_clk),
    .D(_01433_),
    .Q(\cpuregs.regs[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18369_ (.CLK(clknet_leaf_149_clk),
    .D(_01434_),
    .Q(\cpuregs.regs[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18370_ (.CLK(clknet_leaf_138_clk),
    .D(_01435_),
    .Q(\cpuregs.regs[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18371_ (.CLK(clknet_leaf_146_clk),
    .D(_01436_),
    .Q(\cpuregs.regs[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18372_ (.CLK(clknet_leaf_129_clk),
    .D(_01437_),
    .Q(\cpuregs.regs[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18373_ (.CLK(clknet_leaf_141_clk),
    .D(_01438_),
    .Q(\cpuregs.regs[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18374_ (.CLK(clknet_leaf_139_clk),
    .D(_01439_),
    .Q(\cpuregs.regs[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18375_ (.CLK(clknet_leaf_154_clk),
    .D(_01440_),
    .Q(\cpuregs.regs[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18376_ (.CLK(clknet_leaf_180_clk),
    .D(_01441_),
    .Q(\cpuregs.regs[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18377_ (.CLK(clknet_leaf_99_clk),
    .D(_01442_),
    .Q(\cpuregs.regs[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18378_ (.CLK(clknet_leaf_98_clk),
    .D(_01443_),
    .Q(\cpuregs.regs[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18379_ (.CLK(clknet_leaf_118_clk),
    .D(_01444_),
    .Q(\cpuregs.regs[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18380_ (.CLK(clknet_leaf_163_clk),
    .D(_01445_),
    .Q(\cpuregs.regs[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18381_ (.CLK(clknet_leaf_164_clk),
    .D(_01446_),
    .Q(\cpuregs.regs[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18382_ (.CLK(clknet_leaf_111_clk),
    .D(_01447_),
    .Q(\cpuregs.regs[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18383_ (.CLK(clknet_leaf_166_clk),
    .D(_01448_),
    .Q(\cpuregs.regs[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18384_ (.CLK(clknet_leaf_106_clk),
    .D(_01449_),
    .Q(\cpuregs.regs[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18385_ (.CLK(clknet_leaf_113_clk),
    .D(_01450_),
    .Q(\cpuregs.regs[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18386_ (.CLK(clknet_leaf_128_clk),
    .D(_01451_),
    .Q(\cpuregs.regs[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18387_ (.CLK(clknet_leaf_163_clk),
    .D(_01452_),
    .Q(\cpuregs.regs[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18388_ (.CLK(clknet_leaf_168_clk),
    .D(_01453_),
    .Q(\cpuregs.regs[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18389_ (.CLK(clknet_leaf_14_clk),
    .D(_01454_),
    .Q(\cpuregs.regs[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18390_ (.CLK(clknet_leaf_189_clk),
    .D(_01455_),
    .Q(\cpuregs.regs[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18391_ (.CLK(clknet_leaf_12_clk),
    .D(_01456_),
    .Q(\cpuregs.regs[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18392_ (.CLK(clknet_leaf_3_clk),
    .D(_01457_),
    .Q(\cpuregs.regs[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18393_ (.CLK(clknet_leaf_1_clk),
    .D(_01458_),
    .Q(\cpuregs.regs[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18394_ (.CLK(clknet_leaf_170_clk),
    .D(_01459_),
    .Q(\cpuregs.regs[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18395_ (.CLK(clknet_leaf_181_clk),
    .D(_01460_),
    .Q(\cpuregs.regs[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18396_ (.CLK(clknet_leaf_173_clk),
    .D(_01461_),
    .Q(\cpuregs.regs[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18397_ (.CLK(clknet_leaf_183_clk),
    .D(_01462_),
    .Q(\cpuregs.regs[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18398_ (.CLK(clknet_leaf_179_clk),
    .D(_01463_),
    .Q(\cpuregs.regs[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18399_ (.CLK(clknet_leaf_132_clk),
    .D(_01464_),
    .Q(\cpuregs.regs[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18400_ (.CLK(clknet_leaf_159_clk),
    .D(_01465_),
    .Q(\cpuregs.regs[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18401_ (.CLK(clknet_leaf_157_clk),
    .D(_01466_),
    .Q(\cpuregs.regs[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18402_ (.CLK(clknet_leaf_137_clk),
    .D(_01467_),
    .Q(\cpuregs.regs[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18403_ (.CLK(clknet_leaf_147_clk),
    .D(_01468_),
    .Q(\cpuregs.regs[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18404_ (.CLK(clknet_leaf_143_clk),
    .D(_01469_),
    .Q(\cpuregs.regs[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18405_ (.CLK(clknet_leaf_138_clk),
    .D(_01470_),
    .Q(\cpuregs.regs[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18406_ (.CLK(clknet_leaf_140_clk),
    .D(_01471_),
    .Q(\cpuregs.regs[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18407_ (.CLK(clknet_leaf_156_clk),
    .D(_01472_),
    .Q(\cpuregs.regs[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18408_ (.CLK(clknet_leaf_149_clk),
    .D(_01473_),
    .Q(\cpuregs.regs[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18409_ (.CLK(clknet_leaf_99_clk),
    .D(_01474_),
    .Q(\cpuregs.regs[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18410_ (.CLK(clknet_leaf_123_clk),
    .D(_01475_),
    .Q(\cpuregs.regs[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18411_ (.CLK(clknet_leaf_124_clk),
    .D(_01476_),
    .Q(\cpuregs.regs[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18412_ (.CLK(clknet_leaf_109_clk),
    .D(_01477_),
    .Q(\cpuregs.regs[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18413_ (.CLK(clknet_leaf_161_clk),
    .D(_01478_),
    .Q(\cpuregs.regs[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18414_ (.CLK(clknet_leaf_107_clk),
    .D(_01479_),
    .Q(\cpuregs.regs[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18415_ (.CLK(clknet_leaf_109_clk),
    .D(_01480_),
    .Q(\cpuregs.regs[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18416_ (.CLK(clknet_leaf_108_clk),
    .D(_01481_),
    .Q(\cpuregs.regs[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18417_ (.CLK(clknet_leaf_117_clk),
    .D(_01482_),
    .Q(\cpuregs.regs[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18418_ (.CLK(clknet_leaf_127_clk),
    .D(_01483_),
    .Q(\cpuregs.regs[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18419_ (.CLK(clknet_leaf_162_clk),
    .D(_01484_),
    .Q(\cpuregs.regs[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18420_ (.CLK(clknet_leaf_176_clk),
    .D(_01485_),
    .Q(\cpuregs.regs[16][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18421_ (.CLK(clknet_leaf_15_clk),
    .D(_01486_),
    .Q(\cpuregs.regs[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18422_ (.CLK(clknet_leaf_188_clk),
    .D(_01487_),
    .Q(\cpuregs.regs[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18423_ (.CLK(clknet_leaf_14_clk),
    .D(_01488_),
    .Q(\cpuregs.regs[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18424_ (.CLK(clknet_leaf_12_clk),
    .D(_01489_),
    .Q(\cpuregs.regs[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18425_ (.CLK(clknet_leaf_187_clk),
    .D(_01490_),
    .Q(\cpuregs.regs[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18426_ (.CLK(clknet_leaf_166_clk),
    .D(_01491_),
    .Q(\cpuregs.regs[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18427_ (.CLK(clknet_leaf_181_clk),
    .D(_01492_),
    .Q(\cpuregs.regs[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18428_ (.CLK(clknet_leaf_175_clk),
    .D(_01493_),
    .Q(\cpuregs.regs[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18429_ (.CLK(clknet_leaf_184_clk),
    .D(_01494_),
    .Q(\cpuregs.regs[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18430_ (.CLK(clknet_leaf_183_clk),
    .D(_01495_),
    .Q(\cpuregs.regs[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18431_ (.CLK(clknet_leaf_133_clk),
    .D(_01496_),
    .Q(\cpuregs.regs[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18432_ (.CLK(clknet_leaf_143_clk),
    .D(_01497_),
    .Q(\cpuregs.regs[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18433_ (.CLK(clknet_leaf_147_clk),
    .D(_01498_),
    .Q(\cpuregs.regs[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18434_ (.CLK(clknet_leaf_137_clk),
    .D(_01499_),
    .Q(\cpuregs.regs[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18435_ (.CLK(clknet_leaf_145_clk),
    .D(_01500_),
    .Q(\cpuregs.regs[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18436_ (.CLK(clknet_leaf_133_clk),
    .D(_01501_),
    .Q(\cpuregs.regs[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18437_ (.CLK(clknet_leaf_135_clk),
    .D(_01502_),
    .Q(\cpuregs.regs[29][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18438_ (.CLK(clknet_leaf_147_clk),
    .D(_01503_),
    .Q(\cpuregs.regs[29][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18439_ (.CLK(clknet_leaf_151_clk),
    .D(_01504_),
    .Q(\cpuregs.regs[29][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18440_ (.CLK(clknet_leaf_151_clk),
    .D(_01505_),
    .Q(\cpuregs.regs[29][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18441_ (.CLK(clknet_leaf_98_clk),
    .D(_01506_),
    .Q(\cpuregs.regs[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18442_ (.CLK(clknet_leaf_97_clk),
    .D(_01507_),
    .Q(\cpuregs.regs[29][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18443_ (.CLK(clknet_leaf_122_clk),
    .D(_01508_),
    .Q(\cpuregs.regs[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18444_ (.CLK(clknet_leaf_164_clk),
    .D(_01509_),
    .Q(\cpuregs.regs[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18445_ (.CLK(clknet_leaf_160_clk),
    .D(_01510_),
    .Q(\cpuregs.regs[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18446_ (.CLK(clknet_leaf_112_clk),
    .D(_01511_),
    .Q(\cpuregs.regs[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18447_ (.CLK(clknet_leaf_165_clk),
    .D(_01512_),
    .Q(\cpuregs.regs[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18448_ (.CLK(clknet_leaf_113_clk),
    .D(_01513_),
    .Q(\cpuregs.regs[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18449_ (.CLK(clknet_leaf_115_clk),
    .D(_01514_),
    .Q(\cpuregs.regs[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18450_ (.CLK(clknet_leaf_125_clk),
    .D(_01515_),
    .Q(\cpuregs.regs[29][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18451_ (.CLK(clknet_leaf_155_clk),
    .D(_01516_),
    .Q(\cpuregs.regs[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18452_ (.CLK(clknet_leaf_177_clk),
    .D(_01517_),
    .Q(\cpuregs.regs[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18453_ (.CLK(clknet_leaf_14_clk),
    .D(_01518_),
    .Q(\cpuregs.regs[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18454_ (.CLK(clknet_leaf_189_clk),
    .D(_01519_),
    .Q(\cpuregs.regs[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18455_ (.CLK(clknet_leaf_12_clk),
    .D(_01520_),
    .Q(\cpuregs.regs[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18456_ (.CLK(clknet_leaf_11_clk),
    .D(_01521_),
    .Q(\cpuregs.regs[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18457_ (.CLK(clknet_leaf_1_clk),
    .D(_01522_),
    .Q(\cpuregs.regs[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18458_ (.CLK(clknet_leaf_171_clk),
    .D(_01523_),
    .Q(\cpuregs.regs[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18459_ (.CLK(clknet_leaf_181_clk),
    .D(_01524_),
    .Q(\cpuregs.regs[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18460_ (.CLK(clknet_leaf_173_clk),
    .D(_01525_),
    .Q(\cpuregs.regs[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18461_ (.CLK(clknet_leaf_184_clk),
    .D(_01526_),
    .Q(\cpuregs.regs[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18462_ (.CLK(clknet_leaf_182_clk),
    .D(_01527_),
    .Q(\cpuregs.regs[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18463_ (.CLK(clknet_leaf_132_clk),
    .D(_01528_),
    .Q(\cpuregs.regs[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18464_ (.CLK(clknet_leaf_158_clk),
    .D(_01529_),
    .Q(\cpuregs.regs[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18465_ (.CLK(clknet_leaf_157_clk),
    .D(_01530_),
    .Q(\cpuregs.regs[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18466_ (.CLK(clknet_leaf_137_clk),
    .D(_01531_),
    .Q(\cpuregs.regs[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18467_ (.CLK(clknet_leaf_148_clk),
    .D(_01532_),
    .Q(\cpuregs.regs[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18468_ (.CLK(clknet_leaf_143_clk),
    .D(_01533_),
    .Q(\cpuregs.regs[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18469_ (.CLK(clknet_leaf_132_clk),
    .D(_01534_),
    .Q(\cpuregs.regs[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18470_ (.CLK(clknet_leaf_140_clk),
    .D(_01535_),
    .Q(\cpuregs.regs[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18471_ (.CLK(clknet_leaf_156_clk),
    .D(_01536_),
    .Q(\cpuregs.regs[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18472_ (.CLK(clknet_leaf_149_clk),
    .D(_01537_),
    .Q(\cpuregs.regs[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18473_ (.CLK(clknet_leaf_121_clk),
    .D(_01538_),
    .Q(\cpuregs.regs[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18474_ (.CLK(clknet_leaf_123_clk),
    .D(_01539_),
    .Q(\cpuregs.regs[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18475_ (.CLK(clknet_leaf_124_clk),
    .D(_01540_),
    .Q(\cpuregs.regs[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18476_ (.CLK(clknet_leaf_109_clk),
    .D(_01541_),
    .Q(\cpuregs.regs[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18477_ (.CLK(clknet_leaf_161_clk),
    .D(_01542_),
    .Q(\cpuregs.regs[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18478_ (.CLK(clknet_leaf_106_clk),
    .D(_01543_),
    .Q(\cpuregs.regs[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18479_ (.CLK(clknet_leaf_20_clk),
    .D(_01544_),
    .Q(\cpuregs.regs[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18480_ (.CLK(clknet_leaf_108_clk),
    .D(_01545_),
    .Q(\cpuregs.regs[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18481_ (.CLK(clknet_leaf_116_clk),
    .D(_01546_),
    .Q(\cpuregs.regs[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18482_ (.CLK(clknet_leaf_128_clk),
    .D(_01547_),
    .Q(\cpuregs.regs[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18483_ (.CLK(clknet_leaf_155_clk),
    .D(_01548_),
    .Q(\cpuregs.regs[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18484_ (.CLK(clknet_leaf_170_clk),
    .D(_01549_),
    .Q(\cpuregs.regs[17][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18485_ (.CLK(clknet_leaf_14_clk),
    .D(_01550_),
    .Q(\cpuregs.regs[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18486_ (.CLK(clknet_leaf_189_clk),
    .D(_01551_),
    .Q(\cpuregs.regs[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18487_ (.CLK(clknet_leaf_11_clk),
    .D(_01552_),
    .Q(\cpuregs.regs[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18488_ (.CLK(clknet_leaf_3_clk),
    .D(_01553_),
    .Q(\cpuregs.regs[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18489_ (.CLK(clknet_leaf_1_clk),
    .D(_01554_),
    .Q(\cpuregs.regs[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18490_ (.CLK(clknet_leaf_171_clk),
    .D(_01555_),
    .Q(\cpuregs.regs[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18491_ (.CLK(clknet_leaf_181_clk),
    .D(_01556_),
    .Q(\cpuregs.regs[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18492_ (.CLK(clknet_leaf_186_clk),
    .D(_01557_),
    .Q(\cpuregs.regs[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18493_ (.CLK(clknet_leaf_184_clk),
    .D(_01558_),
    .Q(\cpuregs.regs[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18494_ (.CLK(clknet_leaf_182_clk),
    .D(_01559_),
    .Q(\cpuregs.regs[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18495_ (.CLK(clknet_leaf_131_clk),
    .D(_01560_),
    .Q(\cpuregs.regs[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18496_ (.CLK(clknet_leaf_157_clk),
    .D(_01561_),
    .Q(\cpuregs.regs[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18497_ (.CLK(clknet_leaf_156_clk),
    .D(_01562_),
    .Q(\cpuregs.regs[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18498_ (.CLK(clknet_leaf_138_clk),
    .D(_01563_),
    .Q(\cpuregs.regs[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18499_ (.CLK(clknet_leaf_148_clk),
    .D(_01564_),
    .Q(\cpuregs.regs[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18500_ (.CLK(clknet_leaf_143_clk),
    .D(_01565_),
    .Q(\cpuregs.regs[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18501_ (.CLK(clknet_leaf_138_clk),
    .D(_01566_),
    .Q(\cpuregs.regs[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18502_ (.CLK(clknet_leaf_146_clk),
    .D(_01567_),
    .Q(\cpuregs.regs[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18503_ (.CLK(clknet_leaf_154_clk),
    .D(_01568_),
    .Q(\cpuregs.regs[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18504_ (.CLK(clknet_leaf_151_clk),
    .D(_01569_),
    .Q(\cpuregs.regs[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18505_ (.CLK(clknet_leaf_99_clk),
    .D(_01570_),
    .Q(\cpuregs.regs[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18506_ (.CLK(clknet_leaf_121_clk),
    .D(_01571_),
    .Q(\cpuregs.regs[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18507_ (.CLK(clknet_leaf_122_clk),
    .D(_01572_),
    .Q(\cpuregs.regs[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18508_ (.CLK(clknet_leaf_109_clk),
    .D(_01573_),
    .Q(\cpuregs.regs[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18509_ (.CLK(clknet_leaf_162_clk),
    .D(_01574_),
    .Q(\cpuregs.regs[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18510_ (.CLK(clknet_leaf_107_clk),
    .D(_01575_),
    .Q(\cpuregs.regs[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18511_ (.CLK(clknet_leaf_20_clk),
    .D(_01576_),
    .Q(\cpuregs.regs[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18512_ (.CLK(clknet_leaf_108_clk),
    .D(_01577_),
    .Q(\cpuregs.regs[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18513_ (.CLK(clknet_leaf_116_clk),
    .D(_01578_),
    .Q(\cpuregs.regs[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18514_ (.CLK(clknet_leaf_128_clk),
    .D(_01579_),
    .Q(\cpuregs.regs[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18515_ (.CLK(clknet_leaf_155_clk),
    .D(_01580_),
    .Q(\cpuregs.regs[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18516_ (.CLK(clknet_leaf_174_clk),
    .D(_01581_),
    .Q(\cpuregs.regs[18][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18517_ (.CLK(clknet_leaf_17_clk),
    .D(_01582_),
    .Q(\cpuregs.regs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18518_ (.CLK(clknet_leaf_188_clk),
    .D(_01583_),
    .Q(\cpuregs.regs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18519_ (.CLK(clknet_leaf_17_clk),
    .D(_01584_),
    .Q(\cpuregs.regs[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18520_ (.CLK(clknet_leaf_8_clk),
    .D(_01585_),
    .Q(\cpuregs.regs[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18521_ (.CLK(clknet_leaf_2_clk),
    .D(_01586_),
    .Q(\cpuregs.regs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18522_ (.CLK(clknet_leaf_19_clk),
    .D(_01587_),
    .Q(\cpuregs.regs[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18523_ (.CLK(clknet_leaf_178_clk),
    .D(_01588_),
    .Q(\cpuregs.regs[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18524_ (.CLK(clknet_leaf_172_clk),
    .D(_01589_),
    .Q(\cpuregs.regs[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18525_ (.CLK(clknet_leaf_186_clk),
    .D(_01590_),
    .Q(\cpuregs.regs[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18526_ (.CLK(clknet_leaf_175_clk),
    .D(_01591_),
    .Q(\cpuregs.regs[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18527_ (.CLK(clknet_leaf_126_clk),
    .D(_01592_),
    .Q(\cpuregs.regs[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18528_ (.CLK(clknet_leaf_160_clk),
    .D(_01593_),
    .Q(\cpuregs.regs[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18529_ (.CLK(clknet_leaf_157_clk),
    .D(_01594_),
    .Q(\cpuregs.regs[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18530_ (.CLK(clknet_leaf_135_clk),
    .D(_01595_),
    .Q(\cpuregs.regs[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18531_ (.CLK(clknet_leaf_157_clk),
    .D(_01596_),
    .Q(\cpuregs.regs[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18532_ (.CLK(clknet_leaf_116_clk),
    .D(_01597_),
    .Q(\cpuregs.regs[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18533_ (.CLK(clknet_leaf_135_clk),
    .D(_01598_),
    .Q(\cpuregs.regs[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18534_ (.CLK(clknet_leaf_144_clk),
    .D(_01599_),
    .Q(\cpuregs.regs[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18535_ (.CLK(clknet_leaf_156_clk),
    .D(_01600_),
    .Q(\cpuregs.regs[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18536_ (.CLK(clknet_leaf_152_clk),
    .D(_01601_),
    .Q(\cpuregs.regs[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18537_ (.CLK(clknet_leaf_105_clk),
    .D(_01602_),
    .Q(\cpuregs.regs[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18538_ (.CLK(clknet_leaf_98_clk),
    .D(_01603_),
    .Q(\cpuregs.regs[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18539_ (.CLK(clknet_leaf_119_clk),
    .D(_01604_),
    .Q(\cpuregs.regs[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18540_ (.CLK(clknet_leaf_164_clk),
    .D(_01605_),
    .Q(\cpuregs.regs[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18541_ (.CLK(clknet_leaf_114_clk),
    .D(_01606_),
    .Q(\cpuregs.regs[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18542_ (.CLK(clknet_leaf_110_clk),
    .D(_01607_),
    .Q(\cpuregs.regs[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18543_ (.CLK(clknet_leaf_58_clk),
    .D(_01608_),
    .Q(\cpuregs.regs[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18544_ (.CLK(clknet_leaf_105_clk),
    .D(_01609_),
    .Q(\cpuregs.regs[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18545_ (.CLK(clknet_leaf_113_clk),
    .D(_01610_),
    .Q(\cpuregs.regs[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18546_ (.CLK(clknet_leaf_117_clk),
    .D(_01611_),
    .Q(\cpuregs.regs[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18547_ (.CLK(clknet_leaf_162_clk),
    .D(_01612_),
    .Q(\cpuregs.regs[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18548_ (.CLK(clknet_leaf_170_clk),
    .D(_01613_),
    .Q(\cpuregs.regs[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18549_ (.CLK(clknet_leaf_14_clk),
    .D(_01614_),
    .Q(\cpuregs.regs[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18550_ (.CLK(clknet_leaf_189_clk),
    .D(_01615_),
    .Q(\cpuregs.regs[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18551_ (.CLK(clknet_leaf_11_clk),
    .D(_01616_),
    .Q(\cpuregs.regs[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18552_ (.CLK(clknet_leaf_3_clk),
    .D(_01617_),
    .Q(\cpuregs.regs[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18553_ (.CLK(clknet_leaf_1_clk),
    .D(_01618_),
    .Q(\cpuregs.regs[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18554_ (.CLK(clknet_leaf_171_clk),
    .D(_01619_),
    .Q(\cpuregs.regs[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18555_ (.CLK(clknet_leaf_182_clk),
    .D(_01620_),
    .Q(\cpuregs.regs[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18556_ (.CLK(clknet_leaf_187_clk),
    .D(_01621_),
    .Q(\cpuregs.regs[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18557_ (.CLK(clknet_leaf_184_clk),
    .D(_01622_),
    .Q(\cpuregs.regs[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18558_ (.CLK(clknet_leaf_182_clk),
    .D(_01623_),
    .Q(\cpuregs.regs[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18559_ (.CLK(clknet_leaf_131_clk),
    .D(_01624_),
    .Q(\cpuregs.regs[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18560_ (.CLK(clknet_leaf_157_clk),
    .D(_01625_),
    .Q(\cpuregs.regs[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18561_ (.CLK(clknet_leaf_156_clk),
    .D(_01626_),
    .Q(\cpuregs.regs[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18562_ (.CLK(clknet_leaf_138_clk),
    .D(_01627_),
    .Q(\cpuregs.regs[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18563_ (.CLK(clknet_leaf_145_clk),
    .D(_01628_),
    .Q(\cpuregs.regs[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18564_ (.CLK(clknet_leaf_143_clk),
    .D(_01629_),
    .Q(\cpuregs.regs[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18565_ (.CLK(clknet_leaf_138_clk),
    .D(_01630_),
    .Q(\cpuregs.regs[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18566_ (.CLK(clknet_leaf_146_clk),
    .D(_01631_),
    .Q(\cpuregs.regs[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18567_ (.CLK(clknet_leaf_154_clk),
    .D(_01632_),
    .Q(\cpuregs.regs[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18568_ (.CLK(clknet_leaf_151_clk),
    .D(_01633_),
    .Q(\cpuregs.regs[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18569_ (.CLK(clknet_leaf_99_clk),
    .D(_01634_),
    .Q(\cpuregs.regs[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18570_ (.CLK(clknet_leaf_122_clk),
    .D(_01635_),
    .Q(\cpuregs.regs[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18571_ (.CLK(clknet_leaf_122_clk),
    .D(_01636_),
    .Q(\cpuregs.regs[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18572_ (.CLK(clknet_leaf_110_clk),
    .D(_01637_),
    .Q(\cpuregs.regs[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18573_ (.CLK(clknet_leaf_161_clk),
    .D(_01638_),
    .Q(\cpuregs.regs[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18574_ (.CLK(clknet_leaf_107_clk),
    .D(_01639_),
    .Q(\cpuregs.regs[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18575_ (.CLK(clknet_leaf_20_clk),
    .D(_01640_),
    .Q(\cpuregs.regs[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18576_ (.CLK(clknet_leaf_108_clk),
    .D(_01641_),
    .Q(\cpuregs.regs[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18577_ (.CLK(clknet_leaf_119_clk),
    .D(_01642_),
    .Q(\cpuregs.regs[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18578_ (.CLK(clknet_leaf_128_clk),
    .D(_01643_),
    .Q(\cpuregs.regs[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18579_ (.CLK(clknet_leaf_155_clk),
    .D(_01644_),
    .Q(\cpuregs.regs[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18580_ (.CLK(clknet_leaf_174_clk),
    .D(_01645_),
    .Q(\cpuregs.regs[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 _18581_ (.CLK(clknet_leaf_52_clk),
    .D(_01646_),
    .Q(\reg_sh[0] ));
 sky130_fd_sc_hd__dfxtp_1 _18582_ (.CLK(clknet_leaf_52_clk),
    .D(_01647_),
    .Q(\reg_sh[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18583_ (.CLK(clknet_leaf_17_clk),
    .D(_01648_),
    .Q(\cpuregs.regs[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18584_ (.CLK(clknet_leaf_189_clk),
    .D(_01649_),
    .Q(\cpuregs.regs[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18585_ (.CLK(clknet_leaf_10_clk),
    .D(_01650_),
    .Q(\cpuregs.regs[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18586_ (.CLK(clknet_leaf_10_clk),
    .D(_01651_),
    .Q(\cpuregs.regs[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18587_ (.CLK(clknet_leaf_187_clk),
    .D(_01652_),
    .Q(\cpuregs.regs[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18588_ (.CLK(clknet_leaf_166_clk),
    .D(_01653_),
    .Q(\cpuregs.regs[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18589_ (.CLK(clknet_leaf_180_clk),
    .D(_01654_),
    .Q(\cpuregs.regs[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18590_ (.CLK(clknet_leaf_173_clk),
    .D(_01655_),
    .Q(\cpuregs.regs[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18591_ (.CLK(clknet_leaf_185_clk),
    .D(_01656_),
    .Q(\cpuregs.regs[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18592_ (.CLK(clknet_leaf_182_clk),
    .D(_01657_),
    .Q(\cpuregs.regs[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18593_ (.CLK(clknet_leaf_129_clk),
    .D(_01658_),
    .Q(\cpuregs.regs[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18594_ (.CLK(clknet_leaf_159_clk),
    .D(_01659_),
    .Q(\cpuregs.regs[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18595_ (.CLK(clknet_leaf_149_clk),
    .D(_01660_),
    .Q(\cpuregs.regs[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18596_ (.CLK(clknet_leaf_138_clk),
    .D(_01661_),
    .Q(\cpuregs.regs[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18597_ (.CLK(clknet_leaf_146_clk),
    .D(_01662_),
    .Q(\cpuregs.regs[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18598_ (.CLK(clknet_leaf_129_clk),
    .D(_01663_),
    .Q(\cpuregs.regs[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18599_ (.CLK(clknet_leaf_131_clk),
    .D(_01664_),
    .Q(\cpuregs.regs[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18600_ (.CLK(clknet_leaf_138_clk),
    .D(_01665_),
    .Q(\cpuregs.regs[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18601_ (.CLK(clknet_leaf_177_clk),
    .D(_01666_),
    .Q(\cpuregs.regs[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18602_ (.CLK(clknet_leaf_151_clk),
    .D(_01667_),
    .Q(\cpuregs.regs[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18603_ (.CLK(clknet_leaf_99_clk),
    .D(_01668_),
    .Q(\cpuregs.regs[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18604_ (.CLK(clknet_leaf_99_clk),
    .D(_01669_),
    .Q(\cpuregs.regs[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18605_ (.CLK(clknet_leaf_121_clk),
    .D(_01670_),
    .Q(\cpuregs.regs[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18606_ (.CLK(clknet_leaf_163_clk),
    .D(_01671_),
    .Q(\cpuregs.regs[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18607_ (.CLK(clknet_leaf_164_clk),
    .D(_01672_),
    .Q(\cpuregs.regs[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18608_ (.CLK(clknet_leaf_111_clk),
    .D(_01673_),
    .Q(\cpuregs.regs[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18609_ (.CLK(clknet_leaf_165_clk),
    .D(_01674_),
    .Q(\cpuregs.regs[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18610_ (.CLK(clknet_leaf_106_clk),
    .D(_01675_),
    .Q(\cpuregs.regs[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18611_ (.CLK(clknet_leaf_113_clk),
    .D(_01676_),
    .Q(\cpuregs.regs[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18612_ (.CLK(clknet_leaf_117_clk),
    .D(_01677_),
    .Q(\cpuregs.regs[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18613_ (.CLK(clknet_leaf_163_clk),
    .D(_01678_),
    .Q(\cpuregs.regs[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18614_ (.CLK(clknet_leaf_167_clk),
    .D(_01679_),
    .Q(\cpuregs.regs[13][31] ));
 sky130_fd_sc_hd__dfxtp_2 _18615_ (.CLK(clknet_leaf_9_clk),
    .D(_00089_),
    .Q(_00069_));
 sky130_fd_sc_hd__dfxtp_1 _18616_ (.CLK(clknet_leaf_9_clk),
    .D(_00090_),
    .Q(_00070_));
 sky130_fd_sc_hd__dfxtp_4 _18617_ (.CLK(clknet_leaf_16_clk),
    .D(_00091_),
    .Q(_00071_));
 sky130_fd_sc_hd__dfxtp_1 _18618_ (.CLK(clknet_leaf_9_clk),
    .D(_00092_),
    .Q(_00072_));
 sky130_fd_sc_hd__dfxtp_4 _18619_ (.CLK(clknet_leaf_16_clk),
    .D(_00093_),
    .Q(_00073_));
 sky130_fd_sc_hd__dfxtp_1 _18620_ (.CLK(clknet_leaf_17_clk),
    .D(_01680_),
    .Q(\cpuregs.regs[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _18621_ (.CLK(clknet_leaf_189_clk),
    .D(_01681_),
    .Q(\cpuregs.regs[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _18622_ (.CLK(clknet_leaf_10_clk),
    .D(_01682_),
    .Q(\cpuregs.regs[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _18623_ (.CLK(clknet_leaf_10_clk),
    .D(_01683_),
    .Q(\cpuregs.regs[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _18624_ (.CLK(clknet_leaf_1_clk),
    .D(_01684_),
    .Q(\cpuregs.regs[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _18625_ (.CLK(clknet_leaf_18_clk),
    .D(_01685_),
    .Q(\cpuregs.regs[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _18626_ (.CLK(clknet_leaf_179_clk),
    .D(_01686_),
    .Q(\cpuregs.regs[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _18627_ (.CLK(clknet_leaf_174_clk),
    .D(_01687_),
    .Q(\cpuregs.regs[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _18628_ (.CLK(clknet_leaf_184_clk),
    .D(_01688_),
    .Q(\cpuregs.regs[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _18629_ (.CLK(clknet_leaf_182_clk),
    .D(_01689_),
    .Q(\cpuregs.regs[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _18630_ (.CLK(clknet_leaf_129_clk),
    .D(_01690_),
    .Q(\cpuregs.regs[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _18631_ (.CLK(clknet_leaf_160_clk),
    .D(_01691_),
    .Q(\cpuregs.regs[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _18632_ (.CLK(clknet_leaf_149_clk),
    .D(_01692_),
    .Q(\cpuregs.regs[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _18633_ (.CLK(clknet_leaf_138_clk),
    .D(_01693_),
    .Q(\cpuregs.regs[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _18634_ (.CLK(clknet_leaf_146_clk),
    .D(_01694_),
    .Q(\cpuregs.regs[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _18635_ (.CLK(clknet_leaf_129_clk),
    .D(_01695_),
    .Q(\cpuregs.regs[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _18636_ (.CLK(clknet_leaf_131_clk),
    .D(_01696_),
    .Q(\cpuregs.regs[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _18637_ (.CLK(clknet_leaf_140_clk),
    .D(_01697_),
    .Q(\cpuregs.regs[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _18638_ (.CLK(clknet_leaf_178_clk),
    .D(_01698_),
    .Q(\cpuregs.regs[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _18639_ (.CLK(clknet_leaf_180_clk),
    .D(_01699_),
    .Q(\cpuregs.regs[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _18640_ (.CLK(clknet_leaf_99_clk),
    .D(_01700_),
    .Q(\cpuregs.regs[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _18641_ (.CLK(clknet_leaf_99_clk),
    .D(_01701_),
    .Q(\cpuregs.regs[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _18642_ (.CLK(clknet_leaf_119_clk),
    .D(_01702_),
    .Q(\cpuregs.regs[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _18643_ (.CLK(clknet_leaf_163_clk),
    .D(_01703_),
    .Q(\cpuregs.regs[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _18644_ (.CLK(clknet_leaf_164_clk),
    .D(_01704_),
    .Q(\cpuregs.regs[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _18645_ (.CLK(clknet_leaf_111_clk),
    .D(_01705_),
    .Q(\cpuregs.regs[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _18646_ (.CLK(clknet_leaf_168_clk),
    .D(_01706_),
    .Q(\cpuregs.regs[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _18647_ (.CLK(clknet_leaf_112_clk),
    .D(_01707_),
    .Q(\cpuregs.regs[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _18648_ (.CLK(clknet_leaf_113_clk),
    .D(_01708_),
    .Q(\cpuregs.regs[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _18649_ (.CLK(clknet_leaf_117_clk),
    .D(_01709_),
    .Q(\cpuregs.regs[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _18650_ (.CLK(clknet_leaf_163_clk),
    .D(_01710_),
    .Q(\cpuregs.regs[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _18651_ (.CLK(clknet_leaf_167_clk),
    .D(_01711_),
    .Q(\cpuregs.regs[14][31] ));
 sky130_fd_sc_hd__conb_1 alphacore_303 (.LO(net303));
 sky130_fd_sc_hd__conb_1 alphacore_304 (.LO(net304));
 sky130_fd_sc_hd__conb_1 alphacore_305 (.LO(net305));
 sky130_fd_sc_hd__conb_1 alphacore_306 (.LO(net306));
 sky130_fd_sc_hd__conb_1 alphacore_307 (.LO(net307));
 sky130_fd_sc_hd__conb_1 alphacore_308 (.LO(net308));
 sky130_fd_sc_hd__conb_1 alphacore_309 (.LO(net309));
 sky130_fd_sc_hd__conb_1 alphacore_310 (.LO(net310));
 sky130_fd_sc_hd__conb_1 alphacore_311 (.LO(net311));
 sky130_fd_sc_hd__conb_1 alphacore_312 (.LO(net312));
 sky130_fd_sc_hd__conb_1 alphacore_313 (.LO(net313));
 sky130_fd_sc_hd__conb_1 alphacore_314 (.LO(net314));
 sky130_fd_sc_hd__conb_1 alphacore_315 (.LO(net315));
 sky130_fd_sc_hd__conb_1 alphacore_316 (.LO(net316));
 sky130_fd_sc_hd__conb_1 alphacore_317 (.LO(net317));
 sky130_fd_sc_hd__conb_1 alphacore_318 (.LO(net318));
 sky130_fd_sc_hd__conb_1 alphacore_319 (.LO(net319));
 sky130_fd_sc_hd__conb_1 alphacore_320 (.LO(net320));
 sky130_fd_sc_hd__conb_1 alphacore_321 (.LO(net321));
 sky130_fd_sc_hd__conb_1 alphacore_322 (.LO(net322));
 sky130_fd_sc_hd__conb_1 alphacore_323 (.LO(net323));
 sky130_fd_sc_hd__conb_1 alphacore_324 (.LO(net324));
 sky130_fd_sc_hd__conb_1 alphacore_325 (.LO(net325));
 sky130_fd_sc_hd__conb_1 alphacore_326 (.LO(net326));
 sky130_fd_sc_hd__conb_1 alphacore_327 (.LO(net327));
 sky130_fd_sc_hd__conb_1 alphacore_328 (.LO(net328));
 sky130_fd_sc_hd__conb_1 alphacore_329 (.LO(net329));
 sky130_fd_sc_hd__conb_1 alphacore_330 (.LO(net330));
 sky130_fd_sc_hd__conb_1 alphacore_331 (.LO(net331));
 sky130_fd_sc_hd__conb_1 alphacore_332 (.LO(net332));
 sky130_fd_sc_hd__conb_1 alphacore_333 (.LO(net333));
 sky130_fd_sc_hd__conb_1 alphacore_334 (.LO(net334));
 sky130_fd_sc_hd__conb_1 alphacore_335 (.LO(net335));
 sky130_fd_sc_hd__conb_1 alphacore_336 (.LO(net336));
 sky130_fd_sc_hd__conb_1 alphacore_337 (.LO(net337));
 sky130_fd_sc_hd__conb_1 alphacore_338 (.LO(net338));
 sky130_fd_sc_hd__conb_1 alphacore_339 (.LO(net339));
 sky130_fd_sc_hd__conb_1 alphacore_340 (.LO(net340));
 sky130_fd_sc_hd__conb_1 alphacore_341 (.LO(net341));
 sky130_fd_sc_hd__conb_1 alphacore_342 (.LO(net342));
 sky130_fd_sc_hd__conb_1 alphacore_343 (.LO(net343));
 sky130_fd_sc_hd__conb_1 alphacore_344 (.LO(net344));
 sky130_fd_sc_hd__conb_1 alphacore_345 (.LO(net345));
 sky130_fd_sc_hd__conb_1 alphacore_346 (.LO(net346));
 sky130_fd_sc_hd__conb_1 alphacore_347 (.LO(net347));
 sky130_fd_sc_hd__conb_1 alphacore_348 (.LO(net348));
 sky130_fd_sc_hd__conb_1 alphacore_349 (.LO(net349));
 sky130_fd_sc_hd__conb_1 alphacore_350 (.LO(net350));
 sky130_fd_sc_hd__conb_1 alphacore_351 (.LO(net351));
 sky130_fd_sc_hd__conb_1 alphacore_352 (.LO(net352));
 sky130_fd_sc_hd__conb_1 alphacore_353 (.LO(net353));
 sky130_fd_sc_hd__conb_1 alphacore_354 (.LO(net354));
 sky130_fd_sc_hd__conb_1 alphacore_355 (.LO(net355));
 sky130_fd_sc_hd__conb_1 alphacore_356 (.LO(net356));
 sky130_fd_sc_hd__conb_1 alphacore_357 (.LO(net357));
 sky130_fd_sc_hd__conb_1 alphacore_358 (.LO(net358));
 sky130_fd_sc_hd__conb_1 alphacore_359 (.LO(net359));
 sky130_fd_sc_hd__conb_1 alphacore_360 (.LO(net360));
 sky130_fd_sc_hd__conb_1 alphacore_361 (.LO(net361));
 sky130_fd_sc_hd__conb_1 alphacore_362 (.LO(net362));
 sky130_fd_sc_hd__conb_1 alphacore_363 (.LO(net363));
 sky130_fd_sc_hd__conb_1 alphacore_364 (.LO(net364));
 sky130_fd_sc_hd__conb_1 alphacore_365 (.LO(net365));
 sky130_fd_sc_hd__conb_1 alphacore_366 (.LO(net366));
 sky130_fd_sc_hd__conb_1 alphacore_367 (.LO(net367));
 sky130_fd_sc_hd__conb_1 alphacore_368 (.LO(net368));
 sky130_fd_sc_hd__conb_1 alphacore_369 (.LO(net369));
 sky130_fd_sc_hd__conb_1 alphacore_370 (.LO(net370));
 sky130_fd_sc_hd__conb_1 alphacore_371 (.LO(net371));
 sky130_fd_sc_hd__conb_1 alphacore_372 (.LO(net372));
 sky130_fd_sc_hd__conb_1 alphacore_373 (.LO(net373));
 sky130_fd_sc_hd__conb_1 alphacore_374 (.LO(net374));
 sky130_fd_sc_hd__conb_1 alphacore_375 (.LO(net375));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_1 _18726_ (.A(net99),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 _18727_ (.A(net110),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 _18728_ (.A(net121),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 _18729_ (.A(net124),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 _18730_ (.A(net125),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 _18731_ (.A(net126),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 _18732_ (.A(net127),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 _18733_ (.A(net128),
    .X(net254));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3515 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(irq[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(irq[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(irq[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(irq[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(irq[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(irq[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(irq[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(irq[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(irq[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(irq[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(irq[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(irq[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(irq[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(irq[21]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(irq[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(irq[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(irq[24]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(irq[25]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(irq[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(irq[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(irq[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(irq[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(irq[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(irq[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(irq[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input26 (.A(irq[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(irq[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(irq[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input29 (.A(irq[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input30 (.A(irq[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(irq[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(irq[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(mem_rdata[0]),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 input34 (.A(mem_rdata[10]),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(mem_rdata[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(mem_rdata[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(mem_rdata[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(mem_rdata[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(mem_rdata[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(mem_rdata[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_2 input41 (.A(mem_rdata[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(mem_rdata[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(mem_rdata[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(mem_rdata[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(mem_rdata[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(mem_rdata[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input47 (.A(mem_rdata[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input48 (.A(mem_rdata[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_2 input49 (.A(mem_rdata[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input50 (.A(mem_rdata[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input51 (.A(mem_rdata[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input52 (.A(mem_rdata[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input53 (.A(mem_rdata[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_2 input54 (.A(mem_rdata[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(mem_rdata[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(mem_rdata[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_2 input57 (.A(mem_rdata[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(mem_rdata[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(mem_rdata[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(mem_rdata[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(mem_rdata[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(mem_rdata[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(mem_rdata[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(mem_rdata[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 input65 (.A(mem_ready),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_8 input66 (.A(resetn),
    .X(net66));
 sky130_fd_sc_hd__buf_1 output67 (.A(net67),
    .X(cpi_rs1[0]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(cpi_rs1[10]));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(cpi_rs1[11]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(cpi_rs1[12]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .X(cpi_rs1[13]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .X(cpi_rs1[14]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(cpi_rs1[15]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(cpi_rs1[16]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .X(cpi_rs1[17]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(cpi_rs1[18]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(cpi_rs1[19]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(cpi_rs1[1]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(cpi_rs1[20]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net80),
    .X(cpi_rs1[21]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(cpi_rs1[22]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(cpi_rs1[23]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(cpi_rs1[24]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net84),
    .X(cpi_rs1[25]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(cpi_rs1[26]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(cpi_rs1[27]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net87),
    .X(cpi_rs1[28]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net88),
    .X(cpi_rs1[29]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net89),
    .X(cpi_rs1[2]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(cpi_rs1[30]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(cpi_rs1[31]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net92),
    .X(cpi_rs1[3]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(cpi_rs1[4]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(cpi_rs1[5]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net95),
    .X(cpi_rs1[6]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(cpi_rs1[7]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(cpi_rs1[8]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net98),
    .X(cpi_rs1[9]));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net99),
    .X(cpi_rs2[0]));
 sky130_fd_sc_hd__buf_1 output100 (.A(net100),
    .X(cpi_rs2[10]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net101),
    .X(cpi_rs2[11]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net102),
    .X(cpi_rs2[12]));
 sky130_fd_sc_hd__buf_1 output103 (.A(net103),
    .X(cpi_rs2[13]));
 sky130_fd_sc_hd__buf_1 output104 (.A(net104),
    .X(cpi_rs2[14]));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net105),
    .X(cpi_rs2[15]));
 sky130_fd_sc_hd__buf_1 output106 (.A(net106),
    .X(cpi_rs2[16]));
 sky130_fd_sc_hd__buf_1 output107 (.A(net107),
    .X(cpi_rs2[17]));
 sky130_fd_sc_hd__buf_1 output108 (.A(net108),
    .X(cpi_rs2[18]));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net109),
    .X(cpi_rs2[19]));
 sky130_fd_sc_hd__buf_1 output110 (.A(net110),
    .X(cpi_rs2[1]));
 sky130_fd_sc_hd__buf_1 output111 (.A(net111),
    .X(cpi_rs2[20]));
 sky130_fd_sc_hd__buf_1 output112 (.A(net112),
    .X(cpi_rs2[21]));
 sky130_fd_sc_hd__buf_1 output113 (.A(net113),
    .X(cpi_rs2[22]));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net114),
    .X(cpi_rs2[23]));
 sky130_fd_sc_hd__buf_1 output115 (.A(net115),
    .X(cpi_rs2[24]));
 sky130_fd_sc_hd__buf_1 output116 (.A(net116),
    .X(cpi_rs2[25]));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net117),
    .X(cpi_rs2[26]));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(net118),
    .X(cpi_rs2[27]));
 sky130_fd_sc_hd__buf_1 output119 (.A(net119),
    .X(cpi_rs2[28]));
 sky130_fd_sc_hd__buf_1 output120 (.A(net120),
    .X(cpi_rs2[29]));
 sky130_fd_sc_hd__buf_1 output121 (.A(net121),
    .X(cpi_rs2[2]));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(net122),
    .X(cpi_rs2[30]));
 sky130_fd_sc_hd__buf_1 output123 (.A(net123),
    .X(cpi_rs2[31]));
 sky130_fd_sc_hd__buf_1 output124 (.A(net124),
    .X(cpi_rs2[3]));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(net125),
    .X(cpi_rs2[4]));
 sky130_fd_sc_hd__buf_1 output126 (.A(net126),
    .X(cpi_rs2[5]));
 sky130_fd_sc_hd__buf_1 output127 (.A(net127),
    .X(cpi_rs2[6]));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(net128),
    .X(cpi_rs2[7]));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net129),
    .X(cpi_rs2[8]));
 sky130_fd_sc_hd__buf_1 output130 (.A(net130),
    .X(cpi_rs2[9]));
 sky130_fd_sc_hd__buf_1 output131 (.A(net131),
    .X(eoi[0]));
 sky130_fd_sc_hd__buf_1 output132 (.A(net132),
    .X(eoi[10]));
 sky130_fd_sc_hd__buf_1 output133 (.A(net133),
    .X(eoi[11]));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(net134),
    .X(eoi[12]));
 sky130_fd_sc_hd__buf_1 output135 (.A(net135),
    .X(eoi[13]));
 sky130_fd_sc_hd__buf_1 output136 (.A(net136),
    .X(eoi[14]));
 sky130_fd_sc_hd__buf_1 output137 (.A(net137),
    .X(eoi[15]));
 sky130_fd_sc_hd__clkbuf_1 output138 (.A(net138),
    .X(eoi[16]));
 sky130_fd_sc_hd__buf_1 output139 (.A(net139),
    .X(eoi[17]));
 sky130_fd_sc_hd__buf_1 output140 (.A(net140),
    .X(eoi[18]));
 sky130_fd_sc_hd__buf_1 output141 (.A(net141),
    .X(eoi[19]));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net142),
    .X(eoi[1]));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net143),
    .X(eoi[20]));
 sky130_fd_sc_hd__buf_1 output144 (.A(net144),
    .X(eoi[21]));
 sky130_fd_sc_hd__buf_1 output145 (.A(net145),
    .X(eoi[22]));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net146),
    .X(eoi[23]));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net147),
    .X(eoi[24]));
 sky130_fd_sc_hd__buf_1 output148 (.A(net148),
    .X(eoi[25]));
 sky130_fd_sc_hd__buf_1 output149 (.A(net149),
    .X(eoi[26]));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net150),
    .X(eoi[27]));
 sky130_fd_sc_hd__buf_1 output151 (.A(net151),
    .X(eoi[28]));
 sky130_fd_sc_hd__buf_1 output152 (.A(net152),
    .X(eoi[29]));
 sky130_fd_sc_hd__buf_1 output153 (.A(net153),
    .X(eoi[2]));
 sky130_fd_sc_hd__buf_1 output154 (.A(net154),
    .X(eoi[30]));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net155),
    .X(eoi[31]));
 sky130_fd_sc_hd__buf_1 output156 (.A(net156),
    .X(eoi[3]));
 sky130_fd_sc_hd__buf_1 output157 (.A(net157),
    .X(eoi[4]));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net158),
    .X(eoi[5]));
 sky130_fd_sc_hd__buf_1 output159 (.A(net159),
    .X(eoi[6]));
 sky130_fd_sc_hd__buf_1 output160 (.A(net160),
    .X(eoi[7]));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net161),
    .X(eoi[8]));
 sky130_fd_sc_hd__buf_1 output162 (.A(net162),
    .X(eoi[9]));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net163),
    .X(mem_addr[10]));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net164),
    .X(mem_addr[11]));
 sky130_fd_sc_hd__buf_1 output165 (.A(net165),
    .X(mem_addr[12]));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net166),
    .X(mem_addr[13]));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net167),
    .X(mem_addr[14]));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net168),
    .X(mem_addr[15]));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(net169),
    .X(mem_addr[16]));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net170),
    .X(mem_addr[17]));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net171),
    .X(mem_addr[18]));
 sky130_fd_sc_hd__buf_1 output172 (.A(net172),
    .X(mem_addr[19]));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net173),
    .X(mem_addr[20]));
 sky130_fd_sc_hd__buf_1 output174 (.A(net174),
    .X(mem_addr[21]));
 sky130_fd_sc_hd__clkbuf_1 output175 (.A(net175),
    .X(mem_addr[22]));
 sky130_fd_sc_hd__clkbuf_1 output176 (.A(net176),
    .X(mem_addr[23]));
 sky130_fd_sc_hd__clkbuf_1 output177 (.A(net177),
    .X(mem_addr[24]));
 sky130_fd_sc_hd__clkbuf_1 output178 (.A(net178),
    .X(mem_addr[25]));
 sky130_fd_sc_hd__buf_1 output179 (.A(net179),
    .X(mem_addr[26]));
 sky130_fd_sc_hd__clkbuf_1 output180 (.A(net180),
    .X(mem_addr[27]));
 sky130_fd_sc_hd__clkbuf_1 output181 (.A(net181),
    .X(mem_addr[28]));
 sky130_fd_sc_hd__buf_1 output182 (.A(net182),
    .X(mem_addr[29]));
 sky130_fd_sc_hd__clkbuf_1 output183 (.A(net183),
    .X(mem_addr[2]));
 sky130_fd_sc_hd__clkbuf_1 output184 (.A(net184),
    .X(mem_addr[30]));
 sky130_fd_sc_hd__buf_1 output185 (.A(net185),
    .X(mem_addr[31]));
 sky130_fd_sc_hd__clkbuf_1 output186 (.A(net186),
    .X(mem_addr[3]));
 sky130_fd_sc_hd__buf_1 output187 (.A(net187),
    .X(mem_addr[4]));
 sky130_fd_sc_hd__clkbuf_1 output188 (.A(net188),
    .X(mem_addr[5]));
 sky130_fd_sc_hd__buf_1 output189 (.A(net189),
    .X(mem_addr[6]));
 sky130_fd_sc_hd__clkbuf_1 output190 (.A(net190),
    .X(mem_addr[7]));
 sky130_fd_sc_hd__clkbuf_1 output191 (.A(net191),
    .X(mem_addr[8]));
 sky130_fd_sc_hd__buf_1 output192 (.A(net192),
    .X(mem_addr[9]));
 sky130_fd_sc_hd__clkbuf_1 output193 (.A(net193),
    .X(mem_instr));
 sky130_fd_sc_hd__buf_1 output194 (.A(net194),
    .X(mem_la_addr[10]));
 sky130_fd_sc_hd__clkbuf_1 output195 (.A(net195),
    .X(mem_la_addr[11]));
 sky130_fd_sc_hd__buf_1 output196 (.A(net196),
    .X(mem_la_addr[12]));
 sky130_fd_sc_hd__buf_1 output197 (.A(net197),
    .X(mem_la_addr[13]));
 sky130_fd_sc_hd__buf_1 output198 (.A(net198),
    .X(mem_la_addr[14]));
 sky130_fd_sc_hd__clkbuf_1 output199 (.A(net199),
    .X(mem_la_addr[15]));
 sky130_fd_sc_hd__buf_1 output200 (.A(net200),
    .X(mem_la_addr[16]));
 sky130_fd_sc_hd__buf_1 output201 (.A(net201),
    .X(mem_la_addr[17]));
 sky130_fd_sc_hd__buf_1 output202 (.A(net202),
    .X(mem_la_addr[18]));
 sky130_fd_sc_hd__clkbuf_1 output203 (.A(net203),
    .X(mem_la_addr[19]));
 sky130_fd_sc_hd__buf_1 output204 (.A(net204),
    .X(mem_la_addr[20]));
 sky130_fd_sc_hd__buf_1 output205 (.A(net205),
    .X(mem_la_addr[21]));
 sky130_fd_sc_hd__clkbuf_1 output206 (.A(net206),
    .X(mem_la_addr[22]));
 sky130_fd_sc_hd__clkbuf_1 output207 (.A(net207),
    .X(mem_la_addr[23]));
 sky130_fd_sc_hd__buf_1 output208 (.A(net208),
    .X(mem_la_addr[24]));
 sky130_fd_sc_hd__buf_1 output209 (.A(net209),
    .X(mem_la_addr[25]));
 sky130_fd_sc_hd__clkbuf_1 output210 (.A(net210),
    .X(mem_la_addr[26]));
 sky130_fd_sc_hd__buf_1 output211 (.A(net211),
    .X(mem_la_addr[27]));
 sky130_fd_sc_hd__buf_1 output212 (.A(net212),
    .X(mem_la_addr[28]));
 sky130_fd_sc_hd__buf_1 output213 (.A(net213),
    .X(mem_la_addr[29]));
 sky130_fd_sc_hd__buf_1 output214 (.A(net214),
    .X(mem_la_addr[2]));
 sky130_fd_sc_hd__clkbuf_1 output215 (.A(net215),
    .X(mem_la_addr[30]));
 sky130_fd_sc_hd__buf_1 output216 (.A(net216),
    .X(mem_la_addr[31]));
 sky130_fd_sc_hd__buf_1 output217 (.A(net217),
    .X(mem_la_addr[3]));
 sky130_fd_sc_hd__clkbuf_1 output218 (.A(net218),
    .X(mem_la_addr[4]));
 sky130_fd_sc_hd__buf_1 output219 (.A(net219),
    .X(mem_la_addr[5]));
 sky130_fd_sc_hd__buf_1 output220 (.A(net220),
    .X(mem_la_addr[6]));
 sky130_fd_sc_hd__clkbuf_1 output221 (.A(net221),
    .X(mem_la_addr[7]));
 sky130_fd_sc_hd__clkbuf_1 output222 (.A(net222),
    .X(mem_la_addr[8]));
 sky130_fd_sc_hd__buf_1 output223 (.A(net223),
    .X(mem_la_addr[9]));
 sky130_fd_sc_hd__clkbuf_1 output224 (.A(net224),
    .X(mem_la_read));
 sky130_fd_sc_hd__buf_1 output225 (.A(net225),
    .X(mem_la_wdata[0]));
 sky130_fd_sc_hd__clkbuf_1 output226 (.A(net226),
    .X(mem_la_wdata[10]));
 sky130_fd_sc_hd__buf_1 output227 (.A(net227),
    .X(mem_la_wdata[11]));
 sky130_fd_sc_hd__buf_1 output228 (.A(net228),
    .X(mem_la_wdata[12]));
 sky130_fd_sc_hd__clkbuf_1 output229 (.A(net229),
    .X(mem_la_wdata[13]));
 sky130_fd_sc_hd__clkbuf_1 output230 (.A(net230),
    .X(mem_la_wdata[14]));
 sky130_fd_sc_hd__buf_1 output231 (.A(net231),
    .X(mem_la_wdata[15]));
 sky130_fd_sc_hd__buf_1 output232 (.A(net232),
    .X(mem_la_wdata[16]));
 sky130_fd_sc_hd__clkbuf_1 output233 (.A(net233),
    .X(mem_la_wdata[17]));
 sky130_fd_sc_hd__buf_1 output234 (.A(net234),
    .X(mem_la_wdata[18]));
 sky130_fd_sc_hd__buf_1 output235 (.A(net235),
    .X(mem_la_wdata[19]));
 sky130_fd_sc_hd__buf_1 output236 (.A(net236),
    .X(mem_la_wdata[1]));
 sky130_fd_sc_hd__buf_1 output237 (.A(net237),
    .X(mem_la_wdata[20]));
 sky130_fd_sc_hd__clkbuf_1 output238 (.A(net238),
    .X(mem_la_wdata[21]));
 sky130_fd_sc_hd__buf_1 output239 (.A(net239),
    .X(mem_la_wdata[22]));
 sky130_fd_sc_hd__buf_1 output240 (.A(net240),
    .X(mem_la_wdata[23]));
 sky130_fd_sc_hd__clkbuf_1 output241 (.A(net241),
    .X(mem_la_wdata[24]));
 sky130_fd_sc_hd__clkbuf_1 output242 (.A(net242),
    .X(mem_la_wdata[25]));
 sky130_fd_sc_hd__buf_1 output243 (.A(net243),
    .X(mem_la_wdata[26]));
 sky130_fd_sc_hd__buf_1 output244 (.A(net244),
    .X(mem_la_wdata[27]));
 sky130_fd_sc_hd__clkbuf_1 output245 (.A(net245),
    .X(mem_la_wdata[28]));
 sky130_fd_sc_hd__buf_1 output246 (.A(net246),
    .X(mem_la_wdata[29]));
 sky130_fd_sc_hd__clkbuf_1 output247 (.A(net247),
    .X(mem_la_wdata[2]));
 sky130_fd_sc_hd__buf_1 output248 (.A(net248),
    .X(mem_la_wdata[30]));
 sky130_fd_sc_hd__buf_1 output249 (.A(net249),
    .X(mem_la_wdata[31]));
 sky130_fd_sc_hd__buf_1 output250 (.A(net250),
    .X(mem_la_wdata[3]));
 sky130_fd_sc_hd__buf_1 output251 (.A(net251),
    .X(mem_la_wdata[4]));
 sky130_fd_sc_hd__buf_1 output252 (.A(net252),
    .X(mem_la_wdata[5]));
 sky130_fd_sc_hd__clkbuf_1 output253 (.A(net253),
    .X(mem_la_wdata[6]));
 sky130_fd_sc_hd__buf_1 output254 (.A(net254),
    .X(mem_la_wdata[7]));
 sky130_fd_sc_hd__buf_1 output255 (.A(net255),
    .X(mem_la_wdata[8]));
 sky130_fd_sc_hd__clkbuf_1 output256 (.A(net256),
    .X(mem_la_wdata[9]));
 sky130_fd_sc_hd__clkbuf_1 output257 (.A(net257),
    .X(mem_la_write));
 sky130_fd_sc_hd__buf_1 output258 (.A(net258),
    .X(mem_la_wstrb[0]));
 sky130_fd_sc_hd__buf_1 output259 (.A(net259),
    .X(mem_la_wstrb[1]));
 sky130_fd_sc_hd__clkbuf_1 output260 (.A(net260),
    .X(mem_la_wstrb[2]));
 sky130_fd_sc_hd__buf_1 output261 (.A(net261),
    .X(mem_la_wstrb[3]));
 sky130_fd_sc_hd__buf_1 output262 (.A(net262),
    .X(mem_valid));
 sky130_fd_sc_hd__clkbuf_1 output263 (.A(net263),
    .X(mem_wdata[0]));
 sky130_fd_sc_hd__clkbuf_1 output264 (.A(net264),
    .X(mem_wdata[10]));
 sky130_fd_sc_hd__buf_1 output265 (.A(net265),
    .X(mem_wdata[11]));
 sky130_fd_sc_hd__clkbuf_1 output266 (.A(net266),
    .X(mem_wdata[12]));
 sky130_fd_sc_hd__clkbuf_1 output267 (.A(net267),
    .X(mem_wdata[13]));
 sky130_fd_sc_hd__clkbuf_1 output268 (.A(net268),
    .X(mem_wdata[14]));
 sky130_fd_sc_hd__clkbuf_1 output269 (.A(net269),
    .X(mem_wdata[15]));
 sky130_fd_sc_hd__buf_1 output270 (.A(net270),
    .X(mem_wdata[16]));
 sky130_fd_sc_hd__clkbuf_1 output271 (.A(net271),
    .X(mem_wdata[17]));
 sky130_fd_sc_hd__buf_1 output272 (.A(net272),
    .X(mem_wdata[18]));
 sky130_fd_sc_hd__clkbuf_1 output273 (.A(net273),
    .X(mem_wdata[19]));
 sky130_fd_sc_hd__clkbuf_1 output274 (.A(net274),
    .X(mem_wdata[1]));
 sky130_fd_sc_hd__clkbuf_1 output275 (.A(net275),
    .X(mem_wdata[20]));
 sky130_fd_sc_hd__clkbuf_1 output276 (.A(net276),
    .X(mem_wdata[21]));
 sky130_fd_sc_hd__clkbuf_1 output277 (.A(net277),
    .X(mem_wdata[22]));
 sky130_fd_sc_hd__clkbuf_1 output278 (.A(net278),
    .X(mem_wdata[23]));
 sky130_fd_sc_hd__clkbuf_1 output279 (.A(net279),
    .X(mem_wdata[24]));
 sky130_fd_sc_hd__clkbuf_1 output280 (.A(net280),
    .X(mem_wdata[25]));
 sky130_fd_sc_hd__clkbuf_1 output281 (.A(net281),
    .X(mem_wdata[26]));
 sky130_fd_sc_hd__clkbuf_1 output282 (.A(net282),
    .X(mem_wdata[27]));
 sky130_fd_sc_hd__clkbuf_1 output283 (.A(net283),
    .X(mem_wdata[28]));
 sky130_fd_sc_hd__clkbuf_1 output284 (.A(net284),
    .X(mem_wdata[29]));
 sky130_fd_sc_hd__clkbuf_1 output285 (.A(net285),
    .X(mem_wdata[2]));
 sky130_fd_sc_hd__clkbuf_1 output286 (.A(net286),
    .X(mem_wdata[30]));
 sky130_fd_sc_hd__clkbuf_1 output287 (.A(net287),
    .X(mem_wdata[31]));
 sky130_fd_sc_hd__clkbuf_1 output288 (.A(net288),
    .X(mem_wdata[3]));
 sky130_fd_sc_hd__buf_1 output289 (.A(net289),
    .X(mem_wdata[4]));
 sky130_fd_sc_hd__clkbuf_1 output290 (.A(net290),
    .X(mem_wdata[5]));
 sky130_fd_sc_hd__clkbuf_1 output291 (.A(net291),
    .X(mem_wdata[6]));
 sky130_fd_sc_hd__clkbuf_1 output292 (.A(net292),
    .X(mem_wdata[7]));
 sky130_fd_sc_hd__clkbuf_1 output293 (.A(net293),
    .X(mem_wdata[8]));
 sky130_fd_sc_hd__buf_1 output294 (.A(net294),
    .X(mem_wdata[9]));
 sky130_fd_sc_hd__clkbuf_1 output295 (.A(net295),
    .X(mem_wstrb[0]));
 sky130_fd_sc_hd__buf_1 output296 (.A(net296),
    .X(mem_wstrb[1]));
 sky130_fd_sc_hd__buf_1 output297 (.A(net297),
    .X(mem_wstrb[2]));
 sky130_fd_sc_hd__clkbuf_1 output298 (.A(net298),
    .X(mem_wstrb[3]));
 sky130_fd_sc_hd__buf_1 output299 (.A(net299),
    .X(trap));
 sky130_fd_sc_hd__buf_4 max_cap300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__buf_4 max_cap301 (.A(_04099_),
    .X(net301));
 sky130_fd_sc_hd__conb_1 alphacore_302 (.LO(net302));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_3_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_4_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_5_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_6_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_7_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_8_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_9_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_10_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_11_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_12_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_13_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_14_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_15_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_16_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_17_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_18_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_19_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_20_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_21_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_22_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_23_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_24_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_25_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_26_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_27_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_28_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_29_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_30_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_31_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_32_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_33_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_34_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_35_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_36_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_37_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_38_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_39_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_40_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_41_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_42_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_43_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_44_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_45_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_46_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_47_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_48_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_49_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_50_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_51_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_52_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_53_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_54_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_55_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_56_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_57_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_58_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_59_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_60_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_61_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_62_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_63_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_64_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_65_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_66_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_67_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_68_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_69_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_70_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_71_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_72_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_73_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_74_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_75_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_76_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_77_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_78_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_79_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_80_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_81_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_82_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_83_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_84_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_85_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_86_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_87_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_88_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_89_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_90_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_91_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_92_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_93_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_94_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_95_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_96_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_97_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_98_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_99_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_100_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_101_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_102_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_103_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_104_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_105_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_106_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_107_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_108_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_109_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_110_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_111_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_112_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_113_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_114_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_115_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_116_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_117_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_118_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_119_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_120_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_121_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_122_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_123_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_124_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_125_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_126_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_127_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_128_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_129_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_130_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_131_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_132_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_133_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_134_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_135_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_136_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_137_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_138_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_139_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_140_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_141_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_142_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_143_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_144_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_145_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_146_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_147_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_148_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_149_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_150_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_151_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_152_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_153_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_154_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_155_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_156_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_157_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_158_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_159_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_160_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_161_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_162_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_163_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_164_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_165_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_166_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_167_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_168_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_169_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_170_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_171_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_172_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_173_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_174_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_175_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_176_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_177_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_178_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_179_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_180_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_181_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_182_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_183_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_184_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_185_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_186_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_187_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_188_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_189_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_190_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_leaf_191_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__A (.DIODE(_00064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08896__A (.DIODE(_00064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08893__A (.DIODE(_00064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__A (.DIODE(_00064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__A (.DIODE(_00065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08894__A (.DIODE(_00065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__A (.DIODE(_00065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__A (.DIODE(_00065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15415__B1 (.DIODE(_00067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15192__B1 (.DIODE(_00067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15090__C1 (.DIODE(_00067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15082__C1 (.DIODE(_00067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__B1 (.DIODE(_00067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__A (.DIODE(_00067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08889__A (.DIODE(_00067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15627__A1 (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15616__B1 (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15535__B1 (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15395__B1 (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15086__B1 (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__A (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__A (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08874__A (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__S (.DIODE(_00071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__S (.DIODE(_00071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__A (.DIODE(_00071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__A (.DIODE(_00071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__S (.DIODE(_00071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09392__A (.DIODE(_00071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09328__A (.DIODE(_00071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10396__B1 (.DIODE(_00073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__B1 (.DIODE(_00073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__A (.DIODE(_00073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__B1 (.DIODE(_00073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__C1 (.DIODE(_00073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A (.DIODE(_00073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__A (.DIODE(_00073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16947__D (.DIODE(_00075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17696__D (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__C (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18049__D (.DIODE(_01154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18081__D (.DIODE(_01186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18224__D (.DIODE(_01295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15029__B1 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15023__B1 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15021__B1 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14995__B1 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14884__B1 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14869__B1 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14860__B1 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14851__B1 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14842__B1 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14745__A (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14833__B1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14824__B1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14815__B1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14806__B1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14796__B1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14786__B1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14777__B1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__B1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14758__B1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14748__B1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14858__B1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14849__B1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14840__B1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14831__B1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14822__B1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14813__B1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14804__B1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14775__B1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14765__B1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14756__B1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14882__B (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14873__B (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14864__B (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14855__B (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14846__B (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14837__B (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14828__B (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14819__B (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14810__B (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14801__B (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14942__A (.DIODE(_01823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14921__A (.DIODE(_01823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14900__A (.DIODE(_01823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15043__B (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15041__B (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15039__B (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15037__B (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15031__A2 (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15029__A2 (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15023__A2 (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15021__A2 (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14995__A2 (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14972__A (.DIODE(_01863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15044__A2 (.DIODE(_01865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15042__A2 (.DIODE(_01865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15040__A2 (.DIODE(_01865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15038__A2 (.DIODE(_01865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15036__A2 (.DIODE(_01865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15034__A2 (.DIODE(_01865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15028__A2 (.DIODE(_01865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14978__B (.DIODE(_01865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14976__B (.DIODE(_01865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14974__B (.DIODE(_01865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15678__A1 (.DIODE(_01872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14986__A (.DIODE(_01872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15700__A (.DIODE(_01881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15001__A (.DIODE(_01881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15035__B (.DIODE(_01885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15033__B (.DIODE(_01885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15027__B (.DIODE(_01885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15025__B (.DIODE(_01885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15019__B (.DIODE(_01885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15016__B (.DIODE(_01885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15014__B (.DIODE(_01885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15012__B (.DIODE(_01885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15010__B (.DIODE(_01885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15008__B (.DIODE(_01885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15582__A2 (.DIODE(_01905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15566__A2 (.DIODE(_01905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15531__A2 (.DIODE(_01905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15515__A2 (.DIODE(_01905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15477__A2 (.DIODE(_01905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15428__S (.DIODE(_01905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15409__S (.DIODE(_01905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15230__A (.DIODE(_01905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15207__S (.DIODE(_01905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15046__A (.DIODE(_01905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15612__A2 (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15597__A2 (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15391__A2 (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15229__A2 (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15187__A2 (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15156__A2 (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15112__A2 (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15105__A2 (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15099__A2 (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15076__A2 (.DIODE(_01906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15600__S (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15585__S (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15562__S (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15527__S (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15457__S (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15437__S (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15377__S (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15127__A (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15063__A1 (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15053__A1 (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15607__S0 (.DIODE(_01908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15599__S0 (.DIODE(_01908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15598__S0 (.DIODE(_01908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15592__S0 (.DIODE(_01908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15584__S0 (.DIODE(_01908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15583__S0 (.DIODE(_01908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15386__S0 (.DIODE(_01908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15376__S0 (.DIODE(_01908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15375__S0 (.DIODE(_01908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15050__S0 (.DIODE(_01908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15607__S1 (.DIODE(_01909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15599__S1 (.DIODE(_01909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15598__S1 (.DIODE(_01909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15592__S1 (.DIODE(_01909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15584__S1 (.DIODE(_01909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15583__S1 (.DIODE(_01909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15386__S1 (.DIODE(_01909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15376__S1 (.DIODE(_01909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15375__S1 (.DIODE(_01909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15050__S1 (.DIODE(_01909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15573__S0 (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15572__S0 (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15436__S0 (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15435__S0 (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15234__A (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15124__A (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15121__A (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15118__A (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15115__A (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15060__S0 (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15573__S1 (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15572__S1 (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15436__S1 (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15435__S1 (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15235__A (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15125__A (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15122__A (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15119__A (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15116__A (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15060__S1 (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16743__B1 (.DIODE(_01929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15070__B (.DIODE(_01929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15629__B1 (.DIODE(_01932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15372__A (.DIODE(_01932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15110__B2 (.DIODE(_01932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15103__B2 (.DIODE(_01932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15073__A (.DIODE(_01932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15611__A2 (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15548__B1 (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15494__B1 (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15427__B1 (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15408__B1 (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15206__B1 (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15154__A (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15107__B2 (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15098__B2 (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15075__B2 (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15611__C1 (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15596__C1 (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15352__A (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15110__C1 (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15107__C1 (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15106__A (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15103__C1 (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15098__C1 (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15075__C1 (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15414__S0 (.DIODE(_01936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15394__S0 (.DIODE(_01936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15217__A (.DIODE(_01936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15191__S0 (.DIODE(_01936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15168__A (.DIODE(_01936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15159__A (.DIODE(_01936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15135__A (.DIODE(_01936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15130__A (.DIODE(_01936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15087__S0 (.DIODE(_01936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15079__S0 (.DIODE(_01936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15615__S1 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15613__S1 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15534__S1 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15532__S1 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15480__S1 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15478__S1 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15394__S1 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15392__S1 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15223__A (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15079__S1 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15096__B (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16745__B (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15097__B (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15629__A1 (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15611__B1 (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15596__B1 (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15548__A1 (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15494__A1 (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15427__A1 (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15408__A1 (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15206__A1 (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15173__A (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15102__A (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15459__C1 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15443__C1 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15351__C1 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15335__C1 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15300__C1 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15284__C1 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15247__C1 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15227__C1 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15153__C1 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15104__A2 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15105__B1 (.DIODE(_01962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15336__B1 (.DIODE(_01963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15320__B1 (.DIODE(_01963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15301__B1 (.DIODE(_01963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15285__B1 (.DIODE(_01963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15269__B1 (.DIODE(_01963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15248__B1 (.DIODE(_01963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15228__B1 (.DIODE(_01963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15186__B1 (.DIODE(_01963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15155__B1 (.DIODE(_01963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15109__A2 (.DIODE(_01963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15109__B1 (.DIODE(_01965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15610__S0 (.DIODE(_01968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15595__S0 (.DIODE(_01968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15576__B1 (.DIODE(_01968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15539__C1 (.DIODE(_01968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15485__C1 (.DIODE(_01968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15439__B1 (.DIODE(_01968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15399__C1 (.DIODE(_01968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15389__S0 (.DIODE(_01968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15366__B1 (.DIODE(_01968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15114__A (.DIODE(_01968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15564__A1 (.DIODE(_01969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15529__A1 (.DIODE(_01969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15512__C1 (.DIODE(_01969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15475__A1 (.DIODE(_01969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15335__A1 (.DIODE(_01969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15318__C1 (.DIODE(_01969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15267__C1 (.DIODE(_01969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15227__A1 (.DIODE(_01969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15184__C1 (.DIODE(_01969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15153__A1 (.DIODE(_01969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15497__S0 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15355__S0 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15303__S0 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15287__S0 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15271__S0 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15250__S0 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15231__S0 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15209__S0 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15157__S0 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15117__S0 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15497__S1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15355__S1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15303__S1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15287__S1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15271__S1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15250__S1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15231__S1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15209__S1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15157__S1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15117__S1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15569__S0 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15553__S0 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15518__S0 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15464__S0 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15323__S0 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15288__S0 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15272__S0 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15232__S0 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15210__S0 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15120__S0 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15569__S1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15553__S1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15518__S1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15464__S1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15323__S1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15288__S1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15272__S1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15232__S1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15210__S1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15120__S1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15570__S0 (.DIODE(_01976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15448__S0 (.DIODE(_01976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15432__S0 (.DIODE(_01976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15340__S0 (.DIODE(_01976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15324__S0 (.DIODE(_01976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15289__S0 (.DIODE(_01976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15273__S0 (.DIODE(_01976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15233__S0 (.DIODE(_01976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15211__S0 (.DIODE(_01976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15123__S0 (.DIODE(_01976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15570__S1 (.DIODE(_01977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15448__S1 (.DIODE(_01977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15432__S1 (.DIODE(_01977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15340__S1 (.DIODE(_01977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15324__S1 (.DIODE(_01977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15289__S1 (.DIODE(_01977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15273__S1 (.DIODE(_01977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15233__S1 (.DIODE(_01977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15211__S1 (.DIODE(_01977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15123__S1 (.DIODE(_01977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15567__S0 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15551__S0 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15516__S0 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15462__S0 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15446__S0 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15430__S0 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15338__S0 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15322__S0 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15212__S0 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15126__S0 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15567__S1 (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15551__S1 (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15516__S1 (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15462__S1 (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15446__S1 (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15430__S1 (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15338__S1 (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15322__S1 (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15212__S1 (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15126__S1 (.DIODE(_01980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15500__A1 (.DIODE(_01982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15358__A1 (.DIODE(_01982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15326__S0 (.DIODE(_01982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15306__A1 (.DIODE(_01982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15291__S0 (.DIODE(_01982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15275__S0 (.DIODE(_01982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15253__A1 (.DIODE(_01982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15238__S0 (.DIODE(_01982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15213__S0 (.DIODE(_01982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15128__S0 (.DIODE(_01982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15557__A (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15506__A (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15503__S (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15468__A (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15361__S (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15309__S (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15293__A (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15240__A (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15171__S (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15133__A (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15510__S0 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15368__S0 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15316__S0 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15292__S0 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15276__S0 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15265__S0 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15239__S0 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15215__S0 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15181__S0 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15132__S0 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15510__S1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15368__S1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15316__S1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15292__S1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15276__S1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15265__S1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15239__S1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15215__S1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15181__S1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15132__S1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15508__A1 (.DIODE(_01989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15499__A (.DIODE(_01989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15357__A (.DIODE(_01989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15314__A1 (.DIODE(_01989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15305__A (.DIODE(_01989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15252__A (.DIODE(_01989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15242__A1 (.DIODE(_01989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15179__A1 (.DIODE(_01989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15165__A1 (.DIODE(_01989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15139__A1 (.DIODE(_01989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15505__S0 (.DIODE(_01990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15501__S0 (.DIODE(_01990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15363__S0 (.DIODE(_01990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15359__S0 (.DIODE(_01990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15311__S0 (.DIODE(_01990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15307__S0 (.DIODE(_01990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15258__S0 (.DIODE(_01990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15254__S0 (.DIODE(_01990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15167__S0 (.DIODE(_01990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15138__S0 (.DIODE(_01990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15621__S1 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15540__S1 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15487__S1 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15486__S1 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15420__S1 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15419__S1 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15401__S1 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15218__A (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15199__S1 (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15137__A (.DIODE(_01991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15505__S1 (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15501__S1 (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15363__S1 (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15359__S1 (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15311__S1 (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15307__S1 (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15258__S1 (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15254__S1 (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15167__S1 (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15138__S1 (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15615__S0 (.DIODE(_01995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15613__S0 (.DIODE(_01995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15534__S0 (.DIODE(_01995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15532__S0 (.DIODE(_01995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15480__S0 (.DIODE(_01995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15478__S0 (.DIODE(_01995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15392__S0 (.DIODE(_01995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15222__A (.DIODE(_01995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15144__A (.DIODE(_01995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15141__A (.DIODE(_01995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15577__S0 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15556__S0 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15521__S0 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15467__S0 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15451__S0 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15440__S0 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15343__S0 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15327__S0 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15221__S0 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15143__S0 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15577__S1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15556__S1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15521__S1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15467__S1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15451__S1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15440__S1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15343__S1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15327__S1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15221__S1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15143__S1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15560__S0 (.DIODE(_01999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15525__S0 (.DIODE(_01999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15471__S0 (.DIODE(_01999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15455__S0 (.DIODE(_01999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15347__S0 (.DIODE(_01999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15331__S0 (.DIODE(_01999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15296__S0 (.DIODE(_01999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15280__S0 (.DIODE(_01999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15243__S0 (.DIODE(_01999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15146__S0 (.DIODE(_01999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15560__S1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15525__S1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15471__S1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15455__S1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15347__S1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15331__S1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15296__S1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15280__S1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15243__S1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15146__S1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15511__S (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15369__S (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15349__S (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15333__S (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15317__S (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15298__S (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15282__S (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15266__S (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15182__S (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15148__S (.DIODE(_02002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15579__C1 (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15563__B2 (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15555__S1 (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15474__B2 (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15466__S1 (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15458__C1 (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15407__A1 (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15318__B2 (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15213__S1 (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15152__B2 (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15571__S1 (.DIODE(_02005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15454__B1 (.DIODE(_02005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15426__A1 (.DIODE(_02005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15418__A1 (.DIODE(_02005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15346__B1 (.DIODE(_02005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15279__B1 (.DIODE(_02005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15237__A (.DIODE(_02005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15205__A1 (.DIODE(_02005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15197__A1 (.DIODE(_02005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15151__A (.DIODE(_02005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15528__C1 (.DIODE(_02006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15504__B1 (.DIODE(_02006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15474__C1 (.DIODE(_02006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15358__C1 (.DIODE(_02006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15334__C1 (.DIODE(_02006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15310__B1 (.DIODE(_02006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15257__B1 (.DIODE(_02006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15226__C1 (.DIODE(_02006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15172__B1 (.DIODE(_02006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15152__C1 (.DIODE(_02006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15353__A2 (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15336__A2 (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15320__A2 (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15301__A2 (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15285__A2 (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15269__A2 (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15248__A2 (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15228__A2 (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15186__A2 (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15155__A2 (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15524__A1 (.DIODE(_02012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15454__A1 (.DIODE(_02012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15366__A1 (.DIODE(_02012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15346__A1 (.DIODE(_02012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15330__A1 (.DIODE(_02012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15312__A (.DIODE(_02012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15279__A1 (.DIODE(_02012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15220__A1 (.DIODE(_02012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15175__A (.DIODE(_02012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15162__A (.DIODE(_02012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15507__S0 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15498__S0 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15365__S0 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15356__S0 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15313__S0 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15304__S0 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15262__S0 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15251__S0 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15174__S0 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15161__S0 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15507__S1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15498__S1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15365__S1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15356__S1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15313__S1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15304__S1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15262__S1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15251__S1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15174__S1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15161__S1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15628__A1 (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15539__B2 (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15524__B1 (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15508__B1 (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15399__B2 (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15330__B1 (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15263__B1 (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15220__B1 (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15179__B1 (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15164__A (.DIODE(_02017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15500__C1 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15442__C1 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15362__B1 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15350__C1 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15306__C1 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15299__C1 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15283__C1 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15253__C1 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15246__C1 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15165__C1 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15580__A1 (.DIODE(_02020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15459__A1 (.DIODE(_02020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15443__A1 (.DIODE(_02020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15370__C1 (.DIODE(_02020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15351__A1 (.DIODE(_02020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15300__A1 (.DIODE(_02020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15284__A1 (.DIODE(_02020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15257__A1 (.DIODE(_02020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15247__A1 (.DIODE(_02020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15172__A1 (.DIODE(_02020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15509__S0 (.DIODE(_02022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15502__S0 (.DIODE(_02022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15367__S0 (.DIODE(_02022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15360__S0 (.DIODE(_02022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15315__S0 (.DIODE(_02022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15308__S0 (.DIODE(_02022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15264__S0 (.DIODE(_02022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15255__S0 (.DIODE(_02022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15180__S0 (.DIODE(_02022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15170__S0 (.DIODE(_02022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15509__S1 (.DIODE(_02023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15502__S1 (.DIODE(_02023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15367__S1 (.DIODE(_02023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15360__S1 (.DIODE(_02023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15315__S1 (.DIODE(_02023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15308__S1 (.DIODE(_02023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15264__S1 (.DIODE(_02023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15255__S1 (.DIODE(_02023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15180__S1 (.DIODE(_02023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15170__S1 (.DIODE(_02023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15580__C1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15564__C1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15529__C1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15513__B1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15475__C1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15390__B1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15371__B1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15319__B1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15268__B1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15185__B1 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15575__S0 (.DIODE(_02030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15568__S0 (.DIODE(_02030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15552__S0 (.DIODE(_02030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15517__S0 (.DIODE(_02030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15463__S0 (.DIODE(_02030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15447__S0 (.DIODE(_02030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15438__S0 (.DIODE(_02030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15431__S0 (.DIODE(_02030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15339__S0 (.DIODE(_02030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15178__S0 (.DIODE(_02030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15575__S1 (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15568__S1 (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15552__S1 (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15517__S1 (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15463__S1 (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15447__S1 (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15438__S1 (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15431__S1 (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15339__S1 (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15178__S1 (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15595__S1 (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15528__B2 (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15512__B2 (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15504__A1 (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15389__S1 (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15334__B2 (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15310__A1 (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15267__B2 (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15226__B2 (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15184__B2 (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15187__B1 (.DIODE(_02039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15618__S0 (.DIODE(_02046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15617__S0 (.DIODE(_02046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15537__S0 (.DIODE(_02046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15536__S0 (.DIODE(_02046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15483__S0 (.DIODE(_02046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15482__S0 (.DIODE(_02046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15416__S0 (.DIODE(_02046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15397__S0 (.DIODE(_02046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15396__S0 (.DIODE(_02046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15195__S0 (.DIODE(_02046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15618__S1 (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15617__S1 (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15537__S1 (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15536__S1 (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15483__S1 (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15482__S1 (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15416__S1 (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15397__S1 (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15396__S1 (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15195__S1 (.DIODE(_02047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15206__A2 (.DIODE(_02050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15206__A3 (.DIODE(_02058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15559__A1 (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15470__A1 (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15452__A (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15364__A (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15344__A (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15328__A (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15295__A1 (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15277__A (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15259__A (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15216__A (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15558__S0 (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15523__S0 (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15469__S0 (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15453__S0 (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15345__S0 (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15329__S0 (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15294__S0 (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15278__S0 (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15241__S0 (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15219__S0 (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15558__S1 (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15523__S1 (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15469__S1 (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15453__S1 (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15345__S1 (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15329__S1 (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15294__S1 (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15278__S1 (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15241__S1 (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15219__S1 (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15561__S0 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15526__S0 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15472__S0 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15456__S0 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15348__S0 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15332__S0 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15297__S0 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15281__S0 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15244__S0 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15224__S0 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15561__S1 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15526__S1 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15472__S1 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15456__S1 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15348__S1 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15332__S1 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15297__S1 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15281__S1 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15244__S1 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15224__S1 (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15229__B1 (.DIODE(_02079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15554__S0 (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15519__S0 (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15465__S0 (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15449__S0 (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15433__S0 (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15341__S0 (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15325__S0 (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15290__S0 (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15274__S0 (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15236__S0 (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15554__S1 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15519__S1 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15465__S1 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15449__S1 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15433__S1 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15341__S1 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15325__S1 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15290__S1 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15274__S1 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15236__S1 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15579__A1 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15563__C1 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15442__A1 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15434__S1 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15370__B2 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15342__S1 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15299__B2 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15275__S1 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15246__B2 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15238__S1 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15249__B1 (.DIODE(_02098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15609__S (.DIODE(_02110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15606__S (.DIODE(_02110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15603__S (.DIODE(_02110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15594__S (.DIODE(_02110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15591__S (.DIODE(_02110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15588__S (.DIODE(_02110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15388__S (.DIODE(_02110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15385__S (.DIODE(_02110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15382__S (.DIODE(_02110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15261__A (.DIODE(_02110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15576__A1 (.DIODE(_02111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15571__S0 (.DIODE(_02111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15555__S0 (.DIODE(_02111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15520__S0 (.DIODE(_02111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15466__S0 (.DIODE(_02111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15450__S0 (.DIODE(_02111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15439__A1 (.DIODE(_02111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15434__S0 (.DIODE(_02111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15342__S0 (.DIODE(_02111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15263__A1 (.DIODE(_02111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15270__B1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15286__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15302__B1 (.DIODE(_02148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15321__B1 (.DIODE(_02166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15337__B1 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15354__B1 (.DIODE(_02196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15581__B1 (.DIODE(_02197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15565__B1 (.DIODE(_02197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15530__B1 (.DIODE(_02197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15514__B1 (.DIODE(_02197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15476__B1 (.DIODE(_02197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15460__B1 (.DIODE(_02197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15444__B1 (.DIODE(_02197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15390__C1 (.DIODE(_02197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15373__B1 (.DIODE(_02197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15353__B1 (.DIODE(_02197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15374__B1 (.DIODE(_02215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15596__A2 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15581__A2 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15565__A2 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15530__A2 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15514__A2 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15476__A2 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15460__A2 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15444__A2 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15390__A2 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15373__A2 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15608__S0 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15605__S0 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15604__S0 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15593__S0 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15590__S0 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15589__S0 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15387__S0 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15384__S0 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15383__S0 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15380__S0 (.DIODE(_02221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15608__S1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15605__S1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15604__S1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15593__S1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15590__S1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15589__S1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15387__S1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15384__S1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15383__S1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15380__S1 (.DIODE(_02222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15390__B2 (.DIODE(_02232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15391__B1 (.DIODE(_02233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15408__A2 (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15408__A3 (.DIODE(_02249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15409__A1 (.DIODE(_02250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15427__A2 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15427__A3 (.DIODE(_02267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15428__A1 (.DIODE(_02268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15445__B1 (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15461__B1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15477__B1 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15495__A1 (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15515__B1 (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15531__B1 (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15549__A1 (.DIODE(_02382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15566__B1 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15582__B1 (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15596__B2 (.DIODE(_02426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15597__B1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15611__B2 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15612__B1 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15629__A2 (.DIODE(_02449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15629__A3 (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15630__A1 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15774__C1 (.DIODE(_02476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15754__A (.DIODE(_02476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15747__A (.DIODE(_02476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15735__A (.DIODE(_02476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15728__A (.DIODE(_02476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15716__A (.DIODE(_02476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15705__A2 (.DIODE(_02476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15696__B1 (.DIODE(_02476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15688__B1 (.DIODE(_02476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15653__A (.DIODE(_02476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15763__A1 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15725__A1 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15713__A2 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15701__A1 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15686__A1 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15681__A1 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15675__A2 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15672__A2 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15663__A2 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15658__A1 (.DIODE(_02477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15762__B (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15758__B (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15757__B1 (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15724__B (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15720__B (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15700__B (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15685__B (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15680__B (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15678__A2 (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15656__B (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15770__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15712__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15694__A1 (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15671__A1 (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15664__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15662__B1 (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15778__A2 (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15777__B1 (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15775__A2 (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15772__A2 (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15768__A2 (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15755__A2 (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15698__A2 (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15691__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15690__A2 (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15668__A2 (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15767__C1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15749__B1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15741__B1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15738__B1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15730__B1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15718__B1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15707__B1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15677__B1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15674__B1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15667__B1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15773__B (.DIODE(_02560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15767__A2 (.DIODE(_02560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15765__C (.DIODE(_02560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16067__A (.DIODE(_02610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16064__B (.DIODE(_02610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16031__C (.DIODE(_02610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15971__B (.DIODE(_02610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15915__A (.DIODE(_02610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15897__C (.DIODE(_02610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15862__C (.DIODE(_02610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15856__B (.DIODE(_02610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15851__A (.DIODE(_02610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16063__A2 (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16022__A (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16010__A (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15911__A (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15909__B (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15895__A2 (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15890__B (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15885__A (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15883__A (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15858__A2 (.DIODE(_02611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16048__B2 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15900__C (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15896__A (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15887__A (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15872__A (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15870__A_N (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15867__C (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15865__A (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15860__B_N (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15854__A (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16050__B2 (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15900__B (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15896__C_N (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15887__C_N (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15872__B (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15870__B (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15867__A_N (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15865__B (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15860__A (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15854__B (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15951__A2 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15929__A2 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15928__A2 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15925__A2 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15924__A2 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15923__A2 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15922__A2 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15917__A2 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15904__A2 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15858__B1 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15922__B1 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15909__C (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15885__B (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15864__B1 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15925__B1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15902__B1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15891__B1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15866__B2 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15930__B (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15927__A1 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15926__A1 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15913__A2 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15892__B1 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15869__B2 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16088__B1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16042__C1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16040__C1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16038__C1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16036__C1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16034__C1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16032__A2 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16012__C1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15888__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15882__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15979__A2 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15910__A2 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15905__A2 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15894__A2 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15893__A2 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15892__A2 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15891__A2 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15889__A2 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15886__A2 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15884__A2 (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16087__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16070__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16069__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15973__B1 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15947__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15946__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15943__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15940__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15931__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15913__B1 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15946__B1 (.DIODE(_02659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15940__B1 (.DIODE(_02659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15943__B1 (.DIODE(_02665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15940__B2 (.DIODE(_02665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15947__B1 (.DIODE(_02667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15943__B2 (.DIODE(_02667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15947__B2 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15946__B2 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15979__B1 (.DIODE(_02695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16089__A2 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16043__A2 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16041__A2 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16039__A2 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16037__A2 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16035__A2 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16033__A2 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16021__A2 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16018__A2 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16013__A2 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16185__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16183__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16181__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16179__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16158__A (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16137__A (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16111__A (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16135__S (.DIODE(_02771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16133__S (.DIODE(_02771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16131__S (.DIODE(_02771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16129__S (.DIODE(_02771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16127__S (.DIODE(_02771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16125__S (.DIODE(_02771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16123__S (.DIODE(_02771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16121__S (.DIODE(_02771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16120__B2 (.DIODE(_02771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16112__B1_N (.DIODE(_02771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16286__S (.DIODE(_02859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16284__S (.DIODE(_02859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16282__S (.DIODE(_02859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16280__S (.DIODE(_02859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16278__S (.DIODE(_02859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16276__S (.DIODE(_02859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16274__S (.DIODE(_02859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16272__S (.DIODE(_02859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16270__S (.DIODE(_02859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16268__S (.DIODE(_02859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16307__S (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16305__S (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16303__S (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16301__S (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16299__S (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16297__S (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16295__S (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16293__S (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16291__S (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16289__S (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16328__S (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16326__S (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16324__S (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16322__S (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16320__S (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16318__S (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16316__S (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16314__S (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16312__S (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16310__S (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16401__S (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16399__S (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16378__A (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16357__A (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16336__A (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16355__S (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16353__S (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16351__S (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16349__S (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16347__S (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16345__S (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16343__S (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16341__S (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16339__S (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16337__S (.DIODE(_02896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16376__S (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16374__S (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16372__S (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16370__S (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16368__S (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16366__S (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16364__S (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16362__S (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16360__S (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16358__S (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16397__S (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16395__S (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16393__S (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16391__S (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16389__S (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16387__S (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16385__S (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16383__S (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16381__S (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16379__S (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16469__S (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16467__S (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16446__A (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16425__A (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16404__A (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16423__S (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16421__S (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16419__S (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16417__S (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16415__S (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16413__S (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16411__S (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16409__S (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16407__S (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16405__S (.DIODE(_02932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16444__S (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16442__S (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16440__S (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16438__S (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16436__S (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16434__S (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16432__S (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16430__S (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16428__S (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16426__S (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16465__S (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16463__S (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16461__S (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16459__S (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16457__S (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16455__S (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16453__S (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16451__S (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16449__S (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16447__S (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16537__S (.DIODE(_02967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16535__S (.DIODE(_02967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16514__A (.DIODE(_02967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16493__A (.DIODE(_02967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16472__A (.DIODE(_02967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16491__S (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16489__S (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16487__S (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16485__S (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16483__S (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16481__S (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16479__S (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16477__S (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16475__S (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16473__S (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16512__S (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16510__S (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16508__S (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16506__S (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16504__S (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16502__S (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16500__S (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16498__S (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16496__S (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16494__S (.DIODE(_02979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16533__S (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16531__S (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16529__S (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16527__S (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16525__S (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16523__S (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16521__S (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16519__S (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16517__S (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16515__S (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16605__S (.DIODE(_03003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16603__S (.DIODE(_03003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16582__A (.DIODE(_03003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16561__A (.DIODE(_03003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16540__A (.DIODE(_03003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16559__S (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16557__S (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16555__S (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16553__S (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16551__S (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16549__S (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16547__S (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16545__S (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16543__S (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16541__S (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16580__S (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16578__S (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16576__S (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16574__S (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16572__S (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16570__S (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16568__S (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16566__S (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16564__S (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16562__S (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16601__S (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16599__S (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16597__S (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16595__S (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16593__S (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16591__S (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16589__S (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16587__S (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16585__S (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16583__S (.DIODE(_03026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16673__S (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16671__S (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16650__A (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16629__A (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16608__A (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16627__S (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16625__S (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16623__S (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16621__S (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16619__S (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16617__S (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16615__S (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16613__S (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16611__S (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16609__S (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16648__S (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16646__S (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16644__S (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16642__S (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16640__S (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16638__S (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16636__S (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16634__S (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16632__S (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16630__S (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16669__S (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16667__S (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16665__S (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16663__S (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16661__S (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16659__S (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16657__S (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16655__S (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16653__S (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16651__S (.DIODE(_03062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16741__S (.DIODE(_03075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16739__S (.DIODE(_03075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16718__A (.DIODE(_03075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16697__A (.DIODE(_03075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16676__A (.DIODE(_03075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16695__S (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16693__S (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16691__S (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16689__S (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16687__S (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16685__S (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16683__S (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16681__S (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16679__S (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16677__S (.DIODE(_03076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16716__S (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16714__S (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16712__S (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16710__S (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16708__S (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16706__S (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16704__S (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16702__S (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16700__S (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16698__S (.DIODE(_03087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16737__S (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16735__S (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16733__S (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16731__S (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16729__S (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16727__S (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16725__S (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16723__S (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16721__S (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16719__S (.DIODE(_03098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16769__S (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16767__S (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16765__S (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16763__S (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16761__S (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16759__S (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16757__S (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16755__S (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16753__S (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16751__S (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16790__S (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16788__S (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16786__S (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16784__S (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16782__S (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16780__S (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16778__S (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16776__S (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16774__S (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16772__S (.DIODE(_03127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16811__S (.DIODE(_03138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16809__S (.DIODE(_03138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16807__S (.DIODE(_03138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16805__S (.DIODE(_03138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16803__S (.DIODE(_03138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16801__S (.DIODE(_03138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16799__S (.DIODE(_03138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16797__S (.DIODE(_03138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16795__S (.DIODE(_03138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16793__S (.DIODE(_03138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16837__S (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16835__S (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16833__S (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16831__S (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16829__S (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16827__S (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16825__S (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16823__S (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16821__S (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16819__S (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16858__S (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16856__S (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16854__S (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16852__S (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16850__S (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16848__S (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16846__S (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16844__S (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16842__S (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16840__S (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16879__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16877__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16875__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16873__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16871__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16869__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16867__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16865__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16863__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16861__S (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__C (.DIODE(_03191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08407__A_N (.DIODE(_03191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14682__A1 (.DIODE(_03195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14607__A1 (.DIODE(_03195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__A (.DIODE(_03195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__A3 (.DIODE(_03195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__A (.DIODE(_03195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__A (.DIODE(_03195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__B1 (.DIODE(_03195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15954__A (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14897__A (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14195__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__A (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08510__B (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08504__A_N (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__A (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08452__A (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__D1 (.DIODE(_03196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16117__A2 (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16114__A1 (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15646__A1 (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11355__A (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08867__A (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__A1 (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__A3 (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__B2 (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09028__A (.DIODE(_03206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__A_N (.DIODE(_03206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__B_N (.DIODE(_03206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__A (.DIODE(_03206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__B_N (.DIODE(_03206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08444__A (.DIODE(_03206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__A (.DIODE(_03206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16249__A1 (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16083__A (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11366__B (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__B (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09028__B_N (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__B (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__A (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09022__B (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__A (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__B (.DIODE(_03213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16210__C (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16084__B2 (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15840__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11368__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11354__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__A2 (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16213__A1 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16203__A (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16117__A1 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15958__B (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15648__A1 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__A2 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08499__A (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__A1 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__B (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__A1 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15958__C (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__S (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__S (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11326__S (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11320__S (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__S (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__S (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__A (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__A2 (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__A (.DIODE(_03225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__B2 (.DIODE(_03225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__B2 (.DIODE(_03225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__B1 (.DIODE(_03225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09732__B2 (.DIODE(_03225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__B2 (.DIODE(_03225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__B2 (.DIODE(_03225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09616__B2 (.DIODE(_03225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__B2 (.DIODE(_03225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__A (.DIODE(_03225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15795__A2 (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15787__C1 (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__B2 (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__B2 (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__B2 (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__B2 (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__B2 (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__A1 (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09314__A1 (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08490__A1 (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15961__C (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__S (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__S (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09066__S (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__S (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__S (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__A (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__S (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__B1 (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__A1 (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16090__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15985__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__A2 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11338__A (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__A (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__B (.DIODE(_03229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15634__B (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__B (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__B (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__A3 (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__B (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__B (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15856__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15645__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14747__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14743__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14086__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14012__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08508__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08502__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08456__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15694__B1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15671__B1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15031__B1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15017__A (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14991__A (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14878__B1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14780__B1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14689__A (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14188__B1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__A (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__B1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__B (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__B1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__B1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__B1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__B1 (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__A (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__B1 (.DIODE(_03253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__B2 (.DIODE(_03253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__B2 (.DIODE(_03253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__A (.DIODE(_03253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__A (.DIODE(_03253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__C_N (.DIODE(_03253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15636__B (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08614__B (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__A2 (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__A (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16107__A2 (.DIODE(_03255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__D (.DIODE(_03255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15630__S (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15549__S (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15495__S (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15045__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__C1 (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__C (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13353__B (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13322__B (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08643__B (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08492__A (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13788__C1 (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13779__A1 (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13730__A (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13631__A1 (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13570__B1 (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13561__A1 (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13498__A (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13477__A1 (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__A1 (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__A (.DIODE(_03275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13749__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13722__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13662__A (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13606__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13530__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13405__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13392__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13375__A1 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08518__A2 (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__A (.DIODE(_03276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15914__A (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15637__C1 (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15074__A (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__B (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11469__A (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__A (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__A (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A1 (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__A (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08498__A (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16263__B1 (.DIODE(_03292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15795__A1 (.DIODE(_03292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15790__A2 (.DIODE(_03292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15789__A2 (.DIODE(_03292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13875__A (.DIODE(_03292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08510__A (.DIODE(_03292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14649__A1 (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14596__A (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14534__A (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14408__B2 (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14278__A (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14190__A (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__B1 (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__B (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__A (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14679__A1 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14656__A1 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14635__A1 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14561__A1 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14412__A1 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14340__A1 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14275__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14239__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14206__A (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08512__C1 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__B2 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__B2 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__B2 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__B2 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__B2 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__B2 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B2 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__B2 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__A1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__A1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15783__A1 (.DIODE(_03298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15780__A2 (.DIODE(_03298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15637__A1 (.DIODE(_03298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14966__B (.DIODE(_03298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14195__A (.DIODE(_03298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13872__B (.DIODE(_03298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__A (.DIODE(_03298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__B2 (.DIODE(_03298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__A1 (.DIODE(_03298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08518__A1 (.DIODE(_03298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15661__A (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15651__A (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15643__B2 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15074__B (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14970__A (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13873__A (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__C1 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__C1 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__A (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__A (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15793__A (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__C1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__C1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__C1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__C1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__C1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__C1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__B2 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__C1 (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__A (.DIODE(_03302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15032__A1 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15030__A1 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15024__A1 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15022__A1 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14996__A1 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__A1 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09994__B2 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__C1 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__C1 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__A1 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15897__A (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15862__B (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14799__A (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14712__A (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14070__A (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14016__A (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13957__A (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__C1 (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08620__A1 (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__A (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15950__A (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15855__A (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15795__C1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__C (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11447__A (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__A (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11421__A (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__C (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__C1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__A1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__B (.DIODE(_03308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__A2 (.DIODE(_03308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__B1 (.DIODE(_03308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16107__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16095__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16045__B2 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15862__A (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15858__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15647__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__A (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13683__B1 (.DIODE(_03311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13668__B1 (.DIODE(_03311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13612__B1 (.DIODE(_03311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13584__B1 (.DIODE(_03311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13509__B1 (.DIODE(_03311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13346__B1 (.DIODE(_03311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08865__A (.DIODE(_03311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__B (.DIODE(_03311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13951__A1 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A2 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08545__A (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13898__A1 (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__A2 (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08545__B (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13895__A1 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11560__A2 (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08545__C (.DIODE(_03322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13907__A1 (.DIODE(_03323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11595__A2 (.DIODE(_03323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08545__D (.DIODE(_03323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13885__A1 (.DIODE(_03326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11530__B1 (.DIODE(_03326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__B (.DIODE(_03326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13892__A1 (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__A2 (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__C (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13931__A1 (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__A2 (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__A (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13912__A1 (.DIODE(_03333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11605__A2 (.DIODE(_03333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__D (.DIODE(_03333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13915__A1 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11618__A2 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__A (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13937__A1 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__A2 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__B (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13879__A1 (.DIODE(_03338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__B1 (.DIODE(_03338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__D (.DIODE(_03338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__A1 (.DIODE(_03340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13888__A1 (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__B1 (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__D (.DIODE(_03344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13948__A1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__A2 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__A (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13934__A1 (.DIODE(_03348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11673__A2 (.DIODE(_03348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__C (.DIODE(_03348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13901__A1 (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__A2 (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__D (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13882__A1 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11516__B1 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__A (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__A1 (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__A2 (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__B (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13925__A1 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__A2 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__C (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13928__A1 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__A2 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__A (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13918__A1 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11629__A2 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__B (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13940__A1 (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11691__A2 (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__C (.DIODE(_03358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13904__A1 (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__A2 (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__D (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__A2 (.DIODE(_03361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15785__B (.DIODE(_03364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15640__B1 (.DIODE(_03364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14454__A (.DIODE(_03364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14315__B1 (.DIODE(_03364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14310__A (.DIODE(_03364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12737__A (.DIODE(_03364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08592__C_N (.DIODE(_03364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__A3 (.DIODE(_03364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15792__C (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14495__A1 (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14442__B1 (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14400__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14394__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14383__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14369__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14358__A1 (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14295__B (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08592__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14608__B2 (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14597__B2 (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14408__A1 (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14400__B (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14383__B (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14359__A (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15640__A1 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14595__A1 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14362__A (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14308__A (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__B (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15787__A1 (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__A2 (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__A (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__A (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__A1 (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__A (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__C (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__A1 (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__B (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__A (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15789__A1 (.DIODE(_03385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10272__B2 (.DIODE(_03385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09994__A1 (.DIODE(_03385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__B2 (.DIODE(_03385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09883__A1 (.DIODE(_03385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__B2 (.DIODE(_03385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09733__A1 (.DIODE(_03385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__A (.DIODE(_03385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A1 (.DIODE(_03385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__A2 (.DIODE(_03385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15072__B1 (.DIODE(_03387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14893__B2 (.DIODE(_03387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13604__A1_N (.DIODE(_03387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13575__A (.DIODE(_03387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13475__A (.DIODE(_03387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13460__A (.DIODE(_03387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13367__A1_N (.DIODE(_03387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13345__A1_N (.DIODE(_03387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08621__B (.DIODE(_03387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08613__B (.DIODE(_03387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__B (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08620__B1 (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__A1 (.DIODE(_03407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__A1 (.DIODE(_03407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__A1 (.DIODE(_03407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__A1 (.DIODE(_03407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__A1 (.DIODE(_03407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__A1 (.DIODE(_03407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__A1 (.DIODE(_03407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__A1 (.DIODE(_03407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__A1 (.DIODE(_03407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08640__A1 (.DIODE(_03407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__A (.DIODE(_03412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11426__A (.DIODE(_03412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__A (.DIODE(_03412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__A (.DIODE(_03412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__A2 (.DIODE(_03412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15765__B (.DIODE(_03425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__C_N (.DIODE(_03425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11487__B (.DIODE(_03428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__B (.DIODE(_03428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__B (.DIODE(_03428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__B (.DIODE(_03428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11479__B (.DIODE(_03428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__B (.DIODE(_03428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__B (.DIODE(_03428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__B (.DIODE(_03428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11471__B (.DIODE(_03428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__A2 (.DIODE(_03428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__A1 (.DIODE(_03460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__A2 (.DIODE(_03460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__A1 (.DIODE(_03475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__A2 (.DIODE(_03475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__A (.DIODE(_03509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08746__A (.DIODE(_03509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13540__A1 (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13495__A1 (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13487__A (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__A3 (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10788__A1 (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__A0 (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A3 (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__A (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08786__A2 (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__B (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13465__A (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10788__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__A1 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A0 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__A (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08848__B (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08782__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__A1 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13435__A (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A2 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10743__A1 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__A0 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A3 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A0 (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__A (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__B_N (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__B (.DIODE(_03524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13687__A (.DIODE(_03575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13615__A (.DIODE(_03575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__A1 (.DIODE(_03575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08810__B (.DIODE(_03575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08862__S (.DIODE(_03599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08834__A2 (.DIODE(_03599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__B (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__C (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__A_N (.DIODE(_03604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__C (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15784__A (.DIODE(_03630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15647__A3 (.DIODE(_03630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__B2 (.DIODE(_03630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__A1_N (.DIODE(_03630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14891__A (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13800__A (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13761__A1 (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13703__A1 (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13645__A1 (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13547__B1 (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13489__B1 (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13453__B1 (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13430__A1 (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__D (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16105__S (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16101__A1 (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16085__S (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16004__A1 (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15976__S (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15877__S (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15844__S (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15823__S (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__A (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__A (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16093__A2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16000__A2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15996__A2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15990__A1 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15969__A2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15822__B2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__A2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11378__A2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11358__A2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__B2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16743__B2 (.DIODE(_03638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__A1 (.DIODE(_03638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__A1 (.DIODE(_03638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__A1 (.DIODE(_03638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__A1 (.DIODE(_03638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__A1 (.DIODE(_03638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__B2 (.DIODE(_03638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__A1 (.DIODE(_03638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__A2 (.DIODE(_03638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08917__A1 (.DIODE(_03638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15610__S1 (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15547__A1 (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15520__S1 (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15493__A1 (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15326__S1 (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15314__B1 (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15197__C1 (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15166__A (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15128__S1 (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08912__A1 (.DIODE(_03639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15625__S0 (.DIODE(_03640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15624__S0 (.DIODE(_03640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15544__S0 (.DIODE(_03640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15490__S0 (.DIODE(_03640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15423__S0 (.DIODE(_03640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15404__S0 (.DIODE(_03640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15202__S0 (.DIODE(_03640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__A (.DIODE(_03640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08880__A (.DIODE(_03640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08876__A (.DIODE(_03640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15602__S0 (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15601__S0 (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15587__S0 (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15586__S0 (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15381__S0 (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__S0 (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08931__S0 (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08922__S0 (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__S0 (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__S0 (.DIODE(_03641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15625__S1 (.DIODE(_03642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15624__S1 (.DIODE(_03642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15544__S1 (.DIODE(_03642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15543__S1 (.DIODE(_03642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15490__S1 (.DIODE(_03642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15423__S1 (.DIODE(_03642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15404__S1 (.DIODE(_03642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15202__S1 (.DIODE(_03642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15136__A (.DIODE(_03642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08878__A (.DIODE(_03642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15400__S1 (.DIODE(_03643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15198__S1 (.DIODE(_03643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15160__A (.DIODE(_03643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__S1 (.DIODE(_03643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__S1 (.DIODE(_03643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08945__S1 (.DIODE(_03643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08944__S1 (.DIODE(_03643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08886__S1 (.DIODE(_03643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__S1 (.DIODE(_03643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__S1 (.DIODE(_03643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15622__S0 (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15621__S0 (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15541__S0 (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15540__S0 (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15487__S0 (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15486__S0 (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15420__S0 (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15401__S0 (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15199__S0 (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__S0 (.DIODE(_03645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15194__A (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15092__S1 (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15091__S1 (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15088__S1 (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15084__S1 (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15083__S1 (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15080__S1 (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15078__A (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__A (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08882__A (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15622__S1 (.DIODE(_03647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15541__S1 (.DIODE(_03647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15414__S1 (.DIODE(_03647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15191__S1 (.DIODE(_03647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15169__A (.DIODE(_03647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15145__A (.DIODE(_03647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15142__A (.DIODE(_03647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15131__A (.DIODE(_03647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15087__S1 (.DIODE(_03647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__S1 (.DIODE(_03647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15419__S0 (.DIODE(_03649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15400__S0 (.DIODE(_03649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15198__S0 (.DIODE(_03649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15176__A (.DIODE(_03649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__S0 (.DIODE(_03649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__S0 (.DIODE(_03649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08945__S0 (.DIODE(_03649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08944__S0 (.DIODE(_03649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08886__S0 (.DIODE(_03649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__S0 (.DIODE(_03649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15619__S (.DIODE(_03653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15538__S (.DIODE(_03653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15488__S (.DIODE(_03653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15484__S (.DIODE(_03653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15421__S (.DIODE(_03653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15398__S (.DIODE(_03653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15393__A (.DIODE(_03653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15158__A (.DIODE(_03653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15147__A (.DIODE(_03653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08890__S0 (.DIODE(_03653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15620__C1 (.DIODE(_03654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15425__A1 (.DIODE(_03654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15295__B1 (.DIODE(_03654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15242__B1 (.DIODE(_03654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15204__A1 (.DIODE(_03654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15113__A (.DIODE(_03654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15063__C1 (.DIODE(_03654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15053__C1 (.DIODE(_03654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__A (.DIODE(_03654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08890__S1 (.DIODE(_03654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15627__B1 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15546__B1 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15492__B1 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15406__B1 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15067__A1 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15057__A1 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08952__A1 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08937__A1 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__A1 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__A1 (.DIODE(_03657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15378__A (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15055__S0 (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15054__S0 (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15051__S0 (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__S0 (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08934__S0 (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__S0 (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__S0 (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08902__S0 (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__S0 (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15379__A (.DIODE(_03659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15055__S1 (.DIODE(_03659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15054__S1 (.DIODE(_03659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15051__S1 (.DIODE(_03659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__S1 (.DIODE(_03659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08934__S1 (.DIODE(_03659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__S1 (.DIODE(_03659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__S1 (.DIODE(_03659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08902__S1 (.DIODE(_03659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__S1 (.DIODE(_03659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15543__S0 (.DIODE(_03661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15489__S0 (.DIODE(_03661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15422__S0 (.DIODE(_03661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15403__S0 (.DIODE(_03661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15201__S0 (.DIODE(_03661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__S0 (.DIODE(_03661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08958__S0 (.DIODE(_03661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__S0 (.DIODE(_03661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__S0 (.DIODE(_03661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08898__S0 (.DIODE(_03661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15489__S1 (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15422__S1 (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15403__S1 (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15201__S1 (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__S1 (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08958__S1 (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__S1 (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__S1 (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08920__A (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08898__S1 (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15413__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15260__A (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15190__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15066__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15056__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15047__A (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08936__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__A1 (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08900__S (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15626__S (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15417__A (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15203__S (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15134__A (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15089__A (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15062__A (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15052__A (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08946__A (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__A (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__A (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15193__A (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15140__A (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15092__S0 (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15091__S0 (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15088__S0 (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15084__S0 (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15083__S0 (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15080__S0 (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15077__A (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__A (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15412__S0 (.DIODE(_03670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15411__S0 (.DIODE(_03670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15189__S0 (.DIODE(_03670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15188__S0 (.DIODE(_03670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15065__S0 (.DIODE(_03670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15064__S0 (.DIODE(_03670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15061__S0 (.DIODE(_03670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15058__A (.DIODE(_03670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15048__A (.DIODE(_03670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__S0 (.DIODE(_03670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15412__S1 (.DIODE(_03671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15411__S1 (.DIODE(_03671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15189__S1 (.DIODE(_03671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15188__S1 (.DIODE(_03671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15065__S1 (.DIODE(_03671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15064__S1 (.DIODE(_03671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15061__S1 (.DIODE(_03671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15059__A (.DIODE(_03671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15049__A (.DIODE(_03671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__S1 (.DIODE(_03671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15481__B1 (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15163__A (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15094__B1 (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08910__A (.DIODE(_03674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15620__B2 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15546__A1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15492__A1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15425__B1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15204__B1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15149__A (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15067__B1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__B1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08937__B1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__C1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15104__A1 (.DIODE(_03677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08916__A1 (.DIODE(_03677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15100__B (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15096__A (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15069__A (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__A (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__A (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08916__A2 (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16745__A (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__A1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__A1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__A1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__A1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__A1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__A1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__A1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08916__B1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15458__B2 (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15450__S1 (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15362__A1 (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15350__B2 (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15291__S1 (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15283__B2 (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__A1 (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__A1 (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A1 (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__A1 (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15602__S1 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15601__S1 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15587__S1 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15586__S1 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15381__S1 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15177__A (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__S1 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08931__S1 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08922__S1 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__S1 (.DIODE(_03684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15578__A (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15574__S (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15522__A (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15473__S (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15441__A (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15256__S (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15245__S (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15225__S (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__S (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08924__S (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15559__B1 (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15485__B2 (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15470__B1 (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15418__C1 (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15406__A1 (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15183__A (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15139__B1 (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15057__B1 (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08952__B1 (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__B1 (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15108__A2 (.DIODE(_03703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__A2 (.DIODE(_03703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15623__S (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15614__A (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15542__S (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15533__A (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15479__A (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15395__A1 (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15214__A (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15196__A (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15082__A1 (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__S (.DIODE(_03709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15545__S (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15491__S (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15424__S (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15405__S (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15093__S (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15085__S (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15081__A (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__S (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08956__A (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__S (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15616__A1 (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15535__A1 (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15481__A1 (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15415__A1 (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15402__S (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15200__S (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15192__A1 (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15129__A (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15090__A1 (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__S (.DIODE(_03719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15111__A2 (.DIODE(_03726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__B1 (.DIODE(_03726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16200__A (.DIODE(_03730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09206__A (.DIODE(_03730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__A1 (.DIODE(_03730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__A2 (.DIODE(_03730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09045__S (.DIODE(_03730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__S (.DIODE(_03730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09040__S (.DIODE(_03730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__S (.DIODE(_03730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__S (.DIODE(_03730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__S (.DIODE(_03730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16096__A2 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__D (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__A2 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__D (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__B2 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__B1 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09176__A (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__A1 (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09110__A (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__A (.DIODE(_03736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15988__A2 (.DIODE(_03737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15823__A1 (.DIODE(_03737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15821__B (.DIODE(_03737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A1 (.DIODE(_03737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__A1 (.DIODE(_03737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__B1 (.DIODE(_03737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__A1 (.DIODE(_03737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__B2 (.DIODE(_03737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09088__A2 (.DIODE(_03737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__A1 (.DIODE(_03737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15982__A1 (.DIODE(_03743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__A (.DIODE(_03743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__C_N (.DIODE(_03743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09097__A1 (.DIODE(_03743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09082__A (.DIODE(_03743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__A (.DIODE(_03743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09006__A (.DIODE(_03743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__A (.DIODE(_03743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16097__A1 (.DIODE(_03747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15826__B1 (.DIODE(_03747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__A1 (.DIODE(_03747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09181__A2 (.DIODE(_03747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09020__A (.DIODE(_03747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09006__B (.DIODE(_03747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__A (.DIODE(_03747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15836__B1 (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__A (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A1 (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15959__A1 (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__S (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__S (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09248__S (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__S (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__S (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09193__S (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__S (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__A (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__S (.DIODE(_03757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16096__A1 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__B (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__A (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09175__A (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09065__A (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09014__A (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__A (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16004__A2 (.DIODE(_03763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15999__B1 (.DIODE(_03763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15805__B (.DIODE(_03763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11420__A2 (.DIODE(_03763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__B1_N (.DIODE(_03763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09258__B1 (.DIODE(_03763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__A1 (.DIODE(_03763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__A1 (.DIODE(_03763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09149__A1 (.DIODE(_03763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09016__A2 (.DIODE(_03763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16084__A1 (.DIODE(_03767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15987__A1 (.DIODE(_03767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15980__A2 (.DIODE(_03767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11399__A1 (.DIODE(_03767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__A2 (.DIODE(_03767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__A (.DIODE(_03767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09125__B2 (.DIODE(_03767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A (.DIODE(_03767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09007__A (.DIODE(_03767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16097__A2 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16092__A1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15828__B1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11394__A (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__A (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__B1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__A (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__A1 (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09082__B (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09020__B (.DIODE(_03781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16247__A1 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16102__A1 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16091__D (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15981__A (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__A (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11366__A (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__A (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__A (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09087__A1 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09022__A (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16253__A1 (.DIODE(_03810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15848__A2 (.DIODE(_03810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__A3 (.DIODE(_03810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__A2 (.DIODE(_03810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__B2 (.DIODE(_03810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09113__B1 (.DIODE(_03810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09053__A (.DIODE(_03810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15990__A2 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15811__C (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__A1 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__B2 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__A1 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09065__C (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16002__A1 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15995__B2 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15816__A1 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__A1 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A1 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09204__B2 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__A1 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09065__D (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11314__A (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__A (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__A (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__A (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11277__A (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__B (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__B (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__B (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__A (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__A (.DIODE(_03841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16251__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15987__B1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15848__A3 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15840__C (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15809__C (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__B (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A2 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__A1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__B1 (.DIODE(_03864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15994__A1 (.DIODE(_03867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15819__A1 (.DIODE(_03867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__A1 (.DIODE(_03867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__B1 (.DIODE(_03867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__C_N (.DIODE(_03867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11398__A1 (.DIODE(_03867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__A2 (.DIODE(_03867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__B1 (.DIODE(_03867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__A2 (.DIODE(_03867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09108__B_N (.DIODE(_03867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11364__A3 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__A2 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__A1 (.DIODE(_03874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16259__A1 (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16091__A_N (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15839__A_N (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15813__C (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__B (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__A1 (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__C (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__A1 (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09148__B1 (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__A1 (.DIODE(_03878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15995__A2 (.DIODE(_03880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15993__B1 (.DIODE(_03880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15987__B2 (.DIODE(_03880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11398__B2 (.DIODE(_03880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09213__B (.DIODE(_03880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09149__A2 (.DIODE(_03880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__A3 (.DIODE(_03880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__A2 (.DIODE(_03880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16255__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16101__A3 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15995__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15843__B (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15839__B (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11369__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__B (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09204__A1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__B2 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09128__B1 (.DIODE(_03885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__B2 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09254__B2 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09246__B2 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__B2 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__B2 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__B2 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09191__B2 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__B2 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__B2 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__B2 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16098__C1 (.DIODE(_03891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15980__A1 (.DIODE(_03891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15827__B1 (.DIODE(_03891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__A1 (.DIODE(_03891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A (.DIODE(_03891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__A1 (.DIODE(_03891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09193__A1 (.DIODE(_03891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09181__A1 (.DIODE(_03891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__A1 (.DIODE(_03891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09137__A (.DIODE(_03891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15998__B1 (.DIODE(_03892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15817__A1 (.DIODE(_03892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__A1 (.DIODE(_03892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__B (.DIODE(_03892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09266__A1 (.DIODE(_03892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09260__A1 (.DIODE(_03892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__B (.DIODE(_03892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__A1 (.DIODE(_03892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09175__B (.DIODE(_03892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__A2 (.DIODE(_03892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16257__A1 (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15839__C (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15804__B1 (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__A1 (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__A1 (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A1 (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__A1 (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__A1 (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09141__A1 (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__B1 (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15829__B1 (.DIODE(_03910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__B (.DIODE(_03910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09157__A1 (.DIODE(_03910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16098__A3 (.DIODE(_03916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15982__A2 (.DIODE(_03916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15875__B (.DIODE(_03916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15837__B (.DIODE(_03916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11400__A2 (.DIODE(_03916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A (.DIODE(_03916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09195__A (.DIODE(_03916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09187__B (.DIODE(_03916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09179__A (.DIODE(_03916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09164__A (.DIODE(_03916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15834__C (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__A2 (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__A1 (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16092__A2 (.DIODE(_03935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16084__A2 (.DIODE(_03935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09213__A (.DIODE(_03935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__A (.DIODE(_03935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16052__B2 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15900__A_N (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15896__B (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15872__C (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15870__C (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15867__B (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15865__C_N (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15861__A (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15854__C (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09193__A0 (.DIODE(_03940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15810__B1 (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11390__A (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__A1 (.DIODE(_03954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15974__A (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15812__B1 (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__C_N (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__A1 (.DIODE(_03965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15974__D_N (.DIODE(_03977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15814__B1 (.DIODE(_03977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__A (.DIODE(_03977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__A1 (.DIODE(_03977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15840__B (.DIODE(_03979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__B (.DIODE(_03979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__A (.DIODE(_03979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__A1_N (.DIODE(_03979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15816__B2 (.DIODE(_03987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11390__B (.DIODE(_03987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09248__A1 (.DIODE(_03987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15817__B2 (.DIODE(_03994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__B (.DIODE(_03994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__A1 (.DIODE(_03994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15819__B2 (.DIODE(_04000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__C (.DIODE(_04000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__A1 (.DIODE(_04000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15783__A2 (.DIODE(_04006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15649__C (.DIODE(_04006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__A2 (.DIODE(_04006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__A2 (.DIODE(_04006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09270__A (.DIODE(_04006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10169__A2 (.DIODE(_04008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__A2 (.DIODE(_04008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__A2 (.DIODE(_04008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__A2 (.DIODE(_04008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__A2 (.DIODE(_04008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__B1 (.DIODE(_04008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__B1 (.DIODE(_04008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__B1 (.DIODE(_04008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__A2 (.DIODE(_04008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A2 (.DIODE(_04008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__A1 (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__B1 (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__B1 (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__B1 (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__B1 (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__B1 (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__A (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__B1 (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__B1 (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__A (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__A1 (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__A1 (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10301__A1 (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__A1 (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__B2 (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__A1 (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09724__A1 (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__A1 (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__A1 (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__A1 (.DIODE(_04010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__A2 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10209__B1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10070__B1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__B1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09819__A2 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__A2 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09668__B1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__A2 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09411__A (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15946__A1 (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__A2 (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__A2 (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__A2 (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__B1 (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__A2 (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10039__A2 (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09848__B1 (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A2 (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A2 (.DIODE(_04012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__B2 (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__B1 (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__B2 (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__B1 (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09820__B2 (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__A2 (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__B1 (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__A2 (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__B2 (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__A (.DIODE(_04013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__B1 (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__B1 (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10131__A2 (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__A2 (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09986__B2 (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__B1 (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09702__B2 (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__A2 (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__A2 (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__B2 (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10209__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10175__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09608__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09279__A (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15947__A1 (.DIODE(_04016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10413__A2 (.DIODE(_04016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10280__A2 (.DIODE(_04016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__A2 (.DIODE(_04016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09986__A2 (.DIODE(_04016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09848__A2 (.DIODE(_04016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09820__A2 (.DIODE(_04016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09702__A2 (.DIODE(_04016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__A2 (.DIODE(_04016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__A2 (.DIODE(_04016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__B1 (.DIODE(_04017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__B1 (.DIODE(_04017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10175__B1 (.DIODE(_04017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__B1 (.DIODE(_04017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__A1 (.DIODE(_04017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09819__B1 (.DIODE(_04017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__A1 (.DIODE(_04017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__B1 (.DIODE(_04017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__B1 (.DIODE(_04017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A (.DIODE(_04017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15943__A1 (.DIODE(_04018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__A1 (.DIODE(_04018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__A1 (.DIODE(_04018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__A1 (.DIODE(_04018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__A1 (.DIODE(_04018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__A1 (.DIODE(_04018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__B1 (.DIODE(_04018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__A1 (.DIODE(_04018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__A1 (.DIODE(_04018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__B1 (.DIODE(_04018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__A2 (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__A2 (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10060__A2 (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__A2 (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09911__A2 (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__A2 (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__A2 (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__A2 (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__A2 (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__A (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15973__B2 (.DIODE(_04022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15032__A2 (.DIODE(_04022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15030__A2 (.DIODE(_04022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15024__A2 (.DIODE(_04022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15022__A2 (.DIODE(_04022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14996__A2 (.DIODE(_04022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09984__A2 (.DIODE(_04022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A2 (.DIODE(_04022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__A2 (.DIODE(_04022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__A2 (.DIODE(_04022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__B2 (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__B2 (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__B2 (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10060__B2 (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__B2 (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__B2 (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09688__B2 (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__B2 (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09578__B2 (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__A (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15979__A1 (.DIODE(_04024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15661__B (.DIODE(_04024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__B2 (.DIODE(_04024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__B2 (.DIODE(_04024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09984__B2 (.DIODE(_04024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__B2 (.DIODE(_04024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__B2 (.DIODE(_04024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__B2 (.DIODE(_04024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__B2 (.DIODE(_04024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__B2 (.DIODE(_04024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__C1 (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__C1 (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__C1 (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__C1 (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10060__C1 (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__C1 (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09688__C1 (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__C1 (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09578__C1 (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09290__A (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__C1 (.DIODE(_04027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__C1 (.DIODE(_04027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__C1 (.DIODE(_04027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10020__C1 (.DIODE(_04027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09984__C1 (.DIODE(_04027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__C1 (.DIODE(_04027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__C1 (.DIODE(_04027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__C1 (.DIODE(_04027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__C1 (.DIODE(_04027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__C1 (.DIODE(_04027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13368__A0 (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13363__A (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__A3 (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__A1 (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__A0 (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09614__A (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__A (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09467__A (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13412__A1 (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13365__A1 (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13359__A0 (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13347__A1 (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13346__A1 (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__A2 (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__A (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__A (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__B1 (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09306__A (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__A1 (.DIODE(_04038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__A1 (.DIODE(_04038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A1 (.DIODE(_04038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__A1 (.DIODE(_04038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__A1 (.DIODE(_04038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__A1 (.DIODE(_04038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A1 (.DIODE(_04038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__B (.DIODE(_04038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__B (.DIODE(_04038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09306__B (.DIODE(_04038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13387__A0 (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__A2 (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__A0 (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__A2 (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09532__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__S (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__A (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__A1 (.DIODE(_04040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13376__A0 (.DIODE(_04040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13361__A (.DIODE(_04040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__A1 (.DIODE(_04040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__A1 (.DIODE(_04040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__A1_N (.DIODE(_04040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__A1 (.DIODE(_04040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__A (.DIODE(_04040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__S (.DIODE(_04040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__S (.DIODE(_04040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09314__A2 (.DIODE(_04043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16746__B1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__A1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__A1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__A1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__A1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__A1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__B1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__A1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09616__A1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__B2 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__A2 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10272__A2 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A2 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A2 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__A2 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__A2 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__A2 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__C1 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__C1 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09314__C1 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__B2 (.DIODE(_04050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__A (.DIODE(_04051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A (.DIODE(_04051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09983__A (.DIODE(_04051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__A (.DIODE(_04051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A (.DIODE(_04051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__A (.DIODE(_04051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__A (.DIODE(_04051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__A (.DIODE(_04051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__A (.DIODE(_04051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09367__A (.DIODE(_04051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10396__A1 (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__A1 (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__A (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__B2 (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09598__A (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__A (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__A1 (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__B2 (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__A1 (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__A (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__A1 (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__A1 (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__A1 (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__B2 (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__A1 (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__A1 (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__A (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09439__A (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A1 (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09319__A (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13339__A1 (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10430__A1 (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__A (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__A1 (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__A (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__A1 (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__A (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09750__A (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__A (.DIODE(_04054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10323__S0 (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10322__S0 (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__A (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09559__A (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__A (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__A (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__A (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__S0 (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__S0 (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09321__A (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__S0 (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09682__S0 (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__S0 (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09674__S0 (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__S0 (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__S0 (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__S0 (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__S0 (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__S0 (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09322__A (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__S0 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__S0 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__S0 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__S0 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__S0 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__S0 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__S0 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09974__S0 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__S0 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__S0 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10323__S1 (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10322__S1 (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__S1 (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__S1 (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09405__S1 (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__A (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__S1 (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__S1 (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__S1 (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__S1 (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__S1 (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__S1 (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__S1 (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__S1 (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__S1 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__S1 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__S1 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__S1 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__S1 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__S1 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__S1 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09974__S1 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__S1 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__S1 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__S (.DIODE(_04063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__A (.DIODE(_04063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__A (.DIODE(_04063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__S (.DIODE(_04063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__A (.DIODE(_04063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__A (.DIODE(_04063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10460__S (.DIODE(_04064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__S (.DIODE(_04064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10191__S (.DIODE(_04064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__S (.DIODE(_04064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__S (.DIODE(_04064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__S (.DIODE(_04064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09438__S (.DIODE(_04064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__A1 (.DIODE(_04064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__S (.DIODE(_04064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09330__A (.DIODE(_04064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__S (.DIODE(_04065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__S (.DIODE(_04065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__S (.DIODE(_04065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__S (.DIODE(_04065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__S (.DIODE(_04065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10048__S (.DIODE(_04065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__S (.DIODE(_04065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__S (.DIODE(_04065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09556__A (.DIODE(_04065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__S (.DIODE(_04065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__A1 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__A1 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__A1 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__B1 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09863__B1 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__A1 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09482__A (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__B1 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__C1 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09334__A (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10429__A1 (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__A1 (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__B1 (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A1 (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__B1 (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__A1 (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__A1 (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__A1 (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__C1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__A (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__S0 (.DIODE(_04071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10263__S0 (.DIODE(_04071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__S0 (.DIODE(_04071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__S0 (.DIODE(_04071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__S0 (.DIODE(_04071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__S0 (.DIODE(_04071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__S0 (.DIODE(_04071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__S0 (.DIODE(_04071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09394__S0 (.DIODE(_04071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__A (.DIODE(_04071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__S0 (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10006__S0 (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09716__S0 (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__S0 (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__S0 (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__S0 (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09475__A (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09388__S0 (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__S0 (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__S0 (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__S1 (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10263__S1 (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__S1 (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__S1 (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__S1 (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__S1 (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__S1 (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__S1 (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09394__S1 (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A (.DIODE(_04073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__S1 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10006__S1 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09716__S1 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__S1 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__S1 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__S1 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__A (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09388__S1 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__S1 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__S1 (.DIODE(_04074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10395__S (.DIODE(_04077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10317__S (.DIODE(_04077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10313__S (.DIODE(_04077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10264__S (.DIODE(_04077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09834__S (.DIODE(_04077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__S (.DIODE(_04077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__S (.DIODE(_04077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__S (.DIODE(_04077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A (.DIODE(_04077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__A (.DIODE(_04077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__S (.DIODE(_04078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__S (.DIODE(_04078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__S (.DIODE(_04078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09755__S (.DIODE(_04078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__S (.DIODE(_04078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09680__S (.DIODE(_04078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09672__S (.DIODE(_04078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__A (.DIODE(_04078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__S (.DIODE(_04078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__S (.DIODE(_04078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__A2 (.DIODE(_04079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__B1 (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__B1 (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__B1 (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__A (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10389__B1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__B1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__B1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__B1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09718__B1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__B1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09651__B1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__A (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__B1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__A (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10454__B1 (.DIODE(_04082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__B1 (.DIODE(_04082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__B1 (.DIODE(_04082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10049__B1 (.DIODE(_04082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__B1 (.DIODE(_04082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__B1 (.DIODE(_04082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09929__B1 (.DIODE(_04082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__A1 (.DIODE(_04082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__B1 (.DIODE(_04082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__B1 (.DIODE(_04082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__S0 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10311__S0 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10190__S0 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__S0 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09832__S0 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__A (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__A (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__S0 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__S0 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09350__A (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__S0 (.DIODE(_04085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10451__S0 (.DIODE(_04085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09927__S0 (.DIODE(_04085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__S0 (.DIODE(_04085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__S0 (.DIODE(_04085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__S0 (.DIODE(_04085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__S0 (.DIODE(_04085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__S0 (.DIODE(_04085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__S0 (.DIODE(_04085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__S0 (.DIODE(_04085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__S1 (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10311__S1 (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10190__S1 (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__S1 (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09832__S1 (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__A (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__S1 (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__S1 (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__S1 (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__A (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__S1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10451__S1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09927__S1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__S1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__S1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__S1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__S1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__S1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__S1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__S1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__S1 (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__S1 (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09682__S1 (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__S1 (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09674__S1 (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__S1 (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__A (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__S1 (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__S1 (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__S1 (.DIODE(_04091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__B1 (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10429__B1 (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__C1 (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__B1 (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__B1 (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__B1 (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__C1 (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__B1 (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__B1 (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__B1 (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap301_A (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09686__A (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__B1 (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__B1 (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__B1 (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__C1 (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__B1 (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__B1 (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09938__B1 (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__B1 (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__A (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__B1 (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__C1 (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15663__A1 (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14976__A (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13367__A2_N (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09367__B (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__A2 (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__A2 (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10129__A2 (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10070__A2 (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__A2 (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__A2 (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09668__A2 (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__A2 (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__A2 (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__A2 (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__B1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__A1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10280__B1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__A1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10129__B1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__B1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__B1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__A1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__B1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__A2 (.DIODE(_04112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__B2 (.DIODE(_04120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__S (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__S (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10056__S (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10012__S (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09972__S (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__S (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09928__S (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__S (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__S (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__A1 (.DIODE(_04121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10394__S0 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10393__S0 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10320__S0 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__S0 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__S0 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__A (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09405__S0 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__S0 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09400__S0 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09391__S0 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10394__S1 (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10393__S1 (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10320__S1 (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__S1 (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__S1 (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__A (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__A (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__S1 (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09400__S1 (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09391__S1 (.DIODE(_04124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__B1 (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__C1 (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10193__A (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10058__B1 (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__A (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__A (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__B1 (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14978__A (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13385__A (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__B (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10413__B1 (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__A2 (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__A2 (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__A2 (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__A2 (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__A2 (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__A2 (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__B1 (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__B1 (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__A2 (.DIODE(_04145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__C1 (.DIODE(_04149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__C1 (.DIODE(_04149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__C1 (.DIODE(_04149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__C1 (.DIODE(_04149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__C1 (.DIODE(_04149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__A1 (.DIODE(_04149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__C1 (.DIODE(_04149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__C1 (.DIODE(_04149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__C1 (.DIODE(_04149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__A (.DIODE(_04149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14968__B2 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__C1 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10301__C1 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__C1 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10029__A1 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__C1 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09724__C1 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__C1 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__C1 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09417__C1 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16207__A (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15792__A (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15790__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__B1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__B1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09887__B1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__A1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09462__B1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__B1 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__A2 (.DIODE(_04159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13393__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13368__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__A2 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__A1 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__A2 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__B1 (.DIODE(_04163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__A3 (.DIODE(_04164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__B2 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__A2 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10332__A2 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__B2 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10039__B2 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__A2 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__A2 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__A2 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__B1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__B1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15969__A1 (.DIODE(_04168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__A1 (.DIODE(_04168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__A1 (.DIODE(_04168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__A1 (.DIODE(_04168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__A1 (.DIODE(_04168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10021__A1 (.DIODE(_04168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A1 (.DIODE(_04168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__A1 (.DIODE(_04168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__A1 (.DIODE(_04168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__A1 (.DIODE(_04168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15672__A1 (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14981__A (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__A (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13400__A2 (.DIODE(_04186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__A2 (.DIODE(_04186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15651__B (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__B2 (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__B2 (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__B2 (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__B2 (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10020__B2 (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09911__B2 (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__B2 (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__B2 (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__B2 (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__C1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__C1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__C1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__C1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__C1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09911__C1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__C1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__C1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__C1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__C1 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__A2 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13415__A (.DIODE(_04198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13406__A0 (.DIODE(_04198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13387__A1 (.DIODE(_04198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__A1 (.DIODE(_04198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__A0 (.DIODE(_04198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__A0 (.DIODE(_04198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A2 (.DIODE(_04198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__A1 (.DIODE(_04198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__A3 (.DIODE(_04198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__A2 (.DIODE(_04198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__B1 (.DIODE(_04201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__C1 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__C1 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__C1 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__C1 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__C1 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__C1 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__B1 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__B1 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__C1 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__C1 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__A3 (.DIODE(_04203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10486__A1 (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__B2 (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10289__A1 (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__A (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__A (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09719__A1 (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__B2 (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09652__A1 (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__A1 (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__A (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13330__S0 (.DIODE(_04207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13329__S0 (.DIODE(_04207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__S0 (.DIODE(_04207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__S0 (.DIODE(_04207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__S0 (.DIODE(_04207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__S0 (.DIODE(_04207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__S0 (.DIODE(_04207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__S0 (.DIODE(_04207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__S0 (.DIODE(_04207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__S0 (.DIODE(_04207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13330__S1 (.DIODE(_04208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13329__S1 (.DIODE(_04208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__S1 (.DIODE(_04208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__S1 (.DIODE(_04208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__S1 (.DIODE(_04208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__S1 (.DIODE(_04208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__S1 (.DIODE(_04208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__S1 (.DIODE(_04208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__S1 (.DIODE(_04208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__S1 (.DIODE(_04208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13335__S (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13331__S (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__S (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10350__S (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__S (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10254__A1 (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__S (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A1 (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__S (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09480__S (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10397__A1 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10389__A1 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10293__B1 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__A1 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__A (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__A1 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09718__A1 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09651__A1 (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__A (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__A (.DIODE(_04214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13340__A1 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13332__A1 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A1 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__A1 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10147__A1 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10124__A1 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__A1 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__A (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09507__A1 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__A1 (.DIODE(_04215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10383__S0 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__S0 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10252__S0 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09897__S0 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__S0 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__S0 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__S0 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__S0 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__S0 (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09485__A (.DIODE(_04216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__S0 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__S0 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__S0 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__S0 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__S0 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09583__S0 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__S0 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__S0 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__S0 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__S0 (.DIODE(_04217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__S1 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__S1 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__S1 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__S1 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__S1 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__S1 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__S1 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__S1 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__S1 (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__A (.DIODE(_04218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__S1 (.DIODE(_04219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__S1 (.DIODE(_04219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__S1 (.DIODE(_04219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__S1 (.DIODE(_04219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__S1 (.DIODE(_04219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09583__S1 (.DIODE(_04219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__S1 (.DIODE(_04219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__S1 (.DIODE(_04219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__S1 (.DIODE(_04219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__S1 (.DIODE(_04219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10392__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10257__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09602__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__A (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10291__A (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10288__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09714__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09564__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__S (.DIODE(_04223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__A2 (.DIODE(_04224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13332__B1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10486__B1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__B1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10289__B1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10124__B1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__B1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__B1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__B1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__B1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__B1 (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15000__A (.DIODE(_04227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14985__A (.DIODE(_04227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13341__B1 (.DIODE(_04227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__B1 (.DIODE(_04227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__C1 (.DIODE(_04227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__C1 (.DIODE(_04227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09909__A (.DIODE(_04227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__A (.DIODE(_04227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09576__A (.DIODE(_04227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__B1 (.DIODE(_04227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10454__A1 (.DIODE(_04231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__A1 (.DIODE(_04231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__B2 (.DIODE(_04231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10049__A1 (.DIODE(_04231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__A1 (.DIODE(_04231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__A1 (.DIODE(_04231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09929__A1 (.DIODE(_04231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__A (.DIODE(_04231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09685__A1 (.DIODE(_04231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__A1 (.DIODE(_04231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__S0 (.DIODE(_04232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__S0 (.DIODE(_04232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10040__A (.DIODE(_04232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09975__S0 (.DIODE(_04232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09931__S0 (.DIODE(_04232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__S0 (.DIODE(_04232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__S0 (.DIODE(_04232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__S0 (.DIODE(_04232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__S0 (.DIODE(_04232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__S0 (.DIODE(_04232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__S1 (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__S1 (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10041__A (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09975__S1 (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09931__S1 (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__S1 (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__S1 (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__S1 (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__S1 (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__S1 (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__B1 (.DIODE(_04237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__B1 (.DIODE(_04237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__B1 (.DIODE(_04237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10086__B1 (.DIODE(_04237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__C1 (.DIODE(_04237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__B1 (.DIODE(_04237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09642__B1 (.DIODE(_04237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__B1 (.DIODE(_04237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__A (.DIODE(_04237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__B1 (.DIODE(_04237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15675__A1 (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14983__A (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09509__A (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13422__A2 (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__A2 (.DIODE(_04241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__A2 (.DIODE(_04250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__A (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13431__A1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__A1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13351__A1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11196__A (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__A2 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A1 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__A3 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__A0 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A2 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__B1 (.DIODE(_04254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__A3 (.DIODE(_04255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13457__A (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13446__A0 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__A (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__A1 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13373__A2 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11200__A0 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A2 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__A1 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__A1 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__A2 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__B1 (.DIODE(_04265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__A1 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__A1 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A1 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__A1 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__A1 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__A1 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__B2 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__A1 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__A1 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__A1 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15632__A (.DIODE(_04271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10498__A1 (.DIODE(_04271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__A1 (.DIODE(_04271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A1 (.DIODE(_04271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__A1 (.DIODE(_04271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__A1 (.DIODE(_04271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__A1 (.DIODE(_04271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__A1 (.DIODE(_04271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09689__A1 (.DIODE(_04271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__A1 (.DIODE(_04271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13328__A (.DIODE(_04272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__A (.DIODE(_04272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__A1 (.DIODE(_04272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__A (.DIODE(_04272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10125__A1 (.DIODE(_04272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10113__A (.DIODE(_04272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09800__A1 (.DIODE(_04272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09792__A1 (.DIODE(_04272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09575__A1 (.DIODE(_04272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__A1 (.DIODE(_04272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__S0 (.DIODE(_04273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__S0 (.DIODE(_04273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__S0 (.DIODE(_04273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__S0 (.DIODE(_04273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10084__S0 (.DIODE(_04273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__S0 (.DIODE(_04273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__S0 (.DIODE(_04273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__A (.DIODE(_04273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__A (.DIODE(_04273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__A (.DIODE(_04273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__S0 (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__S0 (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__S0 (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__S0 (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__S0 (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09636__S0 (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09635__S0 (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09589__S0 (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__S0 (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__A (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10282__S0 (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10119__S0 (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__S0 (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10115__S0 (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__S0 (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10111__S0 (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__S0 (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09569__S0 (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09568__S0 (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__S0 (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10256__S1 (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__S1 (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__S1 (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__S1 (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__S1 (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09892__S1 (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__S1 (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09638__S1 (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__A (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__A (.DIODE(_04276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__S1 (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__S1 (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__S1 (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__S1 (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__S1 (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09796__S1 (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09704__S1 (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09644__S1 (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__S1 (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__A (.DIODE(_04277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10282__S1 (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10119__S1 (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__S1 (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10115__S1 (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__S1 (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10111__S1 (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__S1 (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09569__S1 (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09568__S1 (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__S1 (.DIODE(_04278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__S0 (.DIODE(_04280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__S0 (.DIODE(_04280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__S0 (.DIODE(_04280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__S0 (.DIODE(_04280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__S0 (.DIODE(_04280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__S0 (.DIODE(_04280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__S0 (.DIODE(_04280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__S0 (.DIODE(_04280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09746__A (.DIODE(_04280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A (.DIODE(_04280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10220__S0 (.DIODE(_04281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10219__S0 (.DIODE(_04281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__S0 (.DIODE(_04281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__S0 (.DIODE(_04281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__S0 (.DIODE(_04281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__S0 (.DIODE(_04281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__S0 (.DIODE(_04281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09922__S0 (.DIODE(_04281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__S0 (.DIODE(_04281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A (.DIODE(_04281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13325__S0 (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__S0 (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__S0 (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__S0 (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10121__S0 (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__S0 (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__S0 (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__S0 (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__S0 (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__S0 (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__S1 (.DIODE(_04283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10390__S1 (.DIODE(_04283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__S1 (.DIODE(_04283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__S1 (.DIODE(_04283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10084__S1 (.DIODE(_04283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__S1 (.DIODE(_04283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__S1 (.DIODE(_04283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09788__A (.DIODE(_04283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09587__A (.DIODE(_04283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__A (.DIODE(_04283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13337__S1 (.DIODE(_04284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13336__S1 (.DIODE(_04284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__S1 (.DIODE(_04284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__S1 (.DIODE(_04284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__S1 (.DIODE(_04284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__S1 (.DIODE(_04284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10077__S1 (.DIODE(_04284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10076__S1 (.DIODE(_04284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__S1 (.DIODE(_04284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__A (.DIODE(_04284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13325__S1 (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__S1 (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__S1 (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__S1 (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10121__S1 (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__S1 (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__S1 (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__S1 (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__S1 (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__S1 (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13327__S (.DIODE(_04287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10285__A1 (.DIODE(_04287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__S (.DIODE(_04287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__S (.DIODE(_04287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__S (.DIODE(_04287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__S (.DIODE(_04287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__S (.DIODE(_04287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__S (.DIODE(_04287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__S (.DIODE(_04287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__S (.DIODE(_04287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10494__A1 (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__A (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10285__C1 (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__A (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__A1 (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__A1 (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__A1 (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__A1 (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__A1 (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__A1 (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10390__S0 (.DIODE(_04290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10256__S0 (.DIODE(_04290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__S0 (.DIODE(_04290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__S0 (.DIODE(_04290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__S0 (.DIODE(_04290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__S0 (.DIODE(_04290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09892__S0 (.DIODE(_04290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__S0 (.DIODE(_04290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09638__S0 (.DIODE(_04290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A (.DIODE(_04290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__S0 (.DIODE(_04291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__S0 (.DIODE(_04291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__S0 (.DIODE(_04291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__S0 (.DIODE(_04291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__S0 (.DIODE(_04291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__S0 (.DIODE(_04291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09706__S0 (.DIODE(_04291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__S0 (.DIODE(_04291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__S0 (.DIODE(_04291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__S0 (.DIODE(_04291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__S1 (.DIODE(_04292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__S1 (.DIODE(_04292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__S1 (.DIODE(_04292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__S1 (.DIODE(_04292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__S1 (.DIODE(_04292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__S1 (.DIODE(_04292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09706__S1 (.DIODE(_04292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__S1 (.DIODE(_04292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__S1 (.DIODE(_04292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__S1 (.DIODE(_04292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13339__B1 (.DIODE(_04296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__C1 (.DIODE(_04296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__B1 (.DIODE(_04296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__A1 (.DIODE(_04296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10147__B1 (.DIODE(_04296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__B1 (.DIODE(_04296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__A1 (.DIODE(_04296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__B1 (.DIODE(_04296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__C1 (.DIODE(_04296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__B1 (.DIODE(_04296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13444__A2 (.DIODE(_04307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__A2 (.DIODE(_04307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__A2 (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__A2 (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__A2 (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__A2 (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__A2 (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__A2 (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__A (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09688__A2 (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__A2 (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09578__A2 (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__S1 (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__S1 (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__S1 (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__S1 (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__S1 (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__S1 (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09636__S1 (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09635__S1 (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09589__S1 (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__S1 (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10428__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10388__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A1 (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09979__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09863__A1 (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09852__A (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__S (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__A (.DIODE(_04320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__S (.DIODE(_04321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__S (.DIODE(_04321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10074__S (.DIODE(_04321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__A1 (.DIODE(_04321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09798__S (.DIODE(_04321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09790__S (.DIODE(_04321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__S (.DIODE(_04321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__S (.DIODE(_04321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09637__S (.DIODE(_04321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__S (.DIODE(_04321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__S0 (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__S0 (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__S0 (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__S0 (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__S0 (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09796__S0 (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09704__S0 (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__S0 (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09644__S0 (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__S0 (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__A1 (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10266__A1 (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10254__C1 (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10086__A1 (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__A1 (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09899__A (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09836__A1 (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09642__A1 (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A1 (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__S0 (.DIODE(_04329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__S0 (.DIODE(_04329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__S0 (.DIODE(_04329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__S0 (.DIODE(_04329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__S0 (.DIODE(_04329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__S0 (.DIODE(_04329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09830__S0 (.DIODE(_04329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__S0 (.DIODE(_04329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__S0 (.DIODE(_04329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__S0 (.DIODE(_04329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15680__A (.DIODE(_04335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14988__A (.DIODE(_04335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13460__B (.DIODE(_04335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__B (.DIODE(_04335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A (.DIODE(_04341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13511__A0 (.DIODE(_04342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13471__A (.DIODE(_04342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13463__A0 (.DIODE(_04342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13433__A1 (.DIODE(_04342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__A2 (.DIODE(_04342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11206__A0 (.DIODE(_04342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__A3 (.DIODE(_04342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A0 (.DIODE(_04342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__A2 (.DIODE(_04342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09616__A2 (.DIODE(_04342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09616__B1 (.DIODE(_04345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13527__A1 (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__A1 (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13478__A0 (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__A (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__A1 (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13403__A2 (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11210__A0 (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A0 (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__A3 (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__A2 (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09692__B (.DIODE(_04363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__B1 (.DIODE(_04363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__S (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__A (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__A (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__S (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09906__S (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09861__A (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09831__S (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09823__S (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__A (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09641__S (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10383__S1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__S1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10252__S1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09897__S1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__S1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09830__S1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__S1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__S1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__S1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__S1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15685__A (.DIODE(_04382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14990__A (.DIODE(_04382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13475__B (.DIODE(_04382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__B (.DIODE(_04382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__C1 (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__B1 (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__B1 (.DIODE(_04390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__A1 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10371__A1 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__A1 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A1 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__A1 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10137__A1 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__A1 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__A1 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__A1 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__A1 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__A2 (.DIODE(_04397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14993__A (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__A (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15690__A1 (.DIODE(_04415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13483__A2 (.DIODE(_04415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09689__A2 (.DIODE(_04415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13535__A1 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13499__A1 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13491__A1 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13409__A (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11216__A0 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__A2 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A2 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A1 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A0 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__A2 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__B2 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__B2 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__B2 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__B2 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__B2 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__B2 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__B2 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__B2 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__B2 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__B1 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__B1 (.DIODE(_04425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__B2 (.DIODE(_04426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__B1 (.DIODE(_04427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09724__A2 (.DIODE(_04429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__S (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10293__A1 (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__A (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__S (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__S (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10120__S (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10051__A (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__A1 (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__S (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15695__A1 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14996__A3 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13502__A2 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__A2 (.DIODE(_04447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14970__B (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10020__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A2 (.DIODE(_04448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13559__A1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13512__A1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13506__A (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13504__A0 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13439__A (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__A (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A3 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09732__A2 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09732__B1 (.DIODE(_04458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__B2 (.DIODE(_04460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13573__A1 (.DIODE(_04466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__A1 (.DIODE(_04466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13523__A1 (.DIODE(_04466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13518__A0 (.DIODE(_04466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13455__A (.DIODE(_04466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__A (.DIODE(_04466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A3 (.DIODE(_04466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A0 (.DIODE(_04466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A2 (.DIODE(_04466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__A2 (.DIODE(_04466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__B1 (.DIODE(_04468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__S1 (.DIODE(_04469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__S1 (.DIODE(_04469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__S1 (.DIODE(_04469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09977__S1 (.DIODE(_04469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__S1 (.DIODE(_04469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__S1 (.DIODE(_04469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__S1 (.DIODE(_04469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09763__S1 (.DIODE(_04469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__S1 (.DIODE(_04469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09744__A (.DIODE(_04469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10220__S1 (.DIODE(_04470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10219__S1 (.DIODE(_04470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__S1 (.DIODE(_04470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__S1 (.DIODE(_04470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__S1 (.DIODE(_04470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__S1 (.DIODE(_04470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__S1 (.DIODE(_04470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09966__S1 (.DIODE(_04470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09922__S1 (.DIODE(_04470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__S1 (.DIODE(_04470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__S0 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__S0 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10216__S0 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__S0 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__S0 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10047__S0 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__S0 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10002__S0 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09923__S0 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__S0 (.DIODE(_04472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__S1 (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__S1 (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10216__S1 (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__S1 (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__S1 (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10047__S1 (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__S1 (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10002__S1 (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09923__S1 (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__S1 (.DIODE(_04473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__S0 (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__S0 (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__S0 (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__S0 (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__S0 (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10010__S0 (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__S0 (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__S0 (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__S0 (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__S0 (.DIODE(_04477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__S1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__S1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__S1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__S1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__S1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10010__S1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__S1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__S1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__S1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__S1 (.DIODE(_04478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10450__A (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__A1 (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__A (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__A1 (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10087__A1 (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10005__A (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09937__A1 (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__A (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__A (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09766__A1 (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__S0 (.DIODE(_04487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__S0 (.DIODE(_04487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__S0 (.DIODE(_04487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09977__S0 (.DIODE(_04487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__S0 (.DIODE(_04487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__S0 (.DIODE(_04487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__S0 (.DIODE(_04487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09856__A (.DIODE(_04487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09763__S0 (.DIODE(_04487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__S0 (.DIODE(_04487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14997__A (.DIODE(_04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13514__A (.DIODE(_04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__B (.DIODE(_04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__C1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__B1 (.DIODE(_04507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__S0 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__S0 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__S0 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__S0 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10073__S0 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__S0 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09855__S0 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__S0 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__S0 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__S0 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__S1 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__S1 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__S1 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__S1 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10073__S1 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__S1 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09855__S1 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__S1 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__S1 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__S1 (.DIODE(_04513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__A2 (.DIODE(_04526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__A2 (.DIODE(_04526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__A3 (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13586__A0 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13533__A1 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13531__A0 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13472__A (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__A0 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__A1 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10669__A0 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A1 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A3 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__B2 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__A2 (.DIODE(_04544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15705__A1 (.DIODE(_04561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15003__A (.DIODE(_04561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09838__A (.DIODE(_04561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13601__A1 (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13557__A1 (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13549__A0 (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13480__A (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__A0 (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__A0 (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10669__A1 (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A2 (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10530__A0 (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__A2 (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__B1 (.DIODE(_04568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09846__B2 (.DIODE(_04569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13338__S (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__S (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__S (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__S (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__S (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__S (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10044__A (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__S (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__S (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09853__S (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13337__S0 (.DIODE(_04579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13336__S0 (.DIODE(_04579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__S0 (.DIODE(_04579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__S0 (.DIODE(_04579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__S0 (.DIODE(_04579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__S0 (.DIODE(_04579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10077__S0 (.DIODE(_04579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10076__S0 (.DIODE(_04579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09966__S0 (.DIODE(_04579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__S0 (.DIODE(_04579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__B (.DIODE(_04581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15005__A (.DIODE(_04592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09870__A (.DIODE(_04592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15709__A1 (.DIODE(_04593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13551__A2 (.DIODE(_04593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A2 (.DIODE(_04593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13616__A1 (.DIODE(_04602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13571__A1 (.DIODE(_04602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13563__A0 (.DIODE(_04602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13500__A (.DIODE(_04602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A (.DIODE(_04602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__A1 (.DIODE(_04602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10669__A2 (.DIODE(_04602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A3 (.DIODE(_04602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10530__A1 (.DIODE(_04602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__A2 (.DIODE(_04602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__B1 (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13629__A0 (.DIODE(_04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13587__A1 (.DIODE(_04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13578__A0 (.DIODE(_04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13557__A0 (.DIODE(_04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13511__A1 (.DIODE(_04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__A (.DIODE(_04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__A3 (.DIODE(_04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10669__A3 (.DIODE(_04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10530__A2 (.DIODE(_04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__A2 (.DIODE(_04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__B1 (.DIODE(_04613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09909__B (.DIODE(_04630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15713__A1 (.DIODE(_04631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15008__A (.DIODE(_04631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13575__B (.DIODE(_04631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__B (.DIODE(_04631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__C1 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13636__A0 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13602__A (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__A0 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13526__A (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__A0 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__A2 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10910__A1 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__A0 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10530__A3 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__A2 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15010__A (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13589__A (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__B (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__B1 (.DIODE(_04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__S (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11160__S (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__S (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__S (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10026__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09990__A (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__B1 (.DIODE(_04668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__B1 (.DIODE(_04673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__B1 (.DIODE(_04673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__B1 (.DIODE(_04673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__A (.DIODE(_04673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__B1 (.DIODE(_04673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__B1 (.DIODE(_04673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__C1 (.DIODE(_04674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15720__A (.DIODE(_04702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15012__A (.DIODE(_04702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13604__A2_N (.DIODE(_04702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09983__B (.DIODE(_04702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09994__B1 (.DIODE(_04707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13649__A1 (.DIODE(_04708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13617__A1 (.DIODE(_04708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13607__A0 (.DIODE(_04708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__A (.DIODE(_04708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__A (.DIODE(_04708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__A3 (.DIODE(_04708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__A1 (.DIODE(_04708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10910__A0 (.DIODE(_04708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__A3 (.DIODE(_04708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__A2 (.DIODE(_04708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__A2 (.DIODE(_04710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__A2 (.DIODE(_04710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__A2 (.DIODE(_04710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11173__A2 (.DIODE(_04710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A2 (.DIODE(_04710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__A2 (.DIODE(_04710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__A2 (.DIODE(_04710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__A2 (.DIODE(_04710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__A2 (.DIODE(_04710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__A2 (.DIODE(_04710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__C1 (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15724__A (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15014__A (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__A (.DIODE(_04737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10029__A3 (.DIODE(_04743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13672__A1 (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13628__A1 (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__A0 (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11267__A (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__A2 (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__A1 (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__A0 (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__A0 (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__A1 (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__A2 (.DIODE(_04744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__S (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__S (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__S (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__S (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__A2 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__A2 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A2 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__A2 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10133__A2 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10027__A2 (.DIODE(_04745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__B2 (.DIODE(_04746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10029__B1 (.DIODE(_04747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10063__A2 (.DIODE(_04753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13686__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13635__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13633__A0 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13572__A (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__A0 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__A3 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__A1 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__A0 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__A0 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__A2 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13334__S0 (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13333__S0 (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__S0 (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__S0 (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10344__S0 (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__S0 (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__S0 (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__S0 (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__S0 (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__S0 (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13334__S1 (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13333__S1 (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__S1 (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__S1 (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10344__S1 (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__S1 (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__S1 (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__S1 (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__S1 (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__S1 (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15016__A (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__A (.DIODE(_04776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15729__A1 (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13622__A2 (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__A2 (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10063__C1 (.DIODE(_04780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__A2 (.DIODE(_04788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15019__A (.DIODE(_04805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__A (.DIODE(_04805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15732__A1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13638__A2 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__A2 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13694__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13647__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13646__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13628__A0 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13586__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__A2 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__A0 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__A2 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__B2 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__B2 (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15736__A1 (.DIODE(_04842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15022__A3 (.DIODE(_04842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13650__A2 (.DIODE(_04842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__A2 (.DIODE(_04842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__A3 (.DIODE(_04847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13673__A (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13664__A1 (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13600__A (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11281__A0 (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A3 (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__A1 (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__A2 (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__A0 (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A0 (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__A2 (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__C1 (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__B1 (.DIODE(_04851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15740__A1 (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15024__A3 (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13675__A2 (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__A2 (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13707__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13677__A0 (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13665__A (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A2 (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__A1 (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10994__B (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__A0 (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__A0 (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A1 (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__A2 (.DIODE(_04880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__B2 (.DIODE(_04881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__A2 (.DIODE(_04890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15025__A (.DIODE(_04908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__A (.DIODE(_04908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15744__A1 (.DIODE(_04909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13689__A2 (.DIODE(_04909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__A2 (.DIODE(_04909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13744__A1 (.DIODE(_04913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13701__A1 (.DIODE(_04913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13693__A1 (.DIODE(_04913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13691__A0 (.DIODE(_04913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13674__A1 (.DIODE(_04913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13629__A1 (.DIODE(_04913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__A0 (.DIODE(_04913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11014__A2 (.DIODE(_04913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A1 (.DIODE(_04913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__A2 (.DIODE(_04913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__B2 (.DIODE(_04914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__B2 (.DIODE(_04915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A2 (.DIODE(_04923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15027__A (.DIODE(_04940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__A (.DIODE(_04940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15748__A1 (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13696__A2 (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A2 (.DIODE(_04941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13754__A1 (.DIODE(_04945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13718__A1 (.DIODE(_04945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13704__A1 (.DIODE(_04945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13688__A1 (.DIODE(_04945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13636__A1 (.DIODE(_04945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__A2 (.DIODE(_04945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11022__A1 (.DIODE(_04945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A0 (.DIODE(_04945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__A1 (.DIODE(_04945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__A2 (.DIODE(_04945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__B2 (.DIODE(_04946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__B2 (.DIODE(_04947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13776__A1 (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13732__A1 (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13723__A0 (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13648__A (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__A1 (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__A3 (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__A1 (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11022__A0 (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__A0 (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__A2 (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__B2 (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__A2 (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15751__A1 (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15030__A3 (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__A2 (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__A2 (.DIODE(_04979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__C1 (.DIODE(_04982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15755__A1 (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15032__A3 (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13733__A2 (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__A2 (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13742__A (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13735__A0 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13726__A (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__A0 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__A2 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11051__A1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__A0 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10609__A0 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__A1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__A2 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__B2 (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15758__A (.DIODE(_05037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15033__A (.DIODE(_05037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13746__A (.DIODE(_05037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__B (.DIODE(_05037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13802__A1 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13752__A1 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13750__A0 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13685__A (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11315__A1 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__A3 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__A1 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11051__A0 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__A0 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__A2 (.DIODE(_05044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__B2 (.DIODE(_05045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__B2 (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15762__A (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15035__A (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13755__A (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__B (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14892__B2 (.DIODE(_05076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13774__A1 (.DIODE(_05076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13762__A1 (.DIODE(_05076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13694__A0 (.DIODE(_05076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11320__A0 (.DIODE(_05076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__A2 (.DIODE(_05076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__A1 (.DIODE(_05076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__A0 (.DIODE(_05076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__A1 (.DIODE(_05076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__A2 (.DIODE(_05076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__B2 (.DIODE(_05077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__B2 (.DIODE(_05078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13789__A1 (.DIODE(_05086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13786__A (.DIODE(_05086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13780__A0 (.DIODE(_05086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13717__A (.DIODE(_05086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11326__A0 (.DIODE(_05086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__A3 (.DIODE(_05086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__A1 (.DIODE(_05086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11096__A2 (.DIODE(_05086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__A0 (.DIODE(_05086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__A2 (.DIODE(_05086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__B2 (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15037__A (.DIODE(_05106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10399__A (.DIODE(_05106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15768__A1 (.DIODE(_05107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__A2 (.DIODE(_05107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10401__A2 (.DIODE(_05107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__C1 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15039__A (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__A (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15772__A1 (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13792__A2 (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__A2 (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13801__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13794__A0 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13774__A0 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13731__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__A0 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__A2 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__A1 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__B (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__A0 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__A2 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__B2 (.DIODE(_05144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__A3 (.DIODE(_05145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15041__A (.DIODE(_05169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10464__A (.DIODE(_05169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15775__A1 (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13803__A2 (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__A2 (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14892__A1 (.DIODE(_05174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13805__A0 (.DIODE(_05174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13797__A (.DIODE(_05174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13796__A (.DIODE(_05174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13789__A0 (.DIODE(_05174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13744__A0 (.DIODE(_05174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__A1 (.DIODE(_05174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__A1 (.DIODE(_05174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__A0 (.DIODE(_05174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__A2 (.DIODE(_05174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__B2 (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10471__B2 (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15043__A (.DIODE(_05200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14893__B1 (.DIODE(_05200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__A (.DIODE(_05200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14896__A1 (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14888__A (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13753__A (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__A0 (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__A0 (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10632__B1 (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__B_N (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10613__B1 (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__A1 (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__A2 (.DIODE(_05205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__B2 (.DIODE(_05206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10503__B2 (.DIODE(_05207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13455__B (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13413__A (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10523__A (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__A (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13355__B1 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__A (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11103__B1 (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__A2 (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__B1 (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10917__A2 (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__A (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__C (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11103__A2 (.DIODE(_05215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11025__B1 (.DIODE(_05215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__B1 (.DIODE(_05215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11004__B1 (.DIODE(_05215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__A2 (.DIODE(_05215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10937__B1 (.DIODE(_05215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__B1 (.DIODE(_05215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__B1 (.DIODE(_05215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__A (.DIODE(_05215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__D (.DIODE(_05215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11080__A (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__B1 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10999__B1 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__B1 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10802__A (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10735__B1 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__A (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10515__A (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__A1 (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11108__A1 (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__A1 (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11032__A (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__A (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__A1 (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10876__A1 (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__A1 (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__A1 (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__A2 (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__B1 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__A1_N (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__B (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__B1 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10599__B1 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__A2 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__A2 (.DIODE(_05221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11072__B1 (.DIODE(_05221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__B1 (.DIODE(_05221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11025__A2_N (.DIODE(_05221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__B1 (.DIODE(_05221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__A2_N (.DIODE(_05221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10705__A2 (.DIODE(_05221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A (.DIODE(_05221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10519__A2_N (.DIODE(_05221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11119__A2 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__B1 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__A2 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10937__A2 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10766__A2 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A3 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__A2 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__A2 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__A3 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10519__B1 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11064__A (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__A1 (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__A1 (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10787__A1 (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10660__A (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__A1 (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10625__B2 (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10549__B (.DIODE(_05225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13789__S (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13775__A1 (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13774__S (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13753__B (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13717__B (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13600__B (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13557__S (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__A2 (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10866__B (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10524__B (.DIODE(_05227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11051__S (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11022__S (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__S (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10910__S (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10669__S0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10621__A (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__B (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__S0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10530__S0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__S0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__S1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__S1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10817__S (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__S0 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__S0 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__S (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__S1 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10562__A (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__C (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__S0 (.DIODE(_05235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__S (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__S0 (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__S0 (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__S0 (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__S1 (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__S1 (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__S1 (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10641__A2 (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__S1 (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__S1 (.DIODE(_05237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__S (.DIODE(_05239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__S (.DIODE(_05239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__S (.DIODE(_05239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__S1 (.DIODE(_05239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__S0 (.DIODE(_05239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__S0 (.DIODE(_05239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__S0 (.DIODE(_05239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__S1 (.DIODE(_05239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__S1 (.DIODE(_05239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__A (.DIODE(_05239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__A1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10912__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__S (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10790__S (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__S1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__A (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10541__S1 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__S (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10835__S (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__S (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10739__A1 (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10704__S (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10695__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10650__S (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__S (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__S (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__A (.DIODE(_05246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__C1 (.DIODE(_05251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__B1 (.DIODE(_05251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__C1 (.DIODE(_05251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__C1 (.DIODE(_05251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10976__B2 (.DIODE(_05251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__B2 (.DIODE(_05251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10766__B1 (.DIODE(_05251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__B2 (.DIODE(_05251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10578__A (.DIODE(_05251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__B2 (.DIODE(_05251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__A2 (.DIODE(_05254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A0 (.DIODE(_05254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__A2 (.DIODE(_05254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11119__B2 (.DIODE(_05254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__B1_N (.DIODE(_05254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__B2 (.DIODE(_05254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__B2 (.DIODE(_05254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__A (.DIODE(_05254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10685__A (.DIODE(_05254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__A (.DIODE(_05254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16129__A1 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15112__A1 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10992__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10971__A1 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__A1 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__A1 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__A1 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__A1 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10625__A1 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__A1 (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13671__B (.DIODE(_05257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13457__B (.DIODE(_05257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13454__A (.DIODE(_05257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__S (.DIODE(_05257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13387__S (.DIODE(_05257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13368__S (.DIODE(_05257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__A (.DIODE(_05257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13601__A2 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13587__A2 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13512__A2 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13471__B (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__A2 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__B (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13403__A3 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__A3 (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10736__B (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__A (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13802__A2 (.DIODE(_05260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13752__A2 (.DIODE(_05260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13647__A2 (.DIODE(_05260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13617__A2 (.DIODE(_05260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13499__A2 (.DIODE(_05260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__A2 (.DIODE(_05260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13412__A2 (.DIODE(_05260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13351__C1 (.DIODE(_05260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10685__B (.DIODE(_05260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__A (.DIODE(_05260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13754__A2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13693__A2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13649__A2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13635__A2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__A2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__B (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__A2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__A2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10625__A2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__A2 (.DIODE(_05261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__S0 (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__S0 (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__S0 (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__S (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__S0 (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__S (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__S0 (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__S0 (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__S (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__S (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__A2 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__A0 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__S1 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__A1 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A1 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__S (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10749__S0 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__A1 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10694__S0 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__S0 (.DIODE(_05277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11120__B2 (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__A1 (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__B2 (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11006__A1 (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10989__A1 (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__B2 (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__A1 (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A1 (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__A1 (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__A1 (.DIODE(_05281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16123__A1 (.DIODE(_05286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15099__A1 (.DIODE(_05286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A2 (.DIODE(_05286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__A0 (.DIODE(_05286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__A2 (.DIODE(_05286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__S1 (.DIODE(_05286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__S0 (.DIODE(_05286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__S1 (.DIODE(_05286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__S0 (.DIODE(_05286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__A2 (.DIODE(_05286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__A (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__A1 (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10872__A (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10836__S (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__S (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__A1 (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__S1 (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10696__S1 (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10651__S (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__A (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15109__A1 (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11024__A (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__A1 (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10884__S (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10867__A (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__A1 (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10813__A1 (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__S (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10749__S1 (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__A1 (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__A2 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A0 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10915__A (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10898__A (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10853__A (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__A (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10820__A (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10715__A (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__S (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__A (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11128__B (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11004__A2 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__A2 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__A2 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__A2_N (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__B1 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__B (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__A2 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__B1 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10599__A2 (.DIODE(_05301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__S (.DIODE(_05322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__B1 (.DIODE(_05322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10620__A (.DIODE(_05322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__A1 (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11077__A (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__A1 (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10996__S (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__C1 (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10800__A1 (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__A (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__A (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__S (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__A (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16121__A1 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15076__A1 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__A2 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__A0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__A2 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__S0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__S (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__S0 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__S1 (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__B (.DIODE(_05324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13775__A2 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__B1 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__B (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__B1 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10917__B1 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__B (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10694__A3 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10633__A1 (.DIODE(_05334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__B1 (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__B1 (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10747__B1 (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10705__B1 (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10655__A (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11129__B1 (.DIODE(_05357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__A2 (.DIODE(_05357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__A2 (.DIODE(_05357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10963__A2 (.DIODE(_05357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10887__A2 (.DIODE(_05357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10865__B1 (.DIODE(_05357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__A2 (.DIODE(_05357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__B1 (.DIODE(_05357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__B1 (.DIODE(_05357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__B (.DIODE(_05357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__A1 (.DIODE(_05361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__A1 (.DIODE(_05361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10954__A1 (.DIODE(_05361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A1 (.DIODE(_05361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10907__A1 (.DIODE(_05361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__A1 (.DIODE(_05361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__A1 (.DIODE(_05361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__A1 (.DIODE(_05361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10709__A1 (.DIODE(_05361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__A1 (.DIODE(_05361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__A1 (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11085__S (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__A1 (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__S (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10878__S (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__S (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10810__S (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__S (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10733__S (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10663__S (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__B1 (.DIODE(_05367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__A2_N (.DIODE(_05367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10973__A2 (.DIODE(_05367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10886__B1 (.DIODE(_05367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10864__B (.DIODE(_05367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__B1 (.DIODE(_05367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__B1 (.DIODE(_05367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__A2 (.DIODE(_05367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10747__A2 (.DIODE(_05367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__B (.DIODE(_05367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11096__B1 (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10921__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10894__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10826__C1 (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__S (.DIODE(_05390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10971__A2 (.DIODE(_05394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__A3 (.DIODE(_05394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11072__A2 (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__A2 (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__A2_N (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__A (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11104__A2 (.DIODE(_05398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__A2 (.DIODE(_05398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__B (.DIODE(_05398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10986__A2 (.DIODE(_05398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__A2 (.DIODE(_05398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10916__B (.DIODE(_05398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10886__A2 (.DIODE(_05398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__A2 (.DIODE(_05398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__A (.DIODE(_05398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__A2 (.DIODE(_05398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11087__A2 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10976__A1_N (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10854__A2 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__B2 (.DIODE(_05404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16125__A1 (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15105__A1 (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__A2 (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__A1 (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11102__S (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__S1 (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__S (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__S0 (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__S0 (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__S0 (.DIODE(_05413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16127__A1 (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__A2 (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11087__A1 (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__A1 (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10890__A (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10863__A (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10854__A1 (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__S1 (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__S1 (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__S1 (.DIODE(_05414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__A1 (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__A (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11129__A2 (.DIODE(_05440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__A2 (.DIODE(_05440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__B2 (.DIODE(_05440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__A2 (.DIODE(_05440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10865__A2 (.DIODE(_05440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10833__A2 (.DIODE(_05440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__A2 (.DIODE(_05440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__A2_N (.DIODE(_05440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__A2 (.DIODE(_05440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10748__A2 (.DIODE(_05440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__A1 (.DIODE(_05458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__A3 (.DIODE(_05458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__A1 (.DIODE(_05461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__A0 (.DIODE(_05461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10766__B2 (.DIODE(_05461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__A (.DIODE(_05498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15921__B2 (.DIODE(_05517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11126__A1 (.DIODE(_05517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__A (.DIODE(_05517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11112__B1 (.DIODE(_05517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11097__B1 (.DIODE(_05517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10982__A1 (.DIODE(_05517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__S (.DIODE(_05517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__A1 (.DIODE(_05517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__B1 (.DIODE(_05517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__A1 (.DIODE(_05517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10977__A1 (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10853__B (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__B1 (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16113__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__A2 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__A2 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__A2 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__A2 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__B1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__A3 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__C (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11199__B (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__A2 (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11213__B (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__B (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__B1 (.DIODE(_05851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11213__C (.DIODE(_05851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__B (.DIODE(_05860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__B (.DIODE(_05860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__A2 (.DIODE(_05864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__B (.DIODE(_05864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11229__B (.DIODE(_05864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__B (.DIODE(_05864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__A3 (.DIODE(_05868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__C (.DIODE(_05868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__B (.DIODE(_05868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__B1 (.DIODE(_05871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__D (.DIODE(_05871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__A2 (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__B (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__B (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__B (.DIODE(_05881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__B1 (.DIODE(_05881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__B (.DIODE(_05881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__C (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11257__B (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11254__B (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__D (.DIODE(_05889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__B (.DIODE(_05889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__B (.DIODE(_05894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__B (.DIODE(_05894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__B (.DIODE(_05899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11275__A2 (.DIODE(_05899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__B (.DIODE(_05899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__C (.DIODE(_05902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11275__B1 (.DIODE(_05902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__B (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__A2 (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__B (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__C (.DIODE(_05911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__B1 (.DIODE(_05911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__B (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__A2 (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__B (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__C (.DIODE(_05918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__B1 (.DIODE(_05918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11302__B (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11301__B (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11318__B (.DIODE(_05929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__B (.DIODE(_05929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__A2 (.DIODE(_05929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__B (.DIODE(_05929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11318__C (.DIODE(_05932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__C (.DIODE(_05932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__B1 (.DIODE(_05932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11319__A2 (.DIODE(_05937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11318__D (.DIODE(_05937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11328__B (.DIODE(_05943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11325__B (.DIODE(_05943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11337__B (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11336__A2 (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11331__B (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11337__C (.DIODE(_05952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11336__B1 (.DIODE(_05952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__B (.DIODE(_05957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15969__B1 (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11418__A (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__A1_N (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__C (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11394__B (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16082__B1 (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16002__A2 (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15992__A1 (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15989__B1 (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15842__B1 (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15819__A2 (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15817__A2 (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15816__A2 (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15804__B2 (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__A2 (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16095__C1 (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15794__C1 (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15789__C1 (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15788__C1 (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15725__C1 (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15698__C1 (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15690__C1 (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15686__C1 (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15668__C1 (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__A1 (.DIODE(_06026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14755__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14158__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14097__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13988__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13924__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13891__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13871__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__A3 (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__A (.DIODE(_06053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13985__B1 (.DIODE(_06054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__A1 (.DIODE(_06054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__A1 (.DIODE(_06054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__A1 (.DIODE(_06054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__A1 (.DIODE(_06054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__A1 (.DIODE(_06054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__A1 (.DIODE(_06054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__A1 (.DIODE(_06054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__A1 (.DIODE(_06054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__A1 (.DIODE(_06054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11699__A (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11618__B1 (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__B1 (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11526__A (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__B (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__B (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__A (.DIODE(_06065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11691__B1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__B1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11673__B1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__B1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__B1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__B1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__B1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11629__B1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11522__A1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11503__A1 (.DIODE(_06066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15789__B2 (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11797__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11753__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13872__A (.DIODE(_06072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__A1 (.DIODE(_06072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__A1 (.DIODE(_06072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__A1 (.DIODE(_06072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__A1 (.DIODE(_06072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__A1 (.DIODE(_06072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__B2 (.DIODE(_06072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11530__B2 (.DIODE(_06072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11516__B2 (.DIODE(_06072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__B2 (.DIODE(_06072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16609__A1 (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__A (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__A (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11504__A (.DIODE(_06077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12816__A0 (.DIODE(_06078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__A0 (.DIODE(_06078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12599__A0 (.DIODE(_06078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12462__A0 (.DIODE(_06078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__A0 (.DIODE(_06078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__A0 (.DIODE(_06078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__A0 (.DIODE(_06078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11878__A0 (.DIODE(_06078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11807__A0 (.DIODE(_06078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__A0 (.DIODE(_06078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16471__D (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16334__D (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16209__A1 (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__A_N (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__B_N (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__A_N (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__A (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__B (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__C (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11510__B_N (.DIODE(_06081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16471__B_N (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16334__B_N (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16208__A1 (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__B_N (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__C (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__B (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__B (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__C (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__A_N (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11510__C (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16334__C (.DIODE(_06083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__C (.DIODE(_06083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__D_N (.DIODE(_06083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__A (.DIODE(_06083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__D (.DIODE(_06083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11874__B (.DIODE(_06083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11510__D (.DIODE(_06083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__S (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11592__S (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__S (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11574__S (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__S (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__S (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__S (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11534__S (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11524__S (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__S (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11751__B1 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__B1 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__B1 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__B1 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11643__B1 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__B2 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11532__B2 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11521__B1 (.DIODE(_06093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16611__A1 (.DIODE(_06095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12887__A (.DIODE(_06095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__A (.DIODE(_06095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__A (.DIODE(_06095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__B1 (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__B1 (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11605__B1 (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11595__B1 (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__B1 (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__B1 (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11560__B1 (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__B1 (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__A (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11528__A (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11795__B1 (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11787__B1 (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11778__B1 (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__B1 (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11743__B1 (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__B1 (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__B1 (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11661__B1 (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__C1 (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11530__C1 (.DIODE(_06101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16613__A1 (.DIODE(_06104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12890__A (.DIODE(_06104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12158__A (.DIODE(_06104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__A (.DIODE(_06104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__A0 (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__A0 (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__A0 (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12466__A0 (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12087__A0 (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12019__A0 (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__A0 (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__A0 (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__A0 (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11534__A0 (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16615__A1 (.DIODE(_06113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__A (.DIODE(_06113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__A (.DIODE(_06113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A (.DIODE(_06113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__A0 (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__A0 (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12605__A0 (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12468__A0 (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__A0 (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__A0 (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__A0 (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__A0 (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__A0 (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__A0 (.DIODE(_06114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11799__A1 (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__A1 (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__A1 (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__A1 (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__A1 (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11606__A1 (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__A1 (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__A1 (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__A1 (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__A1 (.DIODE(_06116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11761__B (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__B (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11709__B (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__B (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__B (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11627__B (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11595__C1 (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__C1 (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__C1 (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__C1 (.DIODE(_06118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16617__A1 (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__A (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12164__A (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__A (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16619__A1 (.DIODE(_06131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__A (.DIODE(_06131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__A (.DIODE(_06131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__A (.DIODE(_06131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__A0 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12678__A0 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__A0 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__A0 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__A0 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__A0 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__A0 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__A0 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11817__A0 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__A0 (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16621__A1 (.DIODE(_06140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__A (.DIODE(_06140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12170__A (.DIODE(_06140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11573__A (.DIODE(_06140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16623__A1 (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12905__A (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12173__A (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11583__A (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__A0 (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12682__A0 (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12613__A0 (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12476__A0 (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12097__A0 (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__A0 (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11961__A0 (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__A0 (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__A0 (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__A0 (.DIODE(_06150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16625__A1 (.DIODE(_06156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__A (.DIODE(_06156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12176__A (.DIODE(_06156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11591__A (.DIODE(_06156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16627__A1 (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__A (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__A (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__A (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__A0 (.DIODE(_06166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12686__A0 (.DIODE(_06166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12617__A0 (.DIODE(_06166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12480__A0 (.DIODE(_06166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12101__A0 (.DIODE(_06166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12033__A0 (.DIODE(_06166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11965__A0 (.DIODE(_06166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__A0 (.DIODE(_06166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11825__A0 (.DIODE(_06166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__A0 (.DIODE(_06166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16630__A1 (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12914__A (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12182__A (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__A (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11685__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11649__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11632__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11622__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11613__S (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16632__A1 (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12918__A (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__A (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__A (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__A0 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__A0 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12622__A0 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__A0 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12106__A0 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12038__A0 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11970__A0 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11901__A0 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11830__A0 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11622__A0 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15780__A1 (.DIODE(_06186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15779__B2 (.DIODE(_06186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14966__A (.DIODE(_06186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__A0 (.DIODE(_06186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__A (.DIODE(_06186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__A1 (.DIODE(_06186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A1 (.DIODE(_06186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__A1 (.DIODE(_06186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A1 (.DIODE(_06186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11630__A1 (.DIODE(_06186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16634__A1 (.DIODE(_06192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12921__A (.DIODE(_06192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__A (.DIODE(_06192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__A (.DIODE(_06192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12841__A0 (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__A0 (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12624__A0 (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12487__A0 (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__A0 (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12040__A0 (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11972__A0 (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11903__A0 (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11832__A0 (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11632__A0 (.DIODE(_06193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16636__A1 (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__A (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12192__A (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11640__A (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16638__A1 (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12927__A (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__A (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__A (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16640__A1 (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12930__A (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12198__A (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__A (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12847__A0 (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__A0 (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12630__A0 (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__A0 (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__A0 (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12046__A0 (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__A0 (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__A0 (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__A0 (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__A0 (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16642__A1 (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12933__A (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__A (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11666__A (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16644__A1 (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12936__A (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12204__A (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11675__A (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16646__A1 (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12939__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__A0 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__A0 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__A0 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__A0 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__A0 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__A0 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11984__A0 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__A0 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__A0 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11685__A0 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16648__A1 (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12942__A (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12210__A (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__A (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11781__A1 (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__A1 (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11763__A1 (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__A1 (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__A1 (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11737__A1 (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A1 (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A1 (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__A1 (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11701__A1 (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16651__A1 (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12945__A (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__A (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11703__A (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__A0 (.DIODE(_06257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__A0 (.DIODE(_06257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__A0 (.DIODE(_06257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__A0 (.DIODE(_06257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__A0 (.DIODE(_06257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12057__A0 (.DIODE(_06257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__A0 (.DIODE(_06257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11920__A0 (.DIODE(_06257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11849__A0 (.DIODE(_06257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__A0 (.DIODE(_06257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11784__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11775__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11731__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11723__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11714__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__S (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16653__A1 (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12949__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12217__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11713__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__A0 (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__A0 (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__A0 (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__A0 (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12127__A0 (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12059__A0 (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__A0 (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11922__A0 (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__A0 (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11714__A0 (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16655__A1 (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12952__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16657__A1 (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12955__A (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__A (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__A (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16659__A1 (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__A (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__A (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__A (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16661__A1 (.DIODE(_06296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12961__A (.DIODE(_06296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__A (.DIODE(_06296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__A (.DIODE(_06296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16663__A1 (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12964__A (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12232__A (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__A (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16665__A1 (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__A (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__A (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__A (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12872__A0 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__A0 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12655__A0 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12518__A0 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12139__A0 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__A0 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12003__A0 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__A0 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__A0 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__A0 (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16667__A1 (.DIODE(_06319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__A (.DIODE(_06319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12238__A (.DIODE(_06319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11774__A (.DIODE(_06319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12874__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12657__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12520__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11936__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11775__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16669__A1 (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11783__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12659__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12522__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12007__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11938__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11784__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16671__A1 (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__A (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__A (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11792__A (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12524__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12145__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12077__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12009__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16673__A1 (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12979__A (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__A (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__A (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11825__S (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__S (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__S (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__S (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11817__S (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11815__S (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__S (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__S (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11809__S (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11807__S (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11846__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11832__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11830__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__S (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__S (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__S (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__S (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__S (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11857__S (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__S (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11853__S (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__S (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11849__S (.DIODE(_06370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__S (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__S (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__S (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__S (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__S (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__S (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__S (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__S (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__S (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11878__S (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__S (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__S (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__S (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__S (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__S (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11907__S (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11905__S (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11903__S (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11901__S (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11899__S (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11938__S (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11936__S (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__S (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__S (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__S (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11928__S (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11926__S (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__S (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11922__S (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11920__S (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11965__S (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11963__S (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11961__S (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__S (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__S (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__S (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__S (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__S (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__S (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__S (.DIODE(_06424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11986__S (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11984__S (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11982__S (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11980__S (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__S (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__S (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11974__S (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11972__S (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11970__S (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11968__S (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12007__S (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__S (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12003__S (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12001__S (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11999__S (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__S (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__S (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__S (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__S (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__S (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12033__S (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12031__S (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__S (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12027__S (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__S (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12023__S (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__S (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12019__S (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12017__S (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__S (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__S (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__S (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__S (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__S (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12046__S (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12044__S (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12042__S (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12040__S (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12038__S (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12036__S (.DIODE(_06471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__S (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__S (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__S (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__S (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__S (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__S (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12063__S (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__S (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12059__S (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12057__S (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12101__S (.DIODE(_06496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__S (.DIODE(_06496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12097__S (.DIODE(_06496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__S (.DIODE(_06496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__S (.DIODE(_06496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12091__S (.DIODE(_06496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__S (.DIODE(_06496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12087__S (.DIODE(_06496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12085__S (.DIODE(_06496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__S (.DIODE(_06496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12122__S (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__S (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__S (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__S (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__S (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12112__S (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12110__S (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__S (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12106__S (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__S (.DIODE(_06507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__S (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__S (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12139__S (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__S (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__S (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__S (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__S (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__S (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12127__S (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__S (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__S (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__S (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__A (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12183__A (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12152__A (.DIODE(_06533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12180__S (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__S (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12174__S (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__S (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12168__S (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__S (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12162__S (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__S (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__S (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12153__S (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16821__A0 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16753__A0 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16475__A1 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__A1 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__A1 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__A1 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__A1 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__A1 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12257__A1 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__A1 (.DIODE(_06536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16825__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16757__A0 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16479__A1 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__A1 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__A1 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__A1 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__A1 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12330__A1 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__A1 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12162__A1 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16840__A0 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16772__A0 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16494__A1 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13005__A1 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__A1 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__A1 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12414__A1 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12345__A1 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__A1 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12184__A1 (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__S (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12208__S (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__S (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12202__S (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__S (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__S (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12193__S (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__S (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12187__S (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12184__S (.DIODE(_06555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16850__A0 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16782__A0 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16504__A1 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__A1 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__A1 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__A1 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__A1 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__A1 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__A1 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__A1 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16854__A0 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16786__A0 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16508__A1 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__A1 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__A1 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__A1 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__A1 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__A1 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12290__A1 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__A1 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16856__A0 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16788__A0 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16510__A1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13021__A1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__A1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__A1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12430__A1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__A1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__A1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12208__A1 (.DIODE(_06571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16861__A0 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16793__A0 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16515__A1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__A1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__A1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__A1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12435__A1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12366__A1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12297__A1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__A1 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__S (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12239__S (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__S (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12233__S (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__S (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12227__S (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__S (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__S (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__S (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__S (.DIODE(_06576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16863__A0 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16795__A0 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16517__A1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__A1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12791__A1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12575__A1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__A1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12368__A1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__A1 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16865__A0 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16797__A0 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16519__A1 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__A1 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__A1 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__A1 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__A1 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__A1 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__A1 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__A1 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16867__A0 (.DIODE(_06582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16799__A0 (.DIODE(_06582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16521__A1 (.DIODE(_06582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__A1 (.DIODE(_06582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12795__A1 (.DIODE(_06582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__A1 (.DIODE(_06582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__A1 (.DIODE(_06582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__A1 (.DIODE(_06582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__A1 (.DIODE(_06582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__A1 (.DIODE(_06582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16869__A0 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16801__A0 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16523__A1 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__A1 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__A1 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__A1 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__A1 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__A1 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12305__A1 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12227__A1 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16871__A0 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16803__A0 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16525__A1 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__A1 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__A1 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__A1 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__A1 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__A1 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__A1 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__A1 (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16873__A0 (.DIODE(_06588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16805__A0 (.DIODE(_06588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16527__A1 (.DIODE(_06588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__A1 (.DIODE(_06588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__A1 (.DIODE(_06588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__A1 (.DIODE(_06588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__A1 (.DIODE(_06588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__A1 (.DIODE(_06588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__A1 (.DIODE(_06588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12233__A1 (.DIODE(_06588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16875__A0 (.DIODE(_06590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16807__A0 (.DIODE(_06590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16529__A1 (.DIODE(_06590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13040__A1 (.DIODE(_06590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12803__A1 (.DIODE(_06590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__A1 (.DIODE(_06590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__A1 (.DIODE(_06590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__A1 (.DIODE(_06590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__A1 (.DIODE(_06590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__A1 (.DIODE(_06590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16883__A0 (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16815__A0 (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16537__A1 (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__A1 (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12811__A1 (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__A1 (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__A1 (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__A1 (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__A1 (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__A1 (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__S (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__S (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__A (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__A (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__A (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__S (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12271__S (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__S (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__S (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__S (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__S (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__S (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12259__S (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12257__S (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__S (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12294__S (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__S (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12290__S (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12288__S (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__S (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12284__S (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12282__S (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__S (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__S (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__S (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__S (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__S (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__S (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__S (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__S (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12305__S (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__S (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__S (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__S (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12297__S (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__S (.DIODE(_06640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__S (.DIODE(_06640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__A (.DIODE(_06640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__A (.DIODE(_06640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__A (.DIODE(_06640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__S (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__S (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12338__S (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__S (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12334__S (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12332__S (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12330__S (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__S (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__S (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12324__S (.DIODE(_06641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__S (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__S (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__S (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__S (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__S (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__S (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__S (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__S (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__S (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12345__S (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__S (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__S (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__S (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__S (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__S (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__S (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__S (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__S (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12368__S (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12366__S (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__S (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__S (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12434__A (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12413__A (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__A (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12411__S (.DIODE(_06678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12409__S (.DIODE(_06678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12407__S (.DIODE(_06678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12405__S (.DIODE(_06678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__S (.DIODE(_06678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12401__S (.DIODE(_06678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__S (.DIODE(_06678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__S (.DIODE(_06678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__S (.DIODE(_06678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12393__S (.DIODE(_06678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12432__S (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12430__S (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__S (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__S (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__S (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__S (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__S (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__S (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__S (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12414__S (.DIODE(_06689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__S (.DIODE(_06700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__S (.DIODE(_06700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__S (.DIODE(_06700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__S (.DIODE(_06700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__S (.DIODE(_06700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__S (.DIODE(_06700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__S (.DIODE(_06700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__S (.DIODE(_06700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__S (.DIODE(_06700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12435__S (.DIODE(_06700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12480__S (.DIODE(_06715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__S (.DIODE(_06715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12476__S (.DIODE(_06715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12474__S (.DIODE(_06715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__S (.DIODE(_06715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__S (.DIODE(_06715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12468__S (.DIODE(_06715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12466__S (.DIODE(_06715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12464__S (.DIODE(_06715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12462__S (.DIODE(_06715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__S (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__S (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12497__S (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__S (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__S (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12491__S (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12489__S (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12487__S (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__S (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__S (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12522__S (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12520__S (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12518__S (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12516__S (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12514__S (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__S (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12510__S (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12508__S (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__S (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__S (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__S (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12593__S (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__A (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__A (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12530__A (.DIODE(_06751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12549__S (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__S (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__S (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12543__S (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__S (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12539__S (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__S (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__S (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__S (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__S (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12570__S (.DIODE(_06763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__S (.DIODE(_06763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__S (.DIODE(_06763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__S (.DIODE(_06763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__S (.DIODE(_06763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__S (.DIODE(_06763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12558__S (.DIODE(_06763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__S (.DIODE(_06763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12554__S (.DIODE(_06763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__S (.DIODE(_06763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12591__S (.DIODE(_06774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12589__S (.DIODE(_06774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__S (.DIODE(_06774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__S (.DIODE(_06774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__S (.DIODE(_06774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__S (.DIODE(_06774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__S (.DIODE(_06774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__S (.DIODE(_06774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12575__S (.DIODE(_06774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__S (.DIODE(_06774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12617__S (.DIODE(_06788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__S (.DIODE(_06788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12613__S (.DIODE(_06788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__S (.DIODE(_06788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__S (.DIODE(_06788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__S (.DIODE(_06788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12605__S (.DIODE(_06788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__S (.DIODE(_06788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12601__S (.DIODE(_06788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12599__S (.DIODE(_06788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__S (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__S (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12634__S (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12632__S (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12630__S (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12628__S (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__S (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12624__S (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12622__S (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__S (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12659__S (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12657__S (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12655__S (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12653__S (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12651__S (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__S (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__S (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__S (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__S (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__S (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12686__S (.DIODE(_06825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12684__S (.DIODE(_06825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12682__S (.DIODE(_06825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12680__S (.DIODE(_06825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12678__S (.DIODE(_06825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12676__S (.DIODE(_06825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__S (.DIODE(_06825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__S (.DIODE(_06825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__S (.DIODE(_06825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__S (.DIODE(_06825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__S (.DIODE(_06836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__S (.DIODE(_06836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12703__S (.DIODE(_06836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__S (.DIODE(_06836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__S (.DIODE(_06836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__S (.DIODE(_06836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12695__S (.DIODE(_06836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__S (.DIODE(_06836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__S (.DIODE(_06836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__S (.DIODE(_06836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__S (.DIODE(_06847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__S (.DIODE(_06847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__S (.DIODE(_06847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__S (.DIODE(_06847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__S (.DIODE(_06847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__S (.DIODE(_06847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12716__S (.DIODE(_06847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__S (.DIODE(_06847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__S (.DIODE(_06847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__S (.DIODE(_06847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14455__A (.DIODE(_06860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14319__A (.DIODE(_06860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14313__C1 (.DIODE(_06860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14202__A (.DIODE(_06860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12735__B (.DIODE(_06860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__B2 (.DIODE(_06861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__B2 (.DIODE(_06861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__B2 (.DIODE(_06861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__B1 (.DIODE(_06861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16209__A2 (.DIODE(_06862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16208__A2 (.DIODE(_06862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__A2 (.DIODE(_06862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__A2 (.DIODE(_06862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__A2 (.DIODE(_06862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16207__C (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15792__B (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14482__B2 (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14473__A (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14375__A1 (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14295__A (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__S (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__A2 (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12739__A2 (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__B (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12765__S (.DIODE(_06869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12763__S (.DIODE(_06869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__S (.DIODE(_06869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__S (.DIODE(_06869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__S (.DIODE(_06869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__S (.DIODE(_06869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__S (.DIODE(_06869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12751__S (.DIODE(_06869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__S (.DIODE(_06869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__S (.DIODE(_06869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__S (.DIODE(_06880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__S (.DIODE(_06880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__S (.DIODE(_06880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__S (.DIODE(_06880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__S (.DIODE(_06880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__S (.DIODE(_06880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__S (.DIODE(_06880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__S (.DIODE(_06880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__S (.DIODE(_06880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__S (.DIODE(_06880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__S (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12805__S (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12803__S (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__S (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__S (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__S (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12795__S (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__S (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12791__S (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__S (.DIODE(_06891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__S (.DIODE(_06906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12832__S (.DIODE(_06906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__S (.DIODE(_06906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__S (.DIODE(_06906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__S (.DIODE(_06906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__S (.DIODE(_06906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__S (.DIODE(_06906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__S (.DIODE(_06906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__S (.DIODE(_06906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12816__S (.DIODE(_06906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12855__S (.DIODE(_06917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__S (.DIODE(_06917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12851__S (.DIODE(_06917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12849__S (.DIODE(_06917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12847__S (.DIODE(_06917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12845__S (.DIODE(_06917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__S (.DIODE(_06917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12841__S (.DIODE(_06917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__S (.DIODE(_06917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12837__S (.DIODE(_06917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__S (.DIODE(_06928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12874__S (.DIODE(_06928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12872__S (.DIODE(_06928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12870__S (.DIODE(_06928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12868__S (.DIODE(_06928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12866__S (.DIODE(_06928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12864__S (.DIODE(_06928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12862__S (.DIODE(_06928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__S (.DIODE(_06928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__S (.DIODE(_06928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16677__A0 (.DIODE(_06941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16541__A0 (.DIODE(_06941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16405__A0 (.DIODE(_06941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16337__A0 (.DIODE(_06941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16268__A0 (.DIODE(_06941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__A0 (.DIODE(_06941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13188__A0 (.DIODE(_06941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13120__A0 (.DIODE(_06941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13052__A0 (.DIODE(_06941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12885__A0 (.DIODE(_06941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__S (.DIODE(_06943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12909__S (.DIODE(_06943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__S (.DIODE(_06943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12903__S (.DIODE(_06943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12900__S (.DIODE(_06943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__S (.DIODE(_06943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__S (.DIODE(_06943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12891__S (.DIODE(_06943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__S (.DIODE(_06943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12885__S (.DIODE(_06943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16681__A0 (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16545__A0 (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16409__A0 (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16341__A0 (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16272__A0 (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__A0 (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13192__A0 (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13124__A0 (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13056__A0 (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12891__A0 (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16683__A0 (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16547__A0 (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16411__A0 (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16343__A0 (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16274__A0 (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13262__A0 (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13194__A0 (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13126__A0 (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__A0 (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__A0 (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12943__S (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12940__S (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12937__S (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12934__S (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__S (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12928__S (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__S (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12922__S (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12919__S (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12916__S (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16702__A0 (.DIODE(_06968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16566__A0 (.DIODE(_06968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16430__A0 (.DIODE(_06968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16362__A0 (.DIODE(_06968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16293__A0 (.DIODE(_06968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13281__A0 (.DIODE(_06968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13213__A0 (.DIODE(_06968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13145__A0 (.DIODE(_06968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13077__A0 (.DIODE(_06968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12922__A0 (.DIODE(_06968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16708__A0 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16572__A0 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16436__A0 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16368__A0 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16299__A0 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13287__A0 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13219__A0 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__A0 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13083__A0 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__A0 (.DIODE(_06974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16714__A0 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16578__A0 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16442__A0 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16374__A0 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16305__A0 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13293__A0 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__A0 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__A0 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__A0 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12940__A0 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16719__A0 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16583__A0 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16447__A0 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16379__A0 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16310__A0 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13298__A0 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13230__A0 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__A0 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__A0 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12947__A0 (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__S (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__S (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__S (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__S (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__S (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__S (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__S (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__S (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12950__S (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12947__S (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16721__A0 (.DIODE(_06987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16585__A0 (.DIODE(_06987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16449__A0 (.DIODE(_06987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16381__A0 (.DIODE(_06987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16312__A0 (.DIODE(_06987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13300__A0 (.DIODE(_06987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13232__A0 (.DIODE(_06987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13164__A0 (.DIODE(_06987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13096__A0 (.DIODE(_06987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12950__A0 (.DIODE(_06987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16725__A0 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16589__A0 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16453__A0 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16385__A0 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16316__A0 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13304__A0 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13236__A0 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13168__A0 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13100__A0 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__A0 (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16733__A0 (.DIODE(_06999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16597__A0 (.DIODE(_06999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16461__A0 (.DIODE(_06999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16393__A0 (.DIODE(_06999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16324__A0 (.DIODE(_06999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__A0 (.DIODE(_06999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13244__A0 (.DIODE(_06999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__A0 (.DIODE(_06999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__A0 (.DIODE(_06999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__A0 (.DIODE(_06999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16741__A0 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16605__A0 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16469__A0 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16401__A0 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16332__A0 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__A0 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13252__A0 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13184__A0 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__A0 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__A0 (.DIODE(_07007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__S (.DIODE(_07009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__S (.DIODE(_07009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13025__A (.DIODE(_07009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__A (.DIODE(_07009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__A (.DIODE(_07009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__S (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__S (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__S (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__S (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__S (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__S (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__S (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12988__S (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__S (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__S (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__S (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13021__S (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__S (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__S (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__S (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13013__S (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__S (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13009__S (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13007__S (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13005__S (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__S (.DIODE(_07032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13042__S (.DIODE(_07032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13040__S (.DIODE(_07032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__S (.DIODE(_07032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__S (.DIODE(_07032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__S (.DIODE(_07032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__S (.DIODE(_07032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__S (.DIODE(_07032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__S (.DIODE(_07032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__S (.DIODE(_07032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__S (.DIODE(_07045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13114__S (.DIODE(_07045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__A (.DIODE(_07045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__A (.DIODE(_07045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__A (.DIODE(_07045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13070__S (.DIODE(_07046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13068__S (.DIODE(_07046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__S (.DIODE(_07046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__S (.DIODE(_07046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13062__S (.DIODE(_07046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__S (.DIODE(_07046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__S (.DIODE(_07046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13056__S (.DIODE(_07046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__S (.DIODE(_07046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13052__S (.DIODE(_07046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__S (.DIODE(_07057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__S (.DIODE(_07057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13087__S (.DIODE(_07057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__S (.DIODE(_07057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13083__S (.DIODE(_07057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__S (.DIODE(_07057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13079__S (.DIODE(_07057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13077__S (.DIODE(_07057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__S (.DIODE(_07057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13073__S (.DIODE(_07057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13112__S (.DIODE(_07068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13110__S (.DIODE(_07068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__S (.DIODE(_07068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13106__S (.DIODE(_07068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__S (.DIODE(_07068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13102__S (.DIODE(_07068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13100__S (.DIODE(_07068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__S (.DIODE(_07068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13096__S (.DIODE(_07068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__S (.DIODE(_07068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13184__S (.DIODE(_07081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__S (.DIODE(_07081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13161__A (.DIODE(_07081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13140__A (.DIODE(_07081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__A (.DIODE(_07081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13138__S (.DIODE(_07082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13136__S (.DIODE(_07082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__S (.DIODE(_07082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13132__S (.DIODE(_07082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__S (.DIODE(_07082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13128__S (.DIODE(_07082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13126__S (.DIODE(_07082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13124__S (.DIODE(_07082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13122__S (.DIODE(_07082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13120__S (.DIODE(_07082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13159__S (.DIODE(_07093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__S (.DIODE(_07093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__S (.DIODE(_07093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__S (.DIODE(_07093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__S (.DIODE(_07093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13149__S (.DIODE(_07093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__S (.DIODE(_07093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13145__S (.DIODE(_07093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13143__S (.DIODE(_07093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13141__S (.DIODE(_07093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__S (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13178__S (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__S (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__S (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__S (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13170__S (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13168__S (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13166__S (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13164__S (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__S (.DIODE(_07104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13206__S (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__S (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__S (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__S (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13198__S (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__S (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13194__S (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13192__S (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13190__S (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13188__S (.DIODE(_07118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13227__S (.DIODE(_07129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__S (.DIODE(_07129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13223__S (.DIODE(_07129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13221__S (.DIODE(_07129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13219__S (.DIODE(_07129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__S (.DIODE(_07129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13215__S (.DIODE(_07129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13213__S (.DIODE(_07129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13211__S (.DIODE(_07129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__S (.DIODE(_07129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13248__S (.DIODE(_07140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13246__S (.DIODE(_07140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13244__S (.DIODE(_07140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13242__S (.DIODE(_07140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13240__S (.DIODE(_07140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13238__S (.DIODE(_07140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13236__S (.DIODE(_07140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13234__S (.DIODE(_07140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13232__S (.DIODE(_07140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13230__S (.DIODE(_07140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__S (.DIODE(_07153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__S (.DIODE(_07153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13297__A (.DIODE(_07153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13276__A (.DIODE(_07153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13255__A (.DIODE(_07153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13274__S (.DIODE(_07154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13272__S (.DIODE(_07154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13270__S (.DIODE(_07154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13268__S (.DIODE(_07154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13266__S (.DIODE(_07154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13264__S (.DIODE(_07154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13262__S (.DIODE(_07154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__S (.DIODE(_07154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13258__S (.DIODE(_07154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__S (.DIODE(_07154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13295__S (.DIODE(_07165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13293__S (.DIODE(_07165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13291__S (.DIODE(_07165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13289__S (.DIODE(_07165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13287__S (.DIODE(_07165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13285__S (.DIODE(_07165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13283__S (.DIODE(_07165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13281__S (.DIODE(_07165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13279__S (.DIODE(_07165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13277__S (.DIODE(_07165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__S (.DIODE(_07176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13314__S (.DIODE(_07176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__S (.DIODE(_07176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13310__S (.DIODE(_07176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13308__S (.DIODE(_07176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13306__S (.DIODE(_07176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13304__S (.DIODE(_07176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13302__S (.DIODE(_07176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13300__S (.DIODE(_07176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13298__S (.DIODE(_07176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15656__A (.DIODE(_07208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14974__A (.DIODE(_07208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13345__A2_N (.DIODE(_07208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__A1 (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__A1 (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__A1 (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13442__A (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13418__A (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13400__A1 (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13386__A1 (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13343__B (.DIODE(_07209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__B1 (.DIODE(_07210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13604__B1 (.DIODE(_07210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13400__B1 (.DIODE(_07210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13367__B1 (.DIODE(_07210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13344__A (.DIODE(_07210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__B1 (.DIODE(_07211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__B1 (.DIODE(_07211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13576__A2 (.DIODE(_07211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__B1 (.DIODE(_07211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__B1 (.DIODE(_07211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__A2 (.DIODE(_07211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13443__A (.DIODE(_07211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__A (.DIODE(_07211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13386__B1 (.DIODE(_07211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13345__B1 (.DIODE(_07211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13731__C1 (.DIODE(_07217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13719__A1 (.DIODE(_07217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13686__C1 (.DIODE(_07217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13672__C1 (.DIODE(_07217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13630__B2 (.DIODE(_07217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13616__C1 (.DIODE(_07217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13601__C1 (.DIODE(_07217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__A1 (.DIODE(_07217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__A1 (.DIODE(_07217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13351__B1 (.DIODE(_07217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13803__C1 (.DIODE(_07221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__C1 (.DIODE(_07221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__C1 (.DIODE(_07221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13576__C1 (.DIODE(_07221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__C1 (.DIODE(_07221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__C1 (.DIODE(_07221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13476__C1 (.DIODE(_07221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__C1 (.DIODE(_07221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13420__A (.DIODE(_07221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13355__A2 (.DIODE(_07221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14887__B1 (.DIODE(_07224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13805__S (.DIODE(_07224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13794__S (.DIODE(_07224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13780__S (.DIODE(_07224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13750__S (.DIODE(_07224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13735__S (.DIODE(_07224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13723__S (.DIODE(_07224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13691__S (.DIODE(_07224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13408__A (.DIODE(_07224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13358__A (.DIODE(_07224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13761__B1 (.DIODE(_07225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13663__B1_N (.DIODE(_07225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13504__S (.DIODE(_07225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13478__S (.DIODE(_07225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13463__S (.DIODE(_07225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13446__S (.DIODE(_07225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13406__S (.DIODE(_07225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13393__S (.DIODE(_07225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13376__S (.DIODE(_07225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13359__S (.DIODE(_07225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13804__A1 (.DIODE(_07232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13777__C1 (.DIODE(_07232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13734__A1 (.DIODE(_07232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13721__A1 (.DIODE(_07232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13690__A1 (.DIODE(_07232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13631__C1 (.DIODE(_07232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13501__B1 (.DIODE(_07232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13404__A1 (.DIODE(_07232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13391__A1 (.DIODE(_07232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13374__A1 (.DIODE(_07232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15668__A1 (.DIODE(_07250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13386__A2 (.DIODE(_07250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13762__A2 (.DIODE(_07271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13704__A2 (.DIODE(_07271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13703__B1 (.DIODE(_07271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13664__A2 (.DIODE(_07271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13646__A2 (.DIODE(_07271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13645__B1 (.DIODE(_07271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13491__A2 (.DIODE(_07271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13490__B1 (.DIODE(_07271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13431__A2 (.DIODE(_07271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13430__B1 (.DIODE(_07271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16744__A2 (.DIODE(_07274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14892__B1 (.DIODE(_07274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13754__C1 (.DIODE(_07274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13695__A1 (.DIODE(_07274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13649__C1 (.DIODE(_07274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13637__A1 (.DIODE(_07274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13513__A1 (.DIODE(_07274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13501__A1 (.DIODE(_07274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13482__A1 (.DIODE(_07274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13412__C1 (.DIODE(_07274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13756__C1 (.DIODE(_07283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13733__C1 (.DIODE(_07283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13689__C1 (.DIODE(_07283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13675__C1 (.DIODE(_07283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13650__C1 (.DIODE(_07283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13618__C1 (.DIODE(_07283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13605__B2 (.DIODE(_07283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13502__C1 (.DIODE(_07283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13444__C1 (.DIODE(_07283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13421__A (.DIODE(_07283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13803__A1 (.DIODE(_07304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13792__A1 (.DIODE(_07304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__A1 (.DIODE(_07304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13733__A1 (.DIODE(_07304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13689__A1 (.DIODE(_07304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13675__A1 (.DIODE(_07304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13618__A1 (.DIODE(_07304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__A1 (.DIODE(_07304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13502__A1 (.DIODE(_07304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13444__A1 (.DIODE(_07304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13803__B1 (.DIODE(_07305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13792__B1 (.DIODE(_07305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13733__B1 (.DIODE(_07305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13689__B1 (.DIODE(_07305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13675__B1 (.DIODE(_07305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13618__B1 (.DIODE(_07305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__B1 (.DIODE(_07305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13502__B1 (.DIODE(_07305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13476__A2 (.DIODE(_07305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13444__B1 (.DIODE(_07305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15698__A1 (.DIODE(_07371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13515__A2 (.DIODE(_07371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13677__S (.DIODE(_07374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13633__S (.DIODE(_07374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__S (.DIODE(_07374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13607__S (.DIODE(_07374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__S (.DIODE(_07374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13578__S (.DIODE(_07374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13563__S (.DIODE(_07374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13549__S (.DIODE(_07374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13531__S (.DIODE(_07374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13518__S (.DIODE(_07374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13548__A2 (.DIODE(_07392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15717__A1 (.DIODE(_07441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__A2 (.DIODE(_07441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14876__B1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14867__B1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14691__B1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14116__B1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14103__B1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14039__B1 (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13889__A (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13886__A (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13883__A (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13880__A (.DIODE(_07675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13979__A2 (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13976__A2 (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13943__A (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13910__A (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13874__A (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14967__A1 (.DIODE(_07679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13877__A2 (.DIODE(_07679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13979__B1 (.DIODE(_07681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13976__B1 (.DIODE(_07681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13944__A (.DIODE(_07681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13911__A (.DIODE(_07681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13878__A (.DIODE(_07681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16261__A (.DIODE(_07737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14964__A (.DIODE(_07737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13980__A (.DIODE(_07737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13977__A (.DIODE(_07737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13974__A (.DIODE(_07737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13971__A (.DIODE(_07737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13968__A (.DIODE(_07737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13965__A (.DIODE(_07737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13962__A (.DIODE(_07737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13959__A (.DIODE(_07737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14605__A1 (.DIODE(_07754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14429__B (.DIODE(_07754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13983__B (.DIODE(_07754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14963__S (.DIODE(_07755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13991__D (.DIODE(_07755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13987__C (.DIODE(_07755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13985__A2 (.DIODE(_07755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13984__B (.DIODE(_07755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14030__B1 (.DIODE(_07759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14021__B1 (.DIODE(_07759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14010__B1 (.DIODE(_07759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14007__B1 (.DIODE(_07759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14004__B1 (.DIODE(_07759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14001__B1 (.DIODE(_07759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13998__B1 (.DIODE(_07759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13995__B1 (.DIODE(_07759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13992__B1 (.DIODE(_07759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13989__B1 (.DIODE(_07759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15713__C1 (.DIODE(_07775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15678__C1 (.DIODE(_07775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15675__C1 (.DIODE(_07775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15663__C1 (.DIODE(_07775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14133__C1 (.DIODE(_07775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14077__B1 (.DIODE(_07775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14067__B1 (.DIODE(_07775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14058__B1 (.DIODE(_07775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14023__B1 (.DIODE(_07775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14013__B1 (.DIODE(_07775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16264__B (.DIODE(_07778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15781__A (.DIODE(_07778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15743__A (.DIODE(_07778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15657__A (.DIODE(_07778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15634__A (.DIODE(_07778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14128__A (.DIODE(_07778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14062__B (.DIODE(_07778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14044__B (.DIODE(_07778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14027__B (.DIODE(_07778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14018__B (.DIODE(_07778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14094__B1 (.DIODE(_07790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14084__B1 (.DIODE(_07790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14075__B1 (.DIODE(_07790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14065__B1 (.DIODE(_07790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14056__B1 (.DIODE(_07790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14053__B1 (.DIODE(_07790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14050__B1 (.DIODE(_07790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14047__B1 (.DIODE(_07790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14037__B1 (.DIODE(_07790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14034__B1 (.DIODE(_07790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14704__B (.DIODE(_07815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14695__B (.DIODE(_07815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14180__B (.DIODE(_07815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14171__B (.DIODE(_07815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14149__B (.DIODE(_07815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14121__B (.DIODE(_07815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14108__B (.DIODE(_07815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14091__B (.DIODE(_07815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14081__B (.DIODE(_07815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14072__B (.DIODE(_07815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14737__B1 (.DIODE(_07826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14728__B1 (.DIODE(_07826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14719__B1 (.DIODE(_07826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14709__B1 (.DIODE(_07826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14700__B1 (.DIODE(_07826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14185__B1 (.DIODE(_07826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14176__B1 (.DIODE(_07826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14167__B1 (.DIODE(_07826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14144__B1 (.DIODE(_07826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14087__B1 (.DIODE(_07826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14155__B1 (.DIODE(_07834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14152__B1 (.DIODE(_07834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14142__B1 (.DIODE(_07834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14138__B1 (.DIODE(_07834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14135__B1 (.DIODE(_07834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14124__B1 (.DIODE(_07834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14114__B1 (.DIODE(_07834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14111__B1 (.DIODE(_07834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14101__B1 (.DIODE(_07834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14098__B1 (.DIODE(_07834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14735__B1 (.DIODE(_07877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14726__B1 (.DIODE(_07877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14717__B1 (.DIODE(_07877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14707__B1 (.DIODE(_07877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14698__B1 (.DIODE(_07877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14183__B1 (.DIODE(_07877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14174__B1 (.DIODE(_07877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14165__B1 (.DIODE(_07877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14162__B1 (.DIODE(_07877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14159__B1 (.DIODE(_07877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16207__B (.DIODE(_07898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__A1 (.DIODE(_07898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14607__C1 (.DIODE(_07898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14579__A1 (.DIODE(_07898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14553__A1 (.DIODE(_07898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__A1 (.DIODE(_07898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14523__A1 (.DIODE(_07898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14470__A1 (.DIODE(_07898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14452__A1 (.DIODE(_07898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14191__A (.DIODE(_07898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15779__A2 (.DIODE(_07899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14633__A1 (.DIODE(_07899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14497__A1 (.DIODE(_07899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14446__A1 (.DIODE(_07899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14434__A1 (.DIODE(_07899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14399__A1 (.DIODE(_07899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14388__B2 (.DIODE(_07899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14374__A1 (.DIODE(_07899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14258__A1 (.DIODE(_07899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14199__A1 (.DIODE(_07899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14332__A1 (.DIODE(_07901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14312__B1 (.DIODE(_07901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14235__B1 (.DIODE(_07901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14232__B1 (.DIODE(_07901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14221__A (.DIODE(_07901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14219__B1 (.DIODE(_07901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14216__B1 (.DIODE(_07901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14213__B1 (.DIODE(_07901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14201__A (.DIODE(_07901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14194__B1 (.DIODE(_07901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15649__D_N (.DIODE(_07904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__B1 (.DIODE(_07904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14649__B1 (.DIODE(_07904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14608__A2 (.DIODE(_07904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14579__B1 (.DIODE(_07904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14553__B1 (.DIODE(_07904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14535__A2 (.DIODE(_07904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14323__B1 (.DIODE(_07904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14256__A (.DIODE(_07904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14197__A (.DIODE(_07904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15779__B1 (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15647__A4 (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14549__B1 (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14526__B1 (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14474__B1 (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14388__A2 (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14338__B1 (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14265__A (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14227__A (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14198__A (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14279__A2 (.DIODE(_07906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14226__A2 (.DIODE(_07906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14224__A2 (.DIODE(_07906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14220__A2 (.DIODE(_07906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14217__A2 (.DIODE(_07906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14214__A2 (.DIODE(_07906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14211__A2 (.DIODE(_07906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14207__A2 (.DIODE(_07906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14203__A2 (.DIODE(_07906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14199__B1 (.DIODE(_07906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14493__A (.DIODE(_07934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14492__A1 (.DIODE(_07934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14471__A (.DIODE(_07934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14470__A2 (.DIODE(_07934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14464__B (.DIODE(_07934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14463__B (.DIODE(_07934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14240__B1 (.DIODE(_07934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14615__A (.DIODE(_07942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14528__B (.DIODE(_07942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14527__A1 (.DIODE(_07942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14281__B1 (.DIODE(_07942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14274__B1 (.DIODE(_07942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14272__B1 (.DIODE(_07942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14269__B1 (.DIODE(_07942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14266__B1 (.DIODE(_07942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14253__A (.DIODE(_07942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14251__B1 (.DIODE(_07942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14547__A (.DIODE(_07943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14545__A1 (.DIODE(_07943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14524__A (.DIODE(_07943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14523__A2 (.DIODE(_07943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14517__B (.DIODE(_07943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14516__B (.DIODE(_07943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14252__B1 (.DIODE(_07943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16263__A2 (.DIODE(_07944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14603__B1 (.DIODE(_07944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14534__B (.DIODE(_07944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14293__B1 (.DIODE(_07944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14290__B1 (.DIODE(_07944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14288__B1 (.DIODE(_07944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14286__B1 (.DIODE(_07944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14284__B1 (.DIODE(_07944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14278__B (.DIODE(_07944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14258__A2 (.DIODE(_07944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14632__A2 (.DIODE(_07947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14496__A2 (.DIODE(_07947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14452__B1 (.DIODE(_07947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14445__A2 (.DIODE(_07947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14433__A2 (.DIODE(_07947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14409__A2 (.DIODE(_07947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14398__A2 (.DIODE(_07947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14373__A2 (.DIODE(_07947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14360__A2 (.DIODE(_07947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14257__A (.DIODE(_07947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14688__A2 (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14666__A2 (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14644__A2 (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14624__A2 (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14574__A2 (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14510__A2 (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14484__A2 (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14423__A2 (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14348__A2 (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14258__B1 (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__A2 (.DIODE(_07950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14547__C (.DIODE(_07950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__A2 (.DIODE(_07950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14538__B (.DIODE(_07950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14537__B (.DIODE(_07950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14261__B1 (.DIODE(_07950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14581__A1 (.DIODE(_07952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14566__A2 (.DIODE(_07952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__B1 (.DIODE(_07952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14555__B (.DIODE(_07952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14553__A2 (.DIODE(_07952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14551__A (.DIODE(_07952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14550__A (.DIODE(_07952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14264__B1 (.DIODE(_07952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14587__A1 (.DIODE(_07954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14581__A2 (.DIODE(_07954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14580__A (.DIODE(_07954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14577__A2 (.DIODE(_07954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14572__A (.DIODE(_07954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14562__B (.DIODE(_07954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14561__A2 (.DIODE(_07954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14267__B1 (.DIODE(_07954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14587__A2 (.DIODE(_07956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14581__B1 (.DIODE(_07956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14580__B (.DIODE(_07956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14579__A2 (.DIODE(_07956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14575__B (.DIODE(_07956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14270__B1 (.DIODE(_07956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14613__A1 (.DIODE(_07958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14596__B (.DIODE(_07958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14594__A1 (.DIODE(_07958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14592__A (.DIODE(_07958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14591__A (.DIODE(_07958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14585__B (.DIODE(_07958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14584__B (.DIODE(_07958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14273__B1 (.DIODE(_07958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14613__A2 (.DIODE(_07959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14607__B1 (.DIODE(_07959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14600__B (.DIODE(_07959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14276__B1 (.DIODE(_07959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14510__B2 (.DIODE(_07960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14484__B2 (.DIODE(_07960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14361__A1 (.DIODE(_07960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14294__B2 (.DIODE(_07960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14291__B2 (.DIODE(_07960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14289__B2 (.DIODE(_07960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14287__B2 (.DIODE(_07960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14285__B2 (.DIODE(_07960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14282__B2 (.DIODE(_07960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14276__B2 (.DIODE(_07960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14637__A2 (.DIODE(_07964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14633__A2 (.DIODE(_07964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14628__B (.DIODE(_07964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14625__B (.DIODE(_07964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14282__B1 (.DIODE(_07964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14658__A1 (.DIODE(_07966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14651__A (.DIODE(_07966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14650__A1 (.DIODE(_07966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14646__A2 (.DIODE(_07966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14642__A (.DIODE(_07966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14636__B (.DIODE(_07966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14635__A2 (.DIODE(_07966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14285__B1 (.DIODE(_07966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14658__A2 (.DIODE(_07967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14651__B (.DIODE(_07967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14650__B1 (.DIODE(_07967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14649__A2 (.DIODE(_07967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14645__B (.DIODE(_07967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14287__B1 (.DIODE(_07967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14674__A (.DIODE(_07968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14673__A1 (.DIODE(_07968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14664__A (.DIODE(_07968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14661__B (.DIODE(_07968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14660__B (.DIODE(_07968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14656__A2 (.DIODE(_07968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14289__B1 (.DIODE(_07968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__A2 (.DIODE(_07969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14674__B (.DIODE(_07969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14673__B1 (.DIODE(_07969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14669__B (.DIODE(_07969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14668__B (.DIODE(_07969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14291__B1 (.DIODE(_07969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14684__B (.DIODE(_07971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14682__A3 (.DIODE(_07971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14681__A1 (.DIODE(_07971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14680__A (.DIODE(_07971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14679__A2 (.DIODE(_07971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14294__B1 (.DIODE(_07971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14544__B1_N (.DIODE(_07972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14508__A1 (.DIODE(_07972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14336__A (.DIODE(_07972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14314__A2 (.DIODE(_07972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14316__B (.DIODE(_07983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__B (.DIODE(_07983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15785__C (.DIODE(_07984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14605__A3 (.DIODE(_07984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14594__B2 (.DIODE(_07984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14362__B (.DIODE(_07984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14308__B (.DIODE(_07984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14681__B1 (.DIODE(_07986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14533__A1 (.DIODE(_07986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14494__A1 (.DIODE(_07986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14480__A1 (.DIODE(_07986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14454__B (.DIODE(_07986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14436__B1 (.DIODE(_07986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14379__A1 (.DIODE(_07986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14357__A1 (.DIODE(_07986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14310__B (.DIODE(_07986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14642__B (.DIODE(_07988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14611__A (.DIODE(_07988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14572__B (.DIODE(_07988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14548__A (.DIODE(_07988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14421__B (.DIODE(_07988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14347__A1 (.DIODE(_07988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14330__B1 (.DIODE(_07988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14313__A2 (.DIODE(_07988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15641__A1 (.DIODE(_07992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14596__C (.DIODE(_07992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14497__A3 (.DIODE(_07992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14482__A2 (.DIODE(_07992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14399__A3 (.DIODE(_07992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14374__A3 (.DIODE(_07992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14361__A3 (.DIODE(_07992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14318__A (.DIODE(_07992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15800__B (.DIODE(_07994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15640__A2 (.DIODE(_07994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14594__A2 (.DIODE(_07994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14494__B1 (.DIODE(_07994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14480__B1 (.DIODE(_07994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14397__A2 (.DIODE(_07994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14372__A2 (.DIODE(_07994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14357__B1 (.DIODE(_07994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14318__B (.DIODE(_07994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14656__B1 (.DIODE(_07997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14635__B1 (.DIODE(_07997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14622__B1 (.DIODE(_07997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14561__B1 (.DIODE(_07997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__B1 (.DIODE(_07997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14523__B1 (.DIODE(_07997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14412__B1 (.DIODE(_07997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14340__B1 (.DIODE(_07997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14326__B (.DIODE(_07997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14323__A2 (.DIODE(_07997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14655__A (.DIODE(_07998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14634__A (.DIODE(_07998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14622__A1 (.DIODE(_07998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14560__A (.DIODE(_07998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14545__B1 (.DIODE(_07998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14522__A (.DIODE(_07998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14469__A1 (.DIODE(_07998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14411__A (.DIODE(_07998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14339__A (.DIODE(_07998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14322__S (.DIODE(_07998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14665__A1_N (.DIODE(_08012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14643__A1 (.DIODE(_08012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__A1_N (.DIODE(_08012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14573__A1 (.DIODE(_08012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14521__B1_N (.DIODE(_08012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14483__A1 (.DIODE(_08012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14468__B1 (.DIODE(_08012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14422__A1 (.DIODE(_08012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14347__B2 (.DIODE(_08012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14337__B1 (.DIODE(_08012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15800__A (.DIODE(_08033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15798__S (.DIODE(_08033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14679__B1 (.DIODE(_08033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14632__B2 (.DIODE(_08033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14496__B2 (.DIODE(_08033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14445__B2 (.DIODE(_08033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14433__B2 (.DIODE(_08033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14398__B2 (.DIODE(_08033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14373__B2 (.DIODE(_08033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14360__B2 (.DIODE(_08033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14626__A (.DIODE(_08035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14605__B1 (.DIODE(_08035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14472__A (.DIODE(_08035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14431__A1 (.DIODE(_08035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14407__A1_N (.DIODE(_08035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14396__B2 (.DIODE(_08035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14371__A1 (.DIODE(_08035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14682__B1 (.DIODE(_08050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__A3 (.DIODE(_08050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14627__A (.DIODE(_08050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14579__A3 (.DIODE(_08050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14553__A3 (.DIODE(_08050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14508__B1 (.DIODE(_08050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14452__A3 (.DIODE(_08050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14446__A3 (.DIODE(_08050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14434__A3 (.DIODE(_08050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14379__B1 (.DIODE(_08050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14672__B1 (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14647__B1 (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14557__B1 (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14384__B1 (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14609__A1 (.DIODE(_08071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14589__B1 (.DIODE(_08071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14583__A1 (.DIODE(_08071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14536__A1 (.DIODE(_08071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14458__A1 (.DIODE(_08071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14410__A1 (.DIODE(_08071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14685__B1 (.DIODE(_08097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14630__B1 (.DIODE(_08097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14430__C1 (.DIODE(_08097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16066__A2 (.DIODE(_08232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15836__A1 (.DIODE(_08232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14684__A (.DIODE(_08232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14669__A (.DIODE(_08232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14668__A (.DIODE(_08232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14660__A (.DIODE(_08232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14658__B1 (.DIODE(_08232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14646__A1 (.DIODE(_08232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14637__B1 (.DIODE(_08232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14577__A1 (.DIODE(_08232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15706__A (.DIODE(_08335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14989__C1 (.DIODE(_08335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14987__C1 (.DIODE(_08335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14984__C1 (.DIODE(_08335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14982__C1 (.DIODE(_08335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14979__C1 (.DIODE(_08335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14977__C1 (.DIODE(_08335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14975__C1 (.DIODE(_08335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14969__A (.DIODE(_08335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14690__A (.DIODE(_08335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14794__B (.DIODE(_08350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14790__B (.DIODE(_08350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14784__B (.DIODE(_08350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14771__B (.DIODE(_08350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14762__B (.DIODE(_08350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14752__B (.DIODE(_08350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14741__B (.DIODE(_08350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14732__B (.DIODE(_08350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14723__B (.DIODE(_08350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14714__B (.DIODE(_08350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17921__D (.DIODE(_08380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17922__D (.DIODE(_08391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17923__D (.DIODE(_08394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17924__D (.DIODE(_08395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18136__D (.DIODE(\alu_out[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18137__D (.DIODE(\alu_out[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18139__D (.DIODE(\alu_out[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18140__D (.DIODE(\alu_out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18141__D (.DIODE(\alu_out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18127__D (.DIODE(\alu_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18146__D (.DIODE(\alu_out[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18148__D (.DIODE(\alu_out[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18149__D (.DIODE(\alu_out[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18154__D (.DIODE(\alu_out[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18128__D (.DIODE(\alu_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18157__D (.DIODE(\alu_out[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18129__D (.DIODE(\alu_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18130__D (.DIODE(\alu_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18131__D (.DIODE(\alu_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18132__D (.DIODE(\alu_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18133__D (.DIODE(\alu_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__A1 (.DIODE(\alu_out_q[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__A1 (.DIODE(\alu_out_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11617__A1 (.DIODE(\alu_out_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11628__A1 (.DIODE(\alu_out_q[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__A1 (.DIODE(\alu_out_q[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11645__A1 (.DIODE(\alu_out_q[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11654__A1 (.DIODE(\alu_out_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__A1 (.DIODE(\alu_out_q[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__A1 (.DIODE(\alu_out_q[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11681__A1 (.DIODE(\alu_out_q[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11690__A1 (.DIODE(\alu_out_q[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__A1 (.DIODE(\alu_out_q[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__A1 (.DIODE(\alu_out_q[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__A1 (.DIODE(\alu_out_q[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11753__A1 (.DIODE(\alu_out_q[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__A1 (.DIODE(\alu_out_q[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__A1 (.DIODE(\alu_out_q[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__A1 (.DIODE(\alu_out_q[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__A1 (.DIODE(\alu_out_q[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__A1 (.DIODE(\alu_out_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__A1 (.DIODE(\alu_out_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__A (.DIODE(\cpu_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__B (.DIODE(\cpu_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__B (.DIODE(\cpu_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__A (.DIODE(\cpu_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08499__C_N (.DIODE(\cpu_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__B1 (.DIODE(\cpu_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08491__A (.DIODE(\cpu_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A (.DIODE(\cpu_state[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16607__C_N (.DIODE(\cpuregs.waddr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__A1 (.DIODE(\cpuregs.waddr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12390__B (.DIODE(\cpuregs.waddr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__A (.DIODE(\cpuregs.waddr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12151__B (.DIODE(\cpuregs.waddr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__B_N (.DIODE(\cpuregs.waddr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11873__B (.DIODE(\cpuregs.waddr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__B (.DIODE(\cpuregs.waddr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__A_N (.DIODE(\cpuregs.waddr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16607__B (.DIODE(\cpuregs.waddr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__A1 (.DIODE(\cpuregs.waddr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12390__A (.DIODE(\cpuregs.waddr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__B_N (.DIODE(\cpuregs.waddr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12151__A (.DIODE(\cpuregs.waddr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__A (.DIODE(\cpuregs.waddr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11873__A (.DIODE(\cpuregs.waddr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__A (.DIODE(\cpuregs.waddr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__B (.DIODE(\cpuregs.waddr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16471__A_N (.DIODE(\cpuregs.waddr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16334__A_N (.DIODE(\cpuregs.waddr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__D (.DIODE(\cpuregs.waddr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__A_N (.DIODE(\cpuregs.waddr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__A1 (.DIODE(\cpuregs.waddr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__A (.DIODE(\cpuregs.waddr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A_N (.DIODE(\cpuregs.waddr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__A_N (.DIODE(\cpuregs.waddr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11874__A (.DIODE(\cpuregs.waddr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11510__A_N (.DIODE(\cpuregs.waddr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16013__A1 (.DIODE(\decoded_imm[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15075__B1 (.DIODE(\decoded_imm[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13381__A2 (.DIODE(\decoded_imm[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13365__A2 (.DIODE(\decoded_imm[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13363__B (.DIODE(\decoded_imm[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13347__A2 (.DIODE(\decoded_imm[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13346__A2 (.DIODE(\decoded_imm[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__B (.DIODE(\decoded_imm[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09308__B (.DIODE(\decoded_imm[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16043__A1 (.DIODE(\decoded_imm[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15269__A1 (.DIODE(\decoded_imm[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13541__B (.DIODE(\decoded_imm[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13523__A2 (.DIODE(\decoded_imm[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13507__B (.DIODE(\decoded_imm[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09736__B (.DIODE(\decoded_imm[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__B (.DIODE(\decoded_imm[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16046__A1 (.DIODE(\decoded_imm[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15285__A1 (.DIODE(\decoded_imm[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13542__A2 (.DIODE(\decoded_imm[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13521__B (.DIODE(\decoded_imm[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13520__B (.DIODE(\decoded_imm[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09814__B (.DIODE(\decoded_imm[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__B (.DIODE(\decoded_imm[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__B (.DIODE(\decoded_imm[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16049__A1 (.DIODE(\decoded_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15301__A1 (.DIODE(\decoded_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13544__B (.DIODE(\decoded_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13543__B (.DIODE(\decoded_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09812__B (.DIODE(\decoded_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__B (.DIODE(\decoded_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16051__A1 (.DIODE(\decoded_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15320__A1 (.DIODE(\decoded_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__B (.DIODE(\decoded_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13552__B (.DIODE(\decoded_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__B (.DIODE(\decoded_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09874__B (.DIODE(\decoded_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16053__A1 (.DIODE(\decoded_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15336__A1 (.DIODE(\decoded_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13566__B (.DIODE(\decoded_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13565__B (.DIODE(\decoded_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__B1 (.DIODE(\decoded_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__A2 (.DIODE(\decoded_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__B (.DIODE(\decoded_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16055__A1 (.DIODE(\decoded_imm[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15353__A1 (.DIODE(\decoded_imm[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13581__B (.DIODE(\decoded_imm[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13580__B (.DIODE(\decoded_imm[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09960__A2 (.DIODE(\decoded_imm[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__A2 (.DIODE(\decoded_imm[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__B (.DIODE(\decoded_imm[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16057__A1 (.DIODE(\decoded_imm[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15373__A1 (.DIODE(\decoded_imm[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13595__B (.DIODE(\decoded_imm[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__B (.DIODE(\decoded_imm[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__A2 (.DIODE(\decoded_imm[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__A2 (.DIODE(\decoded_imm[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__B (.DIODE(\decoded_imm[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16059__A1 (.DIODE(\decoded_imm[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15390__A1 (.DIODE(\decoded_imm[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13610__B (.DIODE(\decoded_imm[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13609__B (.DIODE(\decoded_imm[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10100__B (.DIODE(\decoded_imm[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09996__B (.DIODE(\decoded_imm[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__B (.DIODE(\decoded_imm[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16061__A1 (.DIODE(\decoded_imm[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15408__B2 (.DIODE(\decoded_imm[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13624__B (.DIODE(\decoded_imm[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13623__B (.DIODE(\decoded_imm[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__B (.DIODE(\decoded_imm[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10068__A2 (.DIODE(\decoded_imm[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10031__B (.DIODE(\decoded_imm[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16063__A1 (.DIODE(\decoded_imm[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15427__B2 (.DIODE(\decoded_imm[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13641__B (.DIODE(\decoded_imm[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13640__B (.DIODE(\decoded_imm[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__A2 (.DIODE(\decoded_imm[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__B (.DIODE(\decoded_imm[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10065__B (.DIODE(\decoded_imm[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16018__A1 (.DIODE(\decoded_imm[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15098__B1 (.DIODE(\decoded_imm[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13380__B (.DIODE(\decoded_imm[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13362__B (.DIODE(\decoded_imm[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13361__B (.DIODE(\decoded_imm[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09420__B (.DIODE(\decoded_imm[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__B (.DIODE(\decoded_imm[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__B (.DIODE(\decoded_imm[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16069__A1 (.DIODE(\decoded_imm[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15444__A1 (.DIODE(\decoded_imm[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13653__B (.DIODE(\decoded_imm[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13652__B (.DIODE(\decoded_imm[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__B (.DIODE(\decoded_imm[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__B (.DIODE(\decoded_imm[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16070__A1 (.DIODE(\decoded_imm[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15460__A1 (.DIODE(\decoded_imm[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13707__B (.DIODE(\decoded_imm[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13666__B (.DIODE(\decoded_imm[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13665__B (.DIODE(\decoded_imm[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__B (.DIODE(\decoded_imm[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__B (.DIODE(\decoded_imm[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16072__A1 (.DIODE(\decoded_imm[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15476__A1 (.DIODE(\decoded_imm[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13701__A2 (.DIODE(\decoded_imm[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13680__B (.DIODE(\decoded_imm[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13679__B (.DIODE(\decoded_imm[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__B (.DIODE(\decoded_imm[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10170__B (.DIODE(\decoded_imm[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16073__A1 (.DIODE(\decoded_imm[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15494__B2 (.DIODE(\decoded_imm[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13706__B (.DIODE(\decoded_imm[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13699__B (.DIODE(\decoded_imm[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13698__B (.DIODE(\decoded_imm[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__B (.DIODE(\decoded_imm[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__B (.DIODE(\decoded_imm[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10204__B (.DIODE(\decoded_imm[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16074__A1 (.DIODE(\decoded_imm[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15514__A1 (.DIODE(\decoded_imm[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13713__B (.DIODE(\decoded_imm[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13712__B (.DIODE(\decoded_imm[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10244__B (.DIODE(\decoded_imm[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__B (.DIODE(\decoded_imm[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16075__A1 (.DIODE(\decoded_imm[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15530__A1 (.DIODE(\decoded_imm[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13726__B (.DIODE(\decoded_imm[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13725__B (.DIODE(\decoded_imm[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__B (.DIODE(\decoded_imm[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__B (.DIODE(\decoded_imm[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16076__A1 (.DIODE(\decoded_imm[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15548__B2 (.DIODE(\decoded_imm[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13767__B1 (.DIODE(\decoded_imm[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13738__B (.DIODE(\decoded_imm[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13737__B (.DIODE(\decoded_imm[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__B (.DIODE(\decoded_imm[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__B (.DIODE(\decoded_imm[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16077__A1 (.DIODE(\decoded_imm[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15565__A1 (.DIODE(\decoded_imm[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13768__A2 (.DIODE(\decoded_imm[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13767__A2 (.DIODE(\decoded_imm[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13758__B (.DIODE(\decoded_imm[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__B (.DIODE(\decoded_imm[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__B (.DIODE(\decoded_imm[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10340__B (.DIODE(\decoded_imm[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16078__A1 (.DIODE(\decoded_imm[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15581__A1 (.DIODE(\decoded_imm[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13786__B (.DIODE(\decoded_imm[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13771__B (.DIODE(\decoded_imm[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13770__B (.DIODE(\decoded_imm[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10411__B (.DIODE(\decoded_imm[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__A2 (.DIODE(\decoded_imm[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__B (.DIODE(\decoded_imm[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16079__A1 (.DIODE(\decoded_imm[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15596__A1 (.DIODE(\decoded_imm[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13783__B (.DIODE(\decoded_imm[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13782__B (.DIODE(\decoded_imm[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__B (.DIODE(\decoded_imm[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__B (.DIODE(\decoded_imm[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16021__A1 (.DIODE(\decoded_imm[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15103__B1 (.DIODE(\decoded_imm[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13379__B (.DIODE(\decoded_imm[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13378__B (.DIODE(\decoded_imm[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09419__B (.DIODE(\decoded_imm[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__B (.DIODE(\decoded_imm[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16080__A1 (.DIODE(\decoded_imm[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15611__A1 (.DIODE(\decoded_imm[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13797__B (.DIODE(\decoded_imm[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13796__B (.DIODE(\decoded_imm[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10441__B (.DIODE(\decoded_imm[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__B (.DIODE(\decoded_imm[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16081__A1 (.DIODE(\decoded_imm[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15629__B2 (.DIODE(\decoded_imm[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14888__B (.DIODE(\decoded_imm[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__B (.DIODE(\decoded_imm[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16025__A1 (.DIODE(\decoded_imm[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15107__B1 (.DIODE(\decoded_imm[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__B (.DIODE(\decoded_imm[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13395__B (.DIODE(\decoded_imm[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09460__B (.DIODE(\decoded_imm[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__B (.DIODE(\decoded_imm[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16028__A1 (.DIODE(\decoded_imm[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15110__B1 (.DIODE(\decoded_imm[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13425__B (.DIODE(\decoded_imm[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__B (.DIODE(\decoded_imm[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__B (.DIODE(\decoded_imm[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__B (.DIODE(\decoded_imm[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16032__A1 (.DIODE(\decoded_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15155__A1 (.DIODE(\decoded_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__A2 (.DIODE(\decoded_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__B (.DIODE(\decoded_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13435__B (.DIODE(\decoded_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__B (.DIODE(\decoded_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__B (.DIODE(\decoded_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__B (.DIODE(\decoded_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16035__A1 (.DIODE(\decoded_imm[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15186__A1 (.DIODE(\decoded_imm[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13450__B (.DIODE(\decoded_imm[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13449__B (.DIODE(\decoded_imm[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__B (.DIODE(\decoded_imm[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__B (.DIODE(\decoded_imm[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16037__A1 (.DIODE(\decoded_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15206__B2 (.DIODE(\decoded_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13485__B (.DIODE(\decoded_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__B (.DIODE(\decoded_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13465__B (.DIODE(\decoded_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09628__B (.DIODE(\decoded_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__B (.DIODE(\decoded_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16039__A1 (.DIODE(\decoded_imm[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15228__A1 (.DIODE(\decoded_imm[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13540__A2 (.DIODE(\decoded_imm[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13495__A2 (.DIODE(\decoded_imm[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13487__B (.DIODE(\decoded_imm[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__B (.DIODE(\decoded_imm[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09664__B (.DIODE(\decoded_imm[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16041__A1 (.DIODE(\decoded_imm[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15248__A1 (.DIODE(\decoded_imm[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13506__B (.DIODE(\decoded_imm[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13493__B (.DIODE(\decoded_imm[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13492__B (.DIODE(\decoded_imm[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09726__B (.DIODE(\decoded_imm[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__B (.DIODE(\decoded_imm[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16045__A2 (.DIODE(\decoded_imm_j[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15822__B1 (.DIODE(\decoded_imm_j[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14438__A (.DIODE(\decoded_imm_j[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14437__A (.DIODE(\decoded_imm_j[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16048__A2 (.DIODE(\decoded_imm_j[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15823__A0 (.DIODE(\decoded_imm_j[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14460__A (.DIODE(\decoded_imm_j[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14448__A (.DIODE(\decoded_imm_j[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14447__A (.DIODE(\decoded_imm_j[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16050__A2 (.DIODE(\decoded_imm_j[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15826__A1 (.DIODE(\decoded_imm_j[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14464__A (.DIODE(\decoded_imm_j[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14463__A (.DIODE(\decoded_imm_j[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16052__A2 (.DIODE(\decoded_imm_j[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15827__A1 (.DIODE(\decoded_imm_j[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14476__A (.DIODE(\decoded_imm_j[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14475__A (.DIODE(\decoded_imm_j[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16054__A2 (.DIODE(\decoded_imm_j[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15828__A1 (.DIODE(\decoded_imm_j[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14486__A (.DIODE(\decoded_imm_j[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14485__A (.DIODE(\decoded_imm_j[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16056__A2 (.DIODE(\decoded_imm_j[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15829__A1 (.DIODE(\decoded_imm_j[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14514__A1 (.DIODE(\decoded_imm_j[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14503__A (.DIODE(\decoded_imm_j[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14502__A (.DIODE(\decoded_imm_j[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16058__A2 (.DIODE(\decoded_imm_j[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15831__A1 (.DIODE(\decoded_imm_j[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14517__A (.DIODE(\decoded_imm_j[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14516__A (.DIODE(\decoded_imm_j[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16060__A2 (.DIODE(\decoded_imm_j[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15833__A1 (.DIODE(\decoded_imm_j[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14528__A (.DIODE(\decoded_imm_j[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14527__B1 (.DIODE(\decoded_imm_j[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16062__A2 (.DIODE(\decoded_imm_j[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15835__A1 (.DIODE(\decoded_imm_j[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__A1 (.DIODE(\decoded_imm_j[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14538__A (.DIODE(\decoded_imm_j[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14537__A (.DIODE(\decoded_imm_j[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16034__A2 (.DIODE(\decoded_imm_j[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15812__A1 (.DIODE(\decoded_imm_j[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14381__A (.DIODE(\decoded_imm_j[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14380__A (.DIODE(\decoded_imm_j[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16036__A2 (.DIODE(\decoded_imm_j[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15814__A1 (.DIODE(\decoded_imm_j[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14390__A (.DIODE(\decoded_imm_j[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14389__A (.DIODE(\decoded_imm_j[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16038__A2 (.DIODE(\decoded_imm_j[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15815__A (.DIODE(\decoded_imm_j[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14416__A (.DIODE(\decoded_imm_j[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14403__A (.DIODE(\decoded_imm_j[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14402__A (.DIODE(\decoded_imm_j[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15879__B_N (.DIODE(decoder_trigger));
 sky130_fd_sc_hd__diode_2 ANTENNA__15850__B_N (.DIODE(decoder_trigger));
 sky130_fd_sc_hd__diode_2 ANTENNA__15639__A1 (.DIODE(decoder_trigger));
 sky130_fd_sc_hd__diode_2 ANTENNA__14315__A1 (.DIODE(decoder_trigger));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__B (.DIODE(decoder_trigger));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__A1 (.DIODE(decoder_trigger));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__B_N (.DIODE(decoder_trigger));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__C1 (.DIODE(decoder_trigger));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__A1 (.DIODE(decoder_trigger));
 sky130_fd_sc_hd__diode_2 ANTENNA__15858__B2 (.DIODE(instr_beq));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__A (.DIODE(instr_beq));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__A (.DIODE(instr_beq));
 sky130_fd_sc_hd__diode_2 ANTENNA__16066__A1 (.DIODE(instr_jal));
 sky130_fd_sc_hd__diode_2 ANTENNA__16031__A (.DIODE(instr_jal));
 sky130_fd_sc_hd__diode_2 ANTENNA__16015__A (.DIODE(instr_jal));
 sky130_fd_sc_hd__diode_2 ANTENNA__14429__A (.DIODE(instr_jal));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__A (.DIODE(instr_jal));
 sky130_fd_sc_hd__diode_2 ANTENNA__08601__A (.DIODE(instr_jal));
 sky130_fd_sc_hd__diode_2 ANTENNA__08587__A (.DIODE(instr_jal));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__C (.DIODE(instr_jal));
 sky130_fd_sc_hd__diode_2 ANTENNA__16088__C1 (.DIODE(instr_jalr));
 sky130_fd_sc_hd__diode_2 ANTENNA__16011__A (.DIODE(instr_jalr));
 sky130_fd_sc_hd__diode_2 ANTENNA__15877__A0 (.DIODE(instr_jalr));
 sky130_fd_sc_hd__diode_2 ANTENNA__15791__A2 (.DIODE(instr_jalr));
 sky130_fd_sc_hd__diode_2 ANTENNA__15632__B (.DIODE(instr_jalr));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__B (.DIODE(instr_jalr));
 sky130_fd_sc_hd__diode_2 ANTENNA__15842__A1 (.DIODE(instr_lui));
 sky130_fd_sc_hd__diode_2 ANTENNA__13343__A (.DIODE(instr_lui));
 sky130_fd_sc_hd__diode_2 ANTENNA__08473__B (.DIODE(instr_lui));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__A2 (.DIODE(instr_maskirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__09577__A (.DIODE(instr_maskirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__B (.DIODE(instr_maskirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__A (.DIODE(instr_maskirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__B (.DIODE(instr_maskirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__B1 (.DIODE(instr_rdcycleh));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__B1 (.DIODE(instr_rdcycleh));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__B1 (.DIODE(instr_rdcycleh));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__A1 (.DIODE(instr_rdcycleh));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A (.DIODE(instr_rdcycleh));
 sky130_fd_sc_hd__diode_2 ANTENNA__09280__A (.DIODE(instr_rdcycleh));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__C (.DIODE(instr_rdcycleh));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__B1 (.DIODE(instr_rdinstr));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__B1 (.DIODE(instr_rdinstr));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__B1 (.DIODE(instr_rdinstr));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__B1 (.DIODE(instr_rdinstr));
 sky130_fd_sc_hd__diode_2 ANTENNA__09608__B1 (.DIODE(instr_rdinstr));
 sky130_fd_sc_hd__diode_2 ANTENNA__09274__A (.DIODE(instr_rdinstr));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__B (.DIODE(instr_rdinstr));
 sky130_fd_sc_hd__diode_2 ANTENNA__13876__B (.DIODE(instr_retirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__10401__A1 (.DIODE(instr_retirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__A1 (.DIODE(instr_retirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__A1 (.DIODE(instr_retirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A (.DIODE(instr_retirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__09435__A (.DIODE(instr_retirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__09316__A (.DIODE(instr_retirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__C (.DIODE(instr_retirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__C (.DIODE(instr_retirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__15910__A1 (.DIODE(instr_slli));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__A2 (.DIODE(instr_slli));
 sky130_fd_sc_hd__diode_2 ANTENNA__10914__A2 (.DIODE(instr_slli));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__B (.DIODE(instr_slli));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__D (.DIODE(instr_slli));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__A1 (.DIODE(instr_sub));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__A (.DIODE(instr_sub));
 sky130_fd_sc_hd__diode_2 ANTENNA__11014__A1 (.DIODE(instr_sub));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__A (.DIODE(instr_sub));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__A (.DIODE(instr_sub));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__B (.DIODE(instr_sub));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__B2 (.DIODE(instr_timer));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__B2 (.DIODE(instr_timer));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__B2 (.DIODE(instr_timer));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__B2 (.DIODE(instr_timer));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__B2 (.DIODE(instr_timer));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__B2 (.DIODE(instr_timer));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A (.DIODE(instr_timer));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__A (.DIODE(instr_timer));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A (.DIODE(instr_timer));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__A (.DIODE(instr_timer));
 sky130_fd_sc_hd__diode_2 ANTENNA__15976__A0 (.DIODE(instr_waitirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__A_N (.DIODE(instr_waitirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__B1 (.DIODE(instr_waitirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__A (.DIODE(instr_waitirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__B1 (.DIODE(instr_waitirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__B (.DIODE(instr_waitirq));
 sky130_fd_sc_hd__diode_2 ANTENNA__14968__A1_N (.DIODE(irq_active));
 sky130_fd_sc_hd__diode_2 ANTENNA__14963__A1 (.DIODE(irq_active));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__B (.DIODE(irq_active));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__A2 (.DIODE(irq_active));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__A2 (.DIODE(irq_active));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__A (.DIODE(irq_active));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__B (.DIODE(irq_active));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__A2 (.DIODE(irq_active));
 sky130_fd_sc_hd__diode_2 ANTENNA__14977__A1 (.DIODE(\irq_mask[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__B (.DIODE(\irq_mask[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__A1 (.DIODE(\irq_mask[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__A1 (.DIODE(\irq_mask[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A_N (.DIODE(\irq_mask[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__A (.DIODE(\irq_mask[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14979__A1 (.DIODE(\irq_mask[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A1 (.DIODE(\irq_mask[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__A1 (.DIODE(\irq_mask[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__A (.DIODE(\irq_mask[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__A1 (.DIODE(\irq_mask[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__A_N (.DIODE(\irq_mask[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__A1 (.DIODE(\irq_mask[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14301__C (.DIODE(\irq_pending[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__A2 (.DIODE(\irq_pending[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__A1 (.DIODE(\irq_pending[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08554__B (.DIODE(\irq_pending[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14302__C (.DIODE(\irq_pending[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__A2 (.DIODE(\irq_pending[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A1 (.DIODE(\irq_pending[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__B (.DIODE(\irq_pending[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14302__D (.DIODE(\irq_pending[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11454__A2 (.DIODE(\irq_pending[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A1 (.DIODE(\irq_pending[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08577__B (.DIODE(\irq_pending[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14297__A (.DIODE(\irq_pending[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__A2 (.DIODE(\irq_pending[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__B2 (.DIODE(\irq_pending[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__B (.DIODE(\irq_pending[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14297__C (.DIODE(\irq_pending[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11460__A2 (.DIODE(\irq_pending[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__B2 (.DIODE(\irq_pending[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__B (.DIODE(\irq_pending[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14296__A (.DIODE(\irq_pending[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11464__A2 (.DIODE(\irq_pending[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__B2 (.DIODE(\irq_pending[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__B (.DIODE(\irq_pending[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14303__C (.DIODE(\irq_pending[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11434__A2 (.DIODE(\irq_pending[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09624__B1 (.DIODE(\irq_pending[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__B (.DIODE(\irq_pending[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15639__B1_N (.DIODE(\irq_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14254__A2 (.DIODE(\irq_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14209__A (.DIODE(\irq_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14192__B_N (.DIODE(\irq_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__A1 (.DIODE(\irq_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11497__A (.DIODE(\irq_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__B (.DIODE(\irq_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__B (.DIODE(\irq_state[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16100__B2 (.DIODE(is_alu_reg_imm));
 sky130_fd_sc_hd__diode_2 ANTENNA__16088__A1 (.DIODE(is_alu_reg_imm));
 sky130_fd_sc_hd__diode_2 ANTENNA__16011__C (.DIODE(is_alu_reg_imm));
 sky130_fd_sc_hd__diode_2 ANTENNA__15930__A (.DIODE(is_alu_reg_imm));
 sky130_fd_sc_hd__diode_2 ANTENNA__15913__A1 (.DIODE(is_alu_reg_imm));
 sky130_fd_sc_hd__diode_2 ANTENNA__15909__A (.DIODE(is_alu_reg_imm));
 sky130_fd_sc_hd__diode_2 ANTENNA__15897__B (.DIODE(is_alu_reg_imm));
 sky130_fd_sc_hd__diode_2 ANTENNA__15895__A1 (.DIODE(is_alu_reg_imm));
 sky130_fd_sc_hd__diode_2 ANTENNA__16105__A0 (.DIODE(is_alu_reg_reg));
 sky130_fd_sc_hd__diode_2 ANTENNA__15921__A1 (.DIODE(is_alu_reg_reg));
 sky130_fd_sc_hd__diode_2 ANTENNA__15914__B (.DIODE(is_alu_reg_reg));
 sky130_fd_sc_hd__diode_2 ANTENNA__16016__A (.DIODE(is_beq_bne_blt_bge_bltu_bgeu));
 sky130_fd_sc_hd__diode_2 ANTENNA__15791__A1 (.DIODE(is_beq_bne_blt_bge_bltu_bgeu));
 sky130_fd_sc_hd__diode_2 ANTENNA__15784__B_N (.DIODE(is_beq_bne_blt_bge_bltu_bgeu));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__A (.DIODE(is_beq_bne_blt_bge_bltu_bgeu));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__A (.DIODE(is_beq_bne_blt_bge_bltu_bgeu));
 sky130_fd_sc_hd__diode_2 ANTENNA__16085__A0 (.DIODE(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__diode_2 ANTENNA__16011__B (.DIODE(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__diode_2 ANTENNA__15890__A (.DIODE(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__diode_2 ANTENNA__15889__B2 (.DIODE(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__diode_2 ANTENNA__15886__B2 (.DIODE(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__diode_2 ANTENNA__15884__B2 (.DIODE(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__diode_2 ANTENNA__15642__A1 (.DIODE(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__A (.DIODE(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__A (.DIODE(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__diode_2 ANTENNA__16093__A1 (.DIODE(is_sb_sh_sw));
 sky130_fd_sc_hd__diode_2 ANTENNA__16044__A1 (.DIODE(is_sb_sh_sw));
 sky130_fd_sc_hd__diode_2 ANTENNA__16016__B (.DIODE(is_sb_sh_sw));
 sky130_fd_sc_hd__diode_2 ANTENNA__16012__A1 (.DIODE(is_sb_sh_sw));
 sky130_fd_sc_hd__diode_2 ANTENNA__15905__B2 (.DIODE(is_sb_sh_sw));
 sky130_fd_sc_hd__diode_2 ANTENNA__15894__B2 (.DIODE(is_sb_sh_sw));
 sky130_fd_sc_hd__diode_2 ANTENNA__15893__B2 (.DIODE(is_sb_sh_sw));
 sky130_fd_sc_hd__diode_2 ANTENNA__15642__B2 (.DIODE(is_sb_sh_sw));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__B2 (.DIODE(is_sb_sh_sw));
 sky130_fd_sc_hd__diode_2 ANTENNA__08623__A1 (.DIODE(is_sb_sh_sw));
 sky130_fd_sc_hd__diode_2 ANTENNA__15794__A1 (.DIODE(latched_branch));
 sky130_fd_sc_hd__diode_2 ANTENNA__14254__A1 (.DIODE(latched_branch));
 sky130_fd_sc_hd__diode_2 ANTENNA__14192__A (.DIODE(latched_branch));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__A1 (.DIODE(latched_branch));
 sky130_fd_sc_hd__diode_2 ANTENNA__11491__A (.DIODE(latched_branch));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__C1 (.DIODE(latched_branch));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A (.DIODE(latched_branch));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__A (.DIODE(latched_branch));
 sky130_fd_sc_hd__diode_2 ANTENNA__15798__A0 (.DIODE(latched_compr));
 sky130_fd_sc_hd__diode_2 ANTENNA__11518__A (.DIODE(latched_compr));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__B (.DIODE(latched_compr));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__A2 (.DIODE(latched_compr));
 sky130_fd_sc_hd__diode_2 ANTENNA__15788__A1 (.DIODE(latched_store));
 sky130_fd_sc_hd__diode_2 ANTENNA__14254__B1 (.DIODE(latched_store));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__A2 (.DIODE(latched_store));
 sky130_fd_sc_hd__diode_2 ANTENNA__11491__B_N (.DIODE(latched_store));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__B (.DIODE(latched_store));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__B (.DIODE(latched_store));
 sky130_fd_sc_hd__diode_2 ANTENNA__15643__A1 (.DIODE(mem_do_prefetch));
 sky130_fd_sc_hd__diode_2 ANTENNA__15633__A1 (.DIODE(mem_do_prefetch));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__A (.DIODE(mem_do_prefetch));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__A (.DIODE(mem_do_prefetch));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__B (.DIODE(mem_do_prefetch));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__B (.DIODE(mem_do_prefetch));
 sky130_fd_sc_hd__diode_2 ANTENNA__16109__A (.DIODE(mem_do_wdata));
 sky130_fd_sc_hd__diode_2 ANTENNA__15958__A (.DIODE(mem_do_wdata));
 sky130_fd_sc_hd__diode_2 ANTENNA__15650__B2 (.DIODE(mem_do_wdata));
 sky130_fd_sc_hd__diode_2 ANTENNA__15649__A (.DIODE(mem_do_wdata));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__A1 (.DIODE(mem_do_wdata));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__A (.DIODE(mem_do_wdata));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__A (.DIODE(mem_do_wdata));
 sky130_fd_sc_hd__diode_2 ANTENNA__08497__A1 (.DIODE(mem_do_wdata));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__A (.DIODE(mem_do_wdata));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__A1 (.DIODE(mem_do_wdata));
 sky130_fd_sc_hd__diode_2 ANTENNA__16024__B2 (.DIODE(\mem_rdata_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__A0 (.DIODE(\mem_rdata_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09010__A1 (.DIODE(\mem_rdata_q[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16027__B2 (.DIODE(\mem_rdata_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__A0 (.DIODE(\mem_rdata_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__A0 (.DIODE(\mem_rdata_q[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16069__B2 (.DIODE(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16012__B2 (.DIODE(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15944__A (.DIODE(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A0 (.DIODE(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09040__A1 (.DIODE(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16070__B2 (.DIODE(\mem_rdata_q[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16014__A (.DIODE(\mem_rdata_q[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15944__D_N (.DIODE(\mem_rdata_q[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15939__A (.DIODE(\mem_rdata_q[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__A0 (.DIODE(\mem_rdata_q[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09029__A1 (.DIODE(\mem_rdata_q[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16072__B2 (.DIODE(\mem_rdata_q[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16019__A (.DIODE(\mem_rdata_q[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15944__B (.DIODE(\mem_rdata_q[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15939__B (.DIODE(\mem_rdata_q[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09119__A0 (.DIODE(\mem_rdata_q[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__A0 (.DIODE(\mem_rdata_q[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16073__B2 (.DIODE(\mem_rdata_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16023__A (.DIODE(\mem_rdata_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15944__C (.DIODE(\mem_rdata_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15939__C (.DIODE(\mem_rdata_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__A0 (.DIODE(\mem_rdata_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__A0 (.DIODE(\mem_rdata_q[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16074__B2 (.DIODE(\mem_rdata_q[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16026__A (.DIODE(\mem_rdata_q[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15932__B_N (.DIODE(\mem_rdata_q[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09145__A0 (.DIODE(\mem_rdata_q[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09066__A0 (.DIODE(\mem_rdata_q[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16075__B2 (.DIODE(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16033__A1 (.DIODE(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15971__A (.DIODE(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15941__B (.DIODE(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15907__B (.DIODE(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__A0 (.DIODE(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__A1 (.DIODE(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16076__B2 (.DIODE(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16034__B2 (.DIODE(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15978__B_N (.DIODE(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15973__A1 (.DIODE(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15942__B_N (.DIODE(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15907__C (.DIODE(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__A0 (.DIODE(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__A1 (.DIODE(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16077__B2 (.DIODE(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16036__B2 (.DIODE(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15978__C (.DIODE(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15972__A (.DIODE(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15942__C (.DIODE(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15907__D (.DIODE(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__A0 (.DIODE(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08997__A0 (.DIODE(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16078__B2 (.DIODE(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16038__B2 (.DIODE(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15970__B (.DIODE(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15941__A (.DIODE(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15907__A (.DIODE(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09248__A0 (.DIODE(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__A1 (.DIODE(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16079__B2 (.DIODE(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16040__B2 (.DIODE(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15932__A_N (.DIODE(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15918__A (.DIODE(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15906__A (.DIODE(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__A0 (.DIODE(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08982__A0 (.DIODE(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16251__A0 (.DIODE(\mem_rdata_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15970__A (.DIODE(\mem_rdata_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15950__B (.DIODE(\mem_rdata_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15934__A (.DIODE(\mem_rdata_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09050__A1 (.DIODE(\mem_rdata_q[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16080__B2 (.DIODE(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16042__B2 (.DIODE(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15932__D (.DIODE(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15931__B2 (.DIODE(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15920__A (.DIODE(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15906__B (.DIODE(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__A0 (.DIODE(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__A0 (.DIODE(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16081__B2 (.DIODE(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16066__B2 (.DIODE(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16047__A1 (.DIODE(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16044__B1 (.DIODE(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15932__C (.DIODE(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15918__B (.DIODE(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15906__C (.DIODE(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A0 (.DIODE(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__A0 (.DIODE(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16045__B1 (.DIODE(\mem_rdata_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16012__A2 (.DIODE(\mem_rdata_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__A0 (.DIODE(\mem_rdata_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09058__A1 (.DIODE(\mem_rdata_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16020__B2 (.DIODE(\mem_rdata_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__A0 (.DIODE(\mem_rdata_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09061__A1 (.DIODE(\mem_rdata_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16264__A (.DIODE(\reg_next_pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13345__B2 (.DIODE(\reg_next_pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11502__B1 (.DIODE(\reg_next_pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__A (.DIODE(\reg_next_pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09308__A (.DIODE(\reg_next_pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__A (.DIODE(\reg_next_pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14445__A1 (.DIODE(\reg_next_pc[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14232__A1 (.DIODE(\reg_next_pc[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11619__A2 (.DIODE(\reg_next_pc[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__A0 (.DIODE(\reg_next_pc[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14484__A1 (.DIODE(\reg_next_pc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14242__A1 (.DIODE(\reg_next_pc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__A2 (.DIODE(\reg_next_pc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A0 (.DIODE(\reg_next_pc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14496__A1 (.DIODE(\reg_next_pc[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14245__A1 (.DIODE(\reg_next_pc[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A2 (.DIODE(\reg_next_pc[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11253__A0 (.DIODE(\reg_next_pc[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14510__A1 (.DIODE(\reg_next_pc[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14248__A1 (.DIODE(\reg_next_pc[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__A2 (.DIODE(\reg_next_pc[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__A0 (.DIODE(\reg_next_pc[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14535__A1 (.DIODE(\reg_next_pc[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14255__B2 (.DIODE(\reg_next_pc[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11683__A2 (.DIODE(\reg_next_pc[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__A0 (.DIODE(\reg_next_pc[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14323__B2 (.DIODE(\reg_next_pc[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11516__A2 (.DIODE(\reg_next_pc[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__A (.DIODE(\reg_next_pc[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14553__B2 (.DIODE(\reg_next_pc[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14263__A1 (.DIODE(\reg_next_pc[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11702__A2 (.DIODE(\reg_next_pc[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11279__A0 (.DIODE(\reg_next_pc[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14574__A1 (.DIODE(\reg_next_pc[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__A2 (.DIODE(\reg_next_pc[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__A (.DIODE(\reg_next_pc[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14579__B2 (.DIODE(\reg_next_pc[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14269__A1 (.DIODE(\reg_next_pc[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__A2 (.DIODE(\reg_next_pc[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11290__A0 (.DIODE(\reg_next_pc[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14632__A1 (.DIODE(\reg_next_pc[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14281__A1 (.DIODE(\reg_next_pc[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__A2 (.DIODE(\reg_next_pc[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__A0 (.DIODE(\reg_next_pc[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14644__A1 (.DIODE(\reg_next_pc[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14284__A1 (.DIODE(\reg_next_pc[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__A2 (.DIODE(\reg_next_pc[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11317__A0 (.DIODE(\reg_next_pc[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14649__B2 (.DIODE(\reg_next_pc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__A2 (.DIODE(\reg_next_pc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11323__A (.DIODE(\reg_next_pc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14338__B2 (.DIODE(\reg_next_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14200__A0 (.DIODE(\reg_next_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11530__A2 (.DIODE(\reg_next_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__A0 (.DIODE(\reg_next_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__B2 (.DIODE(\reg_next_pc[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__A2 (.DIODE(\reg_next_pc[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11334__A (.DIODE(\reg_next_pc[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14348__A1 (.DIODE(\reg_next_pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14205__A1 (.DIODE(\reg_next_pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__A2 (.DIODE(\reg_next_pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__A0 (.DIODE(\reg_next_pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__A0 (.DIODE(\reg_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14258__B2 (.DIODE(\reg_pc[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13622__B2 (.DIODE(\reg_pc[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11679__B1 (.DIODE(\reg_pc[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__A (.DIODE(\reg_pc[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__A (.DIODE(\reg_pc[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10068__A1 (.DIODE(\reg_pc[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10031__A (.DIODE(\reg_pc[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14276__A1 (.DIODE(\reg_pc[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__B2 (.DIODE(\reg_pc[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__B1 (.DIODE(\reg_pc[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11733__A (.DIODE(\reg_pc[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10244__A (.DIODE(\reg_pc[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__A (.DIODE(\reg_pc[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14279__A1 (.DIODE(\reg_pc[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13733__B2 (.DIODE(\reg_pc[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__A2 (.DIODE(\reg_pc[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11743__A1 (.DIODE(\reg_pc[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__A (.DIODE(\reg_pc[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__A (.DIODE(\reg_pc[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__A (.DIODE(\reg_pc[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14282__A1 (.DIODE(\reg_pc[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__B2 (.DIODE(\reg_pc[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__A1 (.DIODE(\reg_pc[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11759__B (.DIODE(\reg_pc[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11752__A1 (.DIODE(\reg_pc[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11751__A1 (.DIODE(\reg_pc[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__A (.DIODE(\reg_pc[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__A (.DIODE(\reg_pc[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14285__A1 (.DIODE(\reg_pc[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13756__B2 (.DIODE(\reg_pc[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__B1 (.DIODE(\reg_pc[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11759__A (.DIODE(\reg_pc[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__A (.DIODE(\reg_pc[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__A (.DIODE(\reg_pc[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10340__A (.DIODE(\reg_pc[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14287__A1 (.DIODE(\reg_pc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__B2 (.DIODE(\reg_pc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__B (.DIODE(\reg_pc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__A1 (.DIODE(\reg_pc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__A (.DIODE(\reg_pc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10411__A (.DIODE(\reg_pc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__A1 (.DIODE(\reg_pc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__A (.DIODE(\reg_pc[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14289__A1 (.DIODE(\reg_pc[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13792__B2 (.DIODE(\reg_pc[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11778__A1 (.DIODE(\reg_pc[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__A (.DIODE(\reg_pc[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__A (.DIODE(\reg_pc[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A (.DIODE(\reg_pc[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14211__A1 (.DIODE(\reg_pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13422__B2 (.DIODE(\reg_pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__A (.DIODE(\reg_pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__A (.DIODE(\reg_pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__A (.DIODE(\reg_pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__A (.DIODE(\reg_pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14224__A1 (.DIODE(\reg_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13483__B2 (.DIODE(\reg_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__A1 (.DIODE(\reg_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__B (.DIODE(\reg_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__A (.DIODE(\reg_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__A (.DIODE(\reg_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09664__A (.DIODE(\reg_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__C1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__B1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11450__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11454__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11460__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11464__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11428__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11430__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11432__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11434__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11436__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__16211__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__16205__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09010__A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__A0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09532__A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__08983__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__16215__A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__08416__A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__16217__A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10027__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__16219__A0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__A0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__16221__A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__16211__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__16205__A3 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__16223__A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10133__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09040__A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__16225__A0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09029__A0 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__16227__A0 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__16229__A0 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__16231__A0 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09696__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09066__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__16233__A0 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09730__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__A0 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__16235__A0 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__A0 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__16237__A0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10368__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__08997__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__16239__A0 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__A0 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__16241__A0 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09532__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__08982__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09050__A0 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__16243__A0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__16245__A0 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09632__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09045__A0 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__A0 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09030__A0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09058__A0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09696__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__A0 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09730__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__A0 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09061__A0 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__15963__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__A_N (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__15952__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__C (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__13381__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__C1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08844__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08770__A_N (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08460__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08459__B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__13541__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__13507__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__A3 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__A0 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09740__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__13542__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__13521__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__13520__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__A0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__13544__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__13543__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__A3 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A3 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__08791__B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__13552__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08792__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08728__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__13566__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__13565__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08795__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08726__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__13581__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__13580__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__09921__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08797__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08724__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__13595__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09988__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__B_N (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08718__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__13610__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__13609__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__10933__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__10025__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08800__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__13624__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__13623__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__10036__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__B_N (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08714__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__13641__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__13640__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10602__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__08711__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__08710__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__13380__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__13362__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__B_N (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08458__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__13653__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__13652__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10602__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10132__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08698__B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__13680__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__13679__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__A3 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08812__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__13706__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__13699__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__13698__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__13713__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__13712__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08819__B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08692__B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__13725__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08818__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08688__B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__13767__C1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__13738__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__13737__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10609__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__13768__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__13767__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__13758__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__13771__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__13770__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10570__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08828__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__13783__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__13782__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10570__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08678__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08677__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__13379__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__13378__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__A3 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__B (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__B (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__B (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08766__B (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08829__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__08830__B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__08666__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__13395__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__09465__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08840__B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__13425__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A3 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08762__B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08761__B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__13450__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__13449__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10788__A3 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10743__A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09612__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__13485__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08752__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__13493__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__13492__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10788__A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A0 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__08747__B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__18726__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08770__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__15270__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__A_N (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08739__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__15286__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__15302__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08791__A_N (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__15321__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__08792__A_N (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__08728__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__15337__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08795__A_N (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08726__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__15354__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08797__A_N (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08724__B_N (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__15374__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08718__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__15391__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__10933__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08801__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__15409__A0 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08714__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__15428__A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08711__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08710__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__18727__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__15445__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08698__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__15461__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10994__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08810__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08696__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__15477__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11160__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08812__A_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__15495__A0 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__15515__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08819__A_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08692__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__15531__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08688__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__15549__A0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__A_N (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__15566__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__15582__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__11173__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__15597__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__A_N (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08678__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08677__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__18728__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__A_N (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08766__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__15612__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08829__A_N (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__15630__A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08830__A_N (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08666__B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18729__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08764__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__18730__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__A_N (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08762__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08761__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__18731__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__16131__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__15156__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__A0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__18732__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__16133__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__15187__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__11160__A0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__A_N (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__18733__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__16135__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__15207__A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08848__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__15229__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08784__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08743__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__15249__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__A_N (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08747__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__13954__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__13961__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__13964__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_output154_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__13976__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__13979__B2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__14943__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_output176_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__14945__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__14947__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_output178_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__14949__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_output179_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__14951__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_output180_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__14953__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_output181_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__14955__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_output182_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__14957__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_output184_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__14959__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_output185_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__14961__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_output193_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__16113__B2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_output194_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__14917__A0 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_output195_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__14919__A0 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_output196_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__14922__A0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_output197_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__14924__A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_output198_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__14926__A0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_output199_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__14928__A0 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_output200_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__14930__A0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_output201_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__14932__A0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_output202_A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__14934__A0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_output203_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__14936__A0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_output204_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__14938__A0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_output205_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__14940__A0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_output206_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__14943__A0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_output207_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__14945__A0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_output208_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__14947__A0 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_output209_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__14949__A0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_output210_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__14951__A0 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_output211_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__14953__A0 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_output212_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__14955__A0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_output213_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__14957__A0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_output214_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__14901__A0 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_output215_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__14959__A0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_output216_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__14961__A0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_output217_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__14903__A0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_output218_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__14905__A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_output219_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__14907__A0 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_output220_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__14909__A0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_output221_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__14911__A0 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_output222_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__14913__A0 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_output223_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__14915__A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_output224_A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__15964__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__14898__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_output226_A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__16142__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_output227_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__16144__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_output228_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__16146__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_output229_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__16148__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_output230_A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__16150__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_output231_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__16152__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_output232_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__16154__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_output233_A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__16156__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_output234_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__16159__A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_output235_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__16161__A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_output237_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__16163__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_output238_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__16165__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_output239_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__16167__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_output240_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__16169__A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_output241_A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__16171__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_output242_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__16173__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_output243_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__16175__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_output244_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__16177__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_output245_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__16179__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_output246_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__16181__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_output248_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__16183__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_output249_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__16185__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_output255_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__16138__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_output256_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__16140__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_output257_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__16197__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__16195__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__16192__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__16188__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__14898__B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_output258_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__16188__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_output259_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__16192__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_output260_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__16195__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_output261_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__16197__A2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_output262_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__15968__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_output263_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__16121__A0 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_output288_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__16127__A0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_output299_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__16206__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__15954__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__15952__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__14897__B (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__B1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09837__C1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__B1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__B1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap300_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__B1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_191_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_190_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_189_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_188_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_187_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_173_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_186_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_185_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_184_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_183_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_182_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_181_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_180_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_179_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_178_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_177_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_176_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_175_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_174_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_169_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_172_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_171_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_170_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_168_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_167_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_166_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_165_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_163_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_159_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_158_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_157_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_156_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_155_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_154_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_153_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_152_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_151_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_150_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_149_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_148_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_147_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_146_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_145_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_144_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_143_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_142_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_141_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_140_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_139_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_138_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_137_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_136_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_135_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_134_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_133_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_132_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_131_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_164_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_162_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_161_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_160_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_115_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_114_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_113_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_112_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_111_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_110_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_130_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_129_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_128_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_127_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_126_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_125_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_124_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_123_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_122_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_121_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_120_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_119_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_118_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_117_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_116_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_108_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_104_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_101_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_98_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_01990_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_01992_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_02070_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_02166_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_02166_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_03351_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_03428_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_03826_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_03979_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_04065_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_04151_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_04271_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_04397_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_04570_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_04637_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_04743_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_04923_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_04982_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_05313_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_05342_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_05864_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_05864_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_06141_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_07154_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_07944_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(\decoded_imm[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\decoded_imm[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\decoded_imm[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\decoded_imm[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\decoded_imm_j[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(is_alu_reg_reg));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(mem_do_wdata));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(\mem_rdata_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(\reg_next_pc[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_01908_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_01968_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(_03880_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(_04287_));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(_04575_));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(_04754_));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(_05929_));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_07057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(\decoded_imm[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(\reg_next_pc[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_01753_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(_05517_));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(_04342_));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net93));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_812 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_927 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1021 ();
 assign cpi_insn[0] = net302;
 assign cpi_insn[10] = net312;
 assign cpi_insn[11] = net313;
 assign cpi_insn[12] = net314;
 assign cpi_insn[13] = net315;
 assign cpi_insn[14] = net316;
 assign cpi_insn[15] = net317;
 assign cpi_insn[16] = net318;
 assign cpi_insn[17] = net319;
 assign cpi_insn[18] = net320;
 assign cpi_insn[19] = net321;
 assign cpi_insn[1] = net303;
 assign cpi_insn[20] = net322;
 assign cpi_insn[21] = net323;
 assign cpi_insn[22] = net324;
 assign cpi_insn[23] = net325;
 assign cpi_insn[24] = net326;
 assign cpi_insn[25] = net327;
 assign cpi_insn[26] = net328;
 assign cpi_insn[27] = net329;
 assign cpi_insn[28] = net330;
 assign cpi_insn[29] = net331;
 assign cpi_insn[2] = net304;
 assign cpi_insn[30] = net332;
 assign cpi_insn[31] = net333;
 assign cpi_insn[3] = net305;
 assign cpi_insn[4] = net306;
 assign cpi_insn[5] = net307;
 assign cpi_insn[6] = net308;
 assign cpi_insn[7] = net309;
 assign cpi_insn[8] = net310;
 assign cpi_insn[9] = net311;
 assign cpi_valid = net334;
 assign mem_addr[0] = net335;
 assign mem_addr[1] = net336;
 assign mem_la_addr[0] = net337;
 assign mem_la_addr[1] = net338;
 assign trace_data[0] = net339;
 assign trace_data[10] = net349;
 assign trace_data[11] = net350;
 assign trace_data[12] = net351;
 assign trace_data[13] = net352;
 assign trace_data[14] = net353;
 assign trace_data[15] = net354;
 assign trace_data[16] = net355;
 assign trace_data[17] = net356;
 assign trace_data[18] = net357;
 assign trace_data[19] = net358;
 assign trace_data[1] = net340;
 assign trace_data[20] = net359;
 assign trace_data[21] = net360;
 assign trace_data[22] = net361;
 assign trace_data[23] = net362;
 assign trace_data[24] = net363;
 assign trace_data[25] = net364;
 assign trace_data[26] = net365;
 assign trace_data[27] = net366;
 assign trace_data[28] = net367;
 assign trace_data[29] = net368;
 assign trace_data[2] = net341;
 assign trace_data[30] = net369;
 assign trace_data[31] = net370;
 assign trace_data[32] = net371;
 assign trace_data[33] = net372;
 assign trace_data[34] = net373;
 assign trace_data[35] = net374;
 assign trace_data[3] = net342;
 assign trace_data[4] = net343;
 assign trace_data[5] = net344;
 assign trace_data[6] = net345;
 assign trace_data[7] = net346;
 assign trace_data[8] = net347;
 assign trace_data[9] = net348;
 assign trace_valid = net375;
endmodule
